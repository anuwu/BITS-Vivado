`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qbCebIw2n8+gN2UzOmh7axnoM4dwT2xHCHsKSFB0KAVTaTY3VeBTwlUpMviyYkfKO23wp8O7SpGs
0Wn95oRYAQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MOTbFTv/+AMs8CgHaCOhzDGjJY2CXbGvrGa3rJLL400WolIwHStE0ZS9HCf5QwC/qlTKHtSKXPFo
IKgluTeQifTssmpfL3kRH0S67h8DFhFcVbDg7MudxUvt52DgkYpYAzVfSG/nUYQr0UoPZOGdWNek
d5BNE54QoixjvjzvCn0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GWCTcTUIemqhsdR62OeZRXGpfrf7+14v/PYnlQE2+elD/5AQSNezw8Yh5LK7/U0UILMPApnh3/AH
E8gsLq5Dk9JFecIp+TrRarBrPzdkLyp/yDQZefDHIVKK2//cPrCux9IXp+jQExTJ/wMgB3Pk/8bX
EXcTuij9bNakvhh0qqcvPXbXX9LL1qrTKljruNhZ8fj+nzA6ZReUIHP58Y7Ee1d3Xsop4p9lwil6
6qwN+Lhx0npqK6UrnqNlAIb5F4pmCfRi3mvh8/WO2vx/mksFcUOTOjcUSOA9S4Cc2fWFZaEJu2Jk
nSdbTDU9JPBBG1HOZLBI4PeIS07u4kvjL8YxuA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWqfi4eW93XaurdUTFdBvYmgRlNt3IP2HZZVV3EH4zpzhLtjfG9ITAAZ2wgVBZ/ubHVDQNx+f74V
7yqRHt9FI2nIXks1MGER0/CZXcSrokzmAY5FFnm9jVBaptM3nivib//wb+pTYDyqkgJnA/Lik/xE
5N+mBusMskQJf94X2yznI3BP0RzkvftwacL0/QByYbp8e6B4oEzsoFkwinZKNJ2vNWKLPcxUvmlb
PGne9+10W8+J83DqAyg/K8zGYWdHwirFkQalIXh13D6lOtBVr0AzGpUUavift5/tIqjagi8Vba05
wcVi1W96tvqzhLckg0QwF4ZrgLFtGXEYBLEWwA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T2Je2NpQz222u+FkFMUb+rWAcPEE4CQIHwQeLw0xXMrIAVVpaq5m32NeZx1nQkTHVHeERS6BRWqE
5KXKZ5QH/IVcY6HLPbXO3Dm2EHobkpU16emyCApLCsUgcmA/MRWQ1gDfMjS3AeaVHULoQYQW5w5d
K0sQnMkknyB54GHQXbQ9LDcdo6L8t0/QgEyTJQzA+Bh1kz6FgmgpxVnJ2LlXH2CxQ9jph4sAcht8
4D4AliecDgulrafA2JbdAEK/+S1BpiG4ACtXDtpGUomy9jKwXZ35RlimisNF6bqfSQIV4R/H0ItO
J5XFboxTqNvqI4emJgnLzw49Fg7ZKbuwP+cntw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eAGLDWmORjuQiifMQjmPS2N5D50nOZvLtva+eMzhWZqeQDnHdoI+D/Z7CnebSoJv86oC3voi3uQO
SxQ9InTJFQxtvUyucyRaLG3IUGvvgRJVL9/LE3scUCA2tTEFitvwjYXYvUghUxVeN0l5sMqzky5n
zjDXmH8VKNGD/5c9uPE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HEgtpre6H4t2Ov3YueDpHwa/86EaHsc4/+NjKCU7D9Yxbmaq3EsfTvD4TQrIFaVgkWk0x47Z+GXZ
XP5UWE6u3RBO1x/Mh6hoOs07p3vW8f4+CpkxsVphw/PlJLMA6ViCtY1RT/gVyW3EMzdsWyMhYd0a
eBNyTGx/qVPHDSwhb68iLOncdRos4xvixfgQDHKuQsNL+3IolnroIGIVLQcbMlcya/UeqXPqMG2Q
D34oUJHsZe9pFr0sH47g3KLSIk5+85C9v/KjDCDxxt+J5rehkZYhGiFA7BCW9XzXHBd3bdOzeYwe
44cUn3Y1z5xJtLKPPWZMYlyJ9qCWupZE5Vsg3g==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pKyysRDfDRq2uWj2DY9SyBumhMt32UbCuydjdoIBXHnCxoa9K8W0tPBijFY7TxWwxjCKsAj+kEvj
VtrLvHtrCvuITfo+5kyizBYnGecsUq76gq1jiH7ibthaaoTsSZdz/yX2qho4AswTYeBrNIFRKKMe
ytaGu4E3+UdZJ5AmlC2hS9L3lKp0rYpW7/3ga79U0NGN3PYu4ctIQY/piPLQqm3mLXgYEwlLSYSH
bF6Qetk8JiduocsQ5wCC6ymA1HmnZVZWWMFWqekwyt6poHD5G1+Kc09rJ1xRCleye9m4OKUo6xJs
EyY5+aaPBaQftq1EZopQmHLf2tg/+2D1daktcg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
8buQiSTKBblNwnPy6YQcUgphFPd94u3s4FHr3L/jtuf3AQJcIKnjxtS3sBbilLNA8tL9HRwQaGVu
s0AB/zsIBd0V9zUap1ZwFYd+bUfEo42YsyEs6Jn0B4ejtgJsE0sWwqo5VqeDB9JuQehzR+q1mh1d
FpZsOnVdoC5W85A28cZgUgwdXO2QQ6DLCY1YRikBI1+wZVCDk/fVSVZrJqIId/xmUeskxOiWVEs3
V2/P9PPcYbboZlSQYp41HyNEMuHk9K6M+MyGwA0qxSByIIq61kNMdSMd4jw+Pi0mBPvpsnpGA8Fc
2evqQ36hzCZDiyuZMdTjN3OUXLi7hPmGnn2oF67w1HoJFVZfEpXW/LQ4k9/gr6fBrTn3vs0HGThC
9ZWJJH/cXxXhECocdWvt/y6AQtWNsWcclTbaC1pUIVi9gAOVnMRnZbVF/teH7X1IQtOpm2bSZHLf
vbighrVefNXZDuYNTPWRV7OpuSMhc12+InXnXNud7C1KdyxRvPvMShRY4k59lg4W+Qytv7W+Qbmh
lngBfLYNOvnZBvpyPTYOgaQ4SPqAO00PB0n3TXhdg0Ezhva0nACtFYuDeY2vl5LrepssLKtmqG6F
YYTwl66EqWIQrtOBL/w2/LMfYlEBcoI0bW+wWOoEdJo+o2MZibw/ynXOptzbLAJgZr8TFLKHodKu
uXyGEOI5L5nfVlFD65vlJMCJ1b/pqev+jdNoJHfWyjspPABlNLHKCJx5lzUtLF38Iop5KJgVK+F/
Xa1GpqIulgb4iMHZkRRhVe7ba6oO5EiKIg/Re7i3vCoq4whxWrxrtU6gtmMRJysZELXiLtkkNclK
JZlSQFviURui/QOJ46gQUo+wsm4RLQJwTuoZ8J5NGcKMemExPQGeFHzYOUVghEYDWRDRXrNBQWFs
Qi1mSlL+LUcHGhTpV9NF4wdS97PMe8Cvb712zbZbMdjFWc5PfYAPxvnHlQR6KlIry7IGl85C58lP
abFV9bLmApq/Eg5hNJzbZFSCeLC7ylDe3y3jx6jIUCWcc4rAyQWGqMp8mmCbBmR+2plCQpWo5PF7
1tOb0pggoWvh7LmWSCAj80iYJsqf57sF5chPmKBy7PdGd7bxySTRxSNUhjxA9BX9T/+oyxCcXy3p
9Ub5B17x2HNLOZZHn4xLSTp6iLu8yZCUosI7lW1eF52h78dir3ekiOCJ6jHHMVH3proTaxL5oo+g
V1719s3fPaFhBXVV40VVsJNwujKyghmCGKzvPtXI3Zz0Xq3HmnFPUbtK+XK9DEImswkI/aR2YCLy
NugOaWE5MEBqgaupX4ZTUIqzy3NAfq0w9/0dlFZy2ODcQcAg0yCrp0GAa0xBeWTvydp8B+utaDT+
zsPCRbfbRplAxI3h9TmjC59Z0uUdOEcYaa1nru643DxGV7EGqAFlMpLP6vMkllSBapLT1zvGIf2l
Z1Yt0vCcbHjvQRFNSRghc2ogPq9L8Ut9P8sDF4eQmWEhzY/faUvDwuEFVYPfHXP8+n/j2uOvDdHC
Uhsg/JbWbUflkqrYUV9pJ/e0of0ncWKe3+1OVwO0KE6SyPNGT1btxUwFqKcb5o8O8b14iZczcaCV
10ee+71Xp8OGqjgv401kbPLQLbCeWQhey5IIuse1hkmJ6KmkOMAVPy0WSOe/mKG/jdZMvo5NyBhO
4F+WbJGABmc3YJlB35r8PiyMyLX55o8c21lqeZRbpQuLilvJnU/kxaYYueji3aK3Ek9EPhYcBvBu
oW2nAZVLWgu0G5vTGdemebqAMWp1EA9BzDg83w9dEEzEpg7GaGVu3451XsUWnqetksz8hAdkjYT0
NF4F48HOEkK64jbSwyhWYoNpyxYtwHCuo2Bl4oaZUMac8Oqnn+GbvWBlnTkwL4+Jb8DuXLyjcrvQ
HWCwT+27gxM5gH2DBi84HDroOi6Wtl8TVk8NmM3A7uZDRD6m0eO9ms4bY2dPshM4Q8L0TIHDLaHX
BXoiIvku+MyNyrFb1VBKutXIyqktfllt1ZQn9Ke5laJ4YHNT31oPk5VGjXt+R/TmHqoXyLjcKy1I
G1bV2hwdv8I4OUrW8ZccH5raL+CuTznWyAx+IrGi3UWERK0Q+IVUoKyfcNWJ2V3jwFHnqaHpqjsx
rAferNvL7yYvTjuZkgAGu0svzqHUUEKn8lNCWCHSvelhrKCamI7COgUW0O6B1aZ/R4pgjbHuUtRF
c++sAhFwdmTa9U0PfixX8xu7LruKsVGrJngeJqzGC+seg4d2ZEiarMp18amZzaKnhNDbMVC9XhSf
Tca2eAPd/O1+zD1/ZSRmMRlAyUl/Ffux7vFiwCYgciQf1OXru9nlVw7edyp5bmTBAf8OgPybjUIE
cPKSy0Co7KPRsulvcnLz18VXl6UCxNQids885ElXDmV0MIyD4ph9oytkBRjzPHmLULVf5eC9VP7X
vsUD1P3xB8hpQV7rJpWfbQDdGNFkHIpDJyH0bRBghLKs8y6T5k6V8CfYK73E19PNezwAi7Gpeln4
rjn4CVnNq/JaVy0YkqaipUUHxjVnsQt9T/u4eD57+LXPvC9GNM+g7q4AyXLhLj45aJfK3zSysHGx
/fOG3ppronu1Lu8Kz6NsO44S6f9Ed1XdUiMKObN+vPlPyiPUH8CbkjnwbjqJ+P94MDcEKAH28OT+
ebr2lXkVvYBWZei9PSrOZEhVXk0osM4mNGH6qfeS0qY2fNHd3FC2hvzEFOYu5RenXQRQU4n4hE5x
r8KbIsgNvI5b/kGWOybCQcrbO8RUHQtQ5iBIQe7Ul8gHPnXTipsZ99wu7CMBluvVvbFvGs3Ibs3p
LZIORD9uhK/zylLTVc7zsgvCZRZy0hImClylQNASRUTA/WeL6jxoSGWWasujTBNp9ssjVtG7pks3
esG800bk3m1RyPwmzev0kc0SXGVfN6EvN0zCGBsaaFX8agTQcqE+DHrnK2+hYvwZrtXclzYUO0F+
e9tWcdPZ7mPUl/1ucEbs1HjztpVSdi5fVZRV72uifp58lp94+fWEz1k7VkUUuZPEJkwu7JHJ8rDp
KUn7eTmAxd7WIMulLdrtDqMKWydLMGcA5NTkecHRjbIZuymbnwvHmBYjUMBXcgRIKzFVzWwY6UcT
Y71cJk98mHIoVeidAbTKE5Uz5K3C3YhfudQmUR9J3OFYOfBh4CzFs/zvbLG0LNZNZI13Kv5it9wg
hotBPHL8vhBY7UZYIvd0tiKzannkDVFB1dsAmoqenVmBLj2+pZ0mCFp1NMTap1CJNnkEjAePeR0f
S50DjKD+monufkK2CO//6idYAUXI8J2ksb7p++F0h0H0nZNATs5WAOk4T9vqQ930NypKPkYNwGEa
clvHLUYQFe+epNOxabFsZUj27PSIHCmBtLVAq0Ux/ib3kM0xh78eOFwNI0h57fgEdwIu5khN3HFJ
RvWArHgjpbq6fDYkDAumwFJ0BigVD1uAtsf/Y+7oIFYR9zcy8M7htnoV/mE7ZjTwGnF5v5agyiX+
PmPm756CEyLQeMWnat+8MrPvb6NPmCu80L0C7HXaLFzCsJkkSt73JhrAbAr1tn5JYWKY7IWg3gui
fbidfaDB7E6j5H1BchVBILynWmxGeffdjQm1MwSOWGYZHLTlGDHeQxY3nvDYKOnZzj0DRw+IHgxD
CisOaTPrvK7B8sN+X7vhAuMjYpfKok9DFKS8mGkBffHJyejaaJbzDe0Y9Lu3lU9/vBtCA/+ayYNG
DvUqgkRh21+g6g46eDDE4SMJThqCVbqsYEljfIKKkzD1AopH2+vV/o+A7H6/BxmTPADK9L9FdFmP
gi6uU1YlHt8dRYYLvAi/SlnSQxu3mw+JwYD3kyY4pgnTVaYLnNV1+GST/CyDaRm60p88FQNRwDIY
6f80Hki7DA3TqijpftTqsncJpJSk5sBl5NOINlbRmlsINcCWrN8HPcrG/Se77PpMXnLgjJ+tXBY1
WMRfEOPEpUDV74Jac1GzTv6NGsiZMw4r5SfEY+FaM3s4DiHZR2sn0DkD3r5SYkCGkO2MP67r7lSq
i3m/WoLb7zURxFysqTj7sHNATCN6sCoifdjUNN8MAt7Qrowx6rftzQNb9Pm4i99iByorIvDmX63m
DyIkfymjCbYR98vjJCSO4MYhZpM0gAGXvQd316BgfrEj59XV8Oy7DwuY2RB7exJuqnm/SkNWnFvx
yoaA0112K8jw0RQAHQ4sklCZ/Sknqw5xXJDHSUVEg2qYkvBe7mIjVKLAFEL51wx8gejRzMf4aMf/
IHHA8RJ8JofIU/mJPTjtDSWq2OJxex0+6len8stWEjwATNtf0ZTIukqQR/mj+RAb4gYmJtuWJW6U
sOek0JEWXxPGTtY6lQ7WqK/3mbz9aE861GL8sM+Npi3L07LQzklzd4Q12j/Pmr3xspLDGqWXI3ry
wwJprewCXa1w3uR7vroc4iLdweEks9LnHmmX2TmX6SkM5vJMCUcjHRxyX2mrWSLkQE/wqhSTTM8H
A6+MDVQe/W6pdEc40N8PUwmwReIK1+71rOeELO9wqBQ9U7iogRqMcsYgR4UjhJAvnJTYUGLzCChb
jXhjYwR0j3xMkmzN2reM3nMneMoCdgr/rIXcPQSqIwu4Qlwg6hKc0cELJ1z/eDghRzLeqVVi6f4v
WXjjAhhwCLxBh+NbnV65icrmu+oQFd1sUcwBY27g4Sub9c3DMep8NYzVkGv3mwDKxaLzblLqzO72
trXVa4yx9GnlEHCPXzuX+seyZb1VwsyZ5R9REyhsFv+0lXhrwoVWjCls2QgsW6CfhAgvg/Z5N2p0
fQ79Oa5pipNEW6s4EnTWxea03R6rHrfKIO1aBDC8otrYOUabD+kk60y5aa8HrEbL7642Ka7uZpBi
GDNZkJEU0bzufq1xPUxAKQ+KM/Lda09/TkjgVUz4zr9n3Tfb1PYQfpNKhKpuW9dHLZv4MoZc+Aky
LB/sQi43YuE9lJFm/6c+BTY2RSJEOe0TNVKK+Hkcg99LNNYPcxUPy9IZnWqkFqxpgNQ68P1I1xOt
JNIZCUwOxx5oC5fifcPj9YqhpyI/7M9+cCVgVz4oYGGS86JOj5YoWc+AYjelL1JAWd95TruRMtdZ
v26iD265E++vr3e5D6kM2lcijLJbF2A7opZvsQ6wHWn8ZKOLUZ+3EU20SLRF27DvBdVNag3cK9WK
mH685onbDPFsFuuCe24XAO1W3LQqEfS5MQtW4AI9osSyD7fROc0bXmrQrfyHfSWXG0UVzN2kl7bq
Van/Ny2bZaJraV32oFhyuSQm1l66yrgQP/pxhbH8GbITwMx10gCyWQ9R4d52RlvVopw0LVwHdG4j
Entip7xv1EdbTjrlkKEAYFRtN7vt0LoIUF2esTa02d6x8Hijsgxw8wyFO9Jup4PppuVDhkrflkJ8
SrrG/wD5KP0QYX2bcRZEpd3sk+stWtc8+XsHPv8cQ5/pYGNLnzNmIDiVuMGlCbMki9MeAJaoqGWs
rdArsgtudrm8znsXNuyiyNvoYf7PZqQC/bSgy/qFs/pGGKriptaNB3f3QD6ftutUnUutJLiYvMSS
gn2lI9EHAmaaC2q24FyoQ1idoQbHD/IRLbCZmrC7HfO2ofm2QC5pl9pKrsFM9TjQW1ZAW/954Lkh
ZmSR+9F4XH4Qzazo9Uv+1IOKBisctH7NaBtJjCMB5Vmbw+b+0V0aJNdXIlm3dhpNo1IcPC49BhdA
PuwR7UVNFyc0jxERRb9wC90AP+tsubcZr+TtYeJBNyxY7jnfVlnviKP8Ww6CHWy3+pA2vTTNNGe3
ZJGPe89QayymhhjTSbNDNzipOK7mdBszhsYotsmNVr2jbI7zCzsSsXQFWoGCn8/gsZsYcJp+7Y8M
/34xjm/9wnNQVNyyaUv5Id18maWizEYZ811ffthOq3n5ZNbYKb4lErFLOfro2uPZN2dru2pZ9UqE
bz8+e/fhaOdcV0qqm1aqMINMAdi5n9ZPwU615UpYZRKKPPWgebcz1YRnGRPrwSYR4s4K/VhLiD4I
JDoQw1SA6R0UlmORnifeqhKwQlBR74SL7YolPJBfqwzwv/QO9b29mPZ6VnOpWHud7gy/B5GwWmq7
izn95Q455H+ol3C2nGs9Q71Y+fmP/katZ9/xH402QZyw1ByHqBkuJ0N3Id11uAdpLHT7k2gxj6Hd
EOHggGuL2ztkwKenP59/gEMfWjKeb9pwfe0zOXj3lfIHMDcX/dSlZov/ZQNaAvyWN/fKqOaOiCLF
H0S8FwaiLwWO6U/3R7AfVFAkPlXpknwlhkdSS2+sG5l8MPVFylcUUEOjyPhF+Pw6nvJIUU3Iegit
15bfm9M2ROYhk/cW1XJaSPgUa6IxdzUDlNkFZCGMfs2p1/HMtf6x89rmUTZOHtocdN0Skc5ukolN
mncyjLI191Hrmsu+3jgLBNmFEToC5Xh5qxuPVoESlXBzwVI4tLiX84ove3PgNmHwAdCiutUaOw6K
heL2W3VZsv9rx/xTb0+/88dQqT0BZuY4wG7vP3UNX6T1q/lPx6aorQFQgRNFKmaJqBFZMWUvMCzN
0aUshe0fC9ldq7qRoQqkL98gdaCzZecGh+8UslfyoWQPVS72zMoabobU+2WVn1bCDAWl3CppVAyu
39en7TTts2+Mb4AX9hVPHZp2KN7Ahhj3TwsFYpA4d/urwanvYFJWzYsw5qYsiUwQplR+fhMQmc5s
QTsZs582Wf237ftv7PW1K7SbO+aFHgHGoe8mHFJdzv7nTJHvgBxAQjXfCrwnfudXsBIaDCXC2rew
hO/mKc6l+3uQ2IUCckPO8X4lB5gXoNAWeg0Qq00fxGnKs6EHqE4KdVvJPKoBDGdGVzKU8bZBjaQW
ouDs0/uu0AnfVHZmdfGGeIpVKbFLYaI9pxklHdkHOr24H4KMltO0ULenTg6ITnRvxXObwm8y1Gvc
2ijowKgBb3PZ9BiFG391Tn30js3VpvaZ4SR6e6G68G1PHpgwbF0WIuRBV65YlYQ4rmEbzj5wh/W8
VgB/DcyESvl5Bfn+s3ojfrIB6soYxR5pUfLh5GUyXTEXNHCt8JMc5POkRt1kZYKHKQaZDJqX5Xg9
bVNnpfO2Q5XmV2paobVJy5HfnYRLed7aDlnjZz82fgztv8YomodDvj6z+Js2jY0csUNxcbytA5/2
M6sxLWdqyv3nwX//5nsYQsIx3weZLBxxZfLL0Bv/jGIEd3M7FKe+GNuvVrMgDtU5OyfpMFEc0bno
ff8ITMN+d11JpYxpmSCinyA781aexM9Zg6IwYcE0e1P1nCWzncmlWTpF7AXnN4RAtVHk0H/pvT4l
2FlS4BVyA53syt5Emf/ss20U5/KTnbMc2Ow7WimoFxe6+V++eMQiyD3E7Favqi1OYtw5xetieYL5
aBcZ+1vEONDA9mJcyJnzXs7jH6kY+cO8B9gk94QuyRKiNT1nu2ev3SfXk5Ib1mtD+9zKyFX0VM5L
zGi93yc5Ij7KMhBXM5qfBSR7yBNtw9tO4ncZPcPjOkjpGsLUmeoJDpQ8wp0C+FHua2EwRnN/oQNh
fd12E6qAgc24SrTuSQBM88zjiw+wFD6TIXqzdcdgSyNqD7uxSFbFqgbTUeV0x1J2l2ZSHUYgpIpr
ybBB6aIpRkqwGIk9+Voh7GAUEGZ876mXkqtyqLlg6blNKCru6BQKJ7VNHYdFcJsCTlICdsH0T4Y9
w6SRdQwclpL3b0SpOxfumi+4RNeb/rRLuC54ZX4er/+t+TzT2Fn7wcLflGvLOX/SP5Q0hmzEoKum
0z6+TLU2OD3DTceaw6ux8ayyH/g97yz5TJrP3TaVaO+3basnFyUX35DxwHl2DqcFc+okmy9fcL95
e8gutesJfnTq+xo+gSyqJoSkxdBXvSRZdY+vu/gZgvAmnYrtoEPBIYv6gctgx6YA9g6K5uIgIPI3
BdpBWL/wM6K2xbOmpkkqSF6SMxNGVvvS9CBMS6rJkFQENUnC1cnS9JEU/77kG6M7S4oFvUeNky0W
7Q++gpVBHqMJoHxft7k/34RGbI7vt0ajj3dWfBZPzQTAF3MeJRewVumYTKom67LpqPNokWv+deyj
z2CM+ogI3X8epGs3qTs+ez1Z6cSijHi0h4WbPYh8ZjlzcedZVd+EjbfFUvfkauz5jG2cSRBsAPDA
nXedGd4sAKK3lZd40qZ/Uj98epWM9Sh8nLr4UVk91idv714TseuQfm2lCbCopIUm6Dld9UyajzMP
5rbxohwqpCIcVrFU4sIt9ecy2u+fT9/zFsUF62BsdE7MuXPoup6I+Lz0ATFOIk8eSLl16qFq+Gc6
er4IxOg2wuncro0IvmccVrb+0iaprlIqUtzOucoTy6XjrZPwyOqX+F3iuA26ejPI/JgyQoIWQvZG
nM9N/XgsjkTyCRdeBY/IoVIEL6cIjxemHKZmpywVIK2XrrqJjezNN2ShzGxViK1SbAU15MCRuVeJ
7gPJcLTzXn+rS5aRtAAyHfXYjU7BvFHvIi0Obc7eDtzV5K9ksYJHh1udi2V8NOemR/tdd6eHMtKQ
5lstRS+KL4M2mDyNyL+DhOe5eJnM4CUoe/ZUxyz9ZMqsxRDaF0mGUXFxCxbQcctgxN3JqRPiYLz0
rvBi4ZNmSBujPDQJJTQe3dn18EaZdkKXIqi5LG0t4pqmLLL2vNDLz+WnQEHjrjXrSUEMdfHOlPwZ
5lnPDuRae8+V5lg8ztEAtvmAVRSRu2y5qxcCOHrtwh6QXiGf8WY+Q4kMX+8zhBQINGJ2NxdDWt5T
pNBlqSwF9oaxROv5H4KBsSYLiVgXcDKVaGdDEcmsuhtetHHgRAefPO7CMbmYYOgbvfOEcKuZ1ACS
Lb29EdW9qwck0mnZyNj2zPGobQqETftoOsIeSDNMo3UixWg7S4eLY9K51wnZdtM87yabAV9/xTJP
/JXJGg3c9tNarljB8K2J+EqysrYwYfmXMaSNxQ32pmgk5lu6UocYrqI0JpgSrxcK6R3zqqPYCiW3
sddrBqEGiwVICzi8+TMTZBbvbtc5zLcyGU1p8gxMSLNiDr5S/vZc9gkQwZVpzOeuQ6zy+1uZhDLv
Fu2ujFL4nZISstQ1wxeCIs4MihFkgQV6xb+sn8CtkNrN/B68E3l+m0ppZ/Kbg0rnLZBqkPXWku6p
7VOghBK9mkvfbhcA/3JllOyeF49bEshXlzQSpD8Acr1xtx16z3uNiRkc+czLzkkypyGS40Nv+1rZ
GBpLidzHRbRuht9eIkW/GqKlaHMVUBOZ/KDM50Se+Hez1utFIDliD1f1ASvevIJMTSKOEnfJHaWp
dky7BJ+3HfMfXblY6gMpoIfz5+75PniTrbpvrTvKlgel3ZUBLq00Eafiik3CkatY6sLm/7iCg/+W
5Y3ySkcV2qfRGnSmrhewE1Cl1PxFK5TKi2Inqi9WOzoD9HgFCE8vKpn+74rTrEIr7CpY0VRGN4/0
vmAbmQJxnX/sqL1+sibtFvnV5Y0VkkphEQVaWn9oHN3l4QQTPs1aR4HgvxvxYqpRrMqS6DFTZrr6
5XG9p4kTjh03fAfOiEyGHRRUs9LL0cRd8XzAJ9DvhPRSPSIbMRmYmcZTPZ+BIOA3sWSgLKTzw59d
PuDYzwAccUKk38+hToWHEIAmKC13dSGU1yCAJhug+72gI4NzXDz3Y/YtRnSANMUAhFTpDXsdij1u
424GRM/5IEYpcubVnqA2enP4FUTey4DlAPmpGavoT+PN2RYBziVWSxOf7d3+96Gw5KJqH8+toGfY
gZuYBCmwGxLo+JpO48b1AO368UXPmkYKdqHlPjxIYYPO9L6QjZdUa2vPgWx8RUQt+FTibwGRraX1
Y4aP/wV1XAqmx+ZbCZGIQIMntd2VRAbqQ7cPcw8BWuw9C7BCIjBwq3ksecdfWFgyiQ7w9ZKs73Lb
nGuoZQr/lIOB7JcYW4x69DLxQCeh7ONDVQvL6adDNquGw969wyozcPdc6Mr6OkwKhSv+7WEnhvUv
K4vZ8QOZNElMkXJ/z1SE2mS/uR2Fd0Zaldzd2rYLyRwi7OfTagc5fT6H9+kkNf/hNuiu0AiHjvO1
LHiatupgdL4VnKFWM388RzCUfIG1jNWaYNcRBlKQ74MTPu9rfJpljIwysckNTz6iN9rgfkoqaQz3
B8dyano+6cjiXd4GG2S8lZcDjdSpSgNxAXF49HybBvGNT27tlu9fasnM7fj/NQARmhKCkaQ7sHmk
l4bWISlliFPY4Xd70aS9A449Kn21gh0AuHEr10ZMG+qSQfti5IJ/4/CT/ELDc2QYoPYuPkLitsOJ
kLetw1W5rfV0UqU/qyzk8S8uiFkgSJi8PzcsDV/2UOhbnJob5YIXxM3ZB2c3nXfDskyoTI6mQpvx
oCuD9cD2INxG8VByB9Ew/QNH1ioLS/7jdtzomEuenG884XE7CGIUHYixoCrttwXYjkIhCxTjFZo5
e6eGI1wQoaBkbc7hnQxrXCdWim1n9xKeXafTsIHK9tbnyD85epsA7e4k536qngiDHNTWbWoJxgD1
1sX/2d83/C46cRC6FdVi2FlNIGa2A+npULhkOg6nlBRDQNddlEzvGOCFga9vLAbwcuzhT8dtdGBY
EOUt9D5kT6xHi6UwvWl/gJ2KDOasFSY+KITFvUJG2KijCEmxT5sqvFtNeWMC1tCj+hapinkkeX3j
sDtmQHIKhR2ki7Ns2gFcvG/6unoc00Zi6dqVC8Uz9OjLs1MdxsTi8n/hChyZWY5k9GCO1s5wbLxD
aT6P19kQyCGvOVuSYCIK9fwyb2823vCwhQSZWWB/PF8qjQJBciInQX+mt3QgxtaZ6f91aLMOa51F
83I5vXy9+XSsHXtxI8tHjXWH4vG9Mr+qtbxv56X8B8grEPGWlsS62bxflnJBCJQN14wWfSGqkl5V
o73oB6oSglWL/zzPFcvRZvbg1lHymJM9rJmZEKfqub2otaq6cS6cJ54GDq1E+4RzsUcQyrPKG/gx
jVRUpHg2dEFsobObI4IJtdf/23JoSBmMoUVR1XtQ6E/4JP8FQX5DnkZUexwdm5SoLOzV7YvmD8qM
JJm0h2oi61EJ9TkUpSReg3//pDl0eK5KzHcaI08ym2RlClrCG5DKh5qiiH6p0u3m3LmBdcRmJf4v
DPVWTiSMWv/iEnAGL4eWeT1Htr8ZNy2iSkHXOyKm+0FYeAsVWFRKSfwdtFOLIwThcY1tEqFbCRkR
2waLwkntSPL3cDTlsR2VxLLL1UDgf0z2twv+ao6zN9GXkeFFIIW+jI5vQmiKZO/PgMFerrErDkkF
szYD+v24VnWXmKzeN9YO6rp8z/i95wQjifA1tIAqiNUu1CETzadxlz+XKI5+ct0nVgfRqbzniZhu
g21uXW8tjyZR2hclfcdbqo3HbLn0nXGccd4YBM+Sgj200HnMvuKHZ0op5m5ZXULiaLz/oBAGwXZj
kbYYqPu6MzchQie65h0oe4uR6J7HDuDaVcmgftE2AV0KvswwTXkr8D38ti2tCRRIVQwNcaQ8Oy3O
fJu0mGEpHC1dM4TNGXeCiUNbuzFFDeEH1rrYv6gBzkwQ+sduIItFp29SbZjQFZH3sZzu4arGg1wG
pT1tYzCniomsSGCtZeTKJJsbbzKzZbdAlbyiheg92UacHCZd1VcTvd7CIL1b3SR/DjEktQ+VUFs1
l2CEMns3hOzFMhI/LS08B37fm+8JlDlIrB/6vuJU6IJlXXMpgxxBP4iScMCdaHY0R7rv6QP9Ywpq
JVqBQHJN/+BmgSyEeITw9amVgXdUY7jUt91A6dL2uKSLrUaf2BX1rNoCM+Ap+GEhAMEl9POJlQrF
JuT9r/E/B4jgIOG+/bXw1CUrAdC6UCGPOYLKgsAwnV55lOQNEqX0gg9VnGqMbSO4oI3YLJzazvcA
2kP+Mo3vMjfYQ7r3gT1NcfZ0cGPkxiBRZIGTHV0UplzuRKyJEnAd2CQjNoFzHm5Ekh37PXkc/MWK
KRFOppNbDK9uGkDPXwvPaMmwLFuXUapkoYiBeWS7u+hc65dA81a8b52VSBfmLyTsC1L9W7uCBJDg
wSzrdGg0elfIu8syPyYSa62Z+F7MrvnlLWSf370QP+o+XzWGQzGOX/FfcJvdh6gyOPhsULIikRoE
qdrukq+2Dugx+h4dSX4JEvf2txji37Hm4v/pbesRTKsY8pDTTyGYgWV7aoJSG7fPLADOTjk3Gsyf
2NGNpi52xKKzGVZ2waP8UKYAdwYX240Wxkfu1PpXFDuFAjoihOk+Qk9hqagSQMe75MReRH4stu3H
COj34sz1fFfo+Rzogj5shXXPdft4F5X4D2fs58fPrJ0evTuTaZiUkXN4DHGxSVQULWV0yt80Z82l
sGbGWCrxiayp0jeyzgXu87l15HE+8haOXnpx/7mnzjRhYMxr5xa8ymZj2aYz2FquHDta7GuTCEhD
wVY810wYwXz9Qode/STmjP/nBWjRYuuSXpbJ4LMYm1kdDPpznmzwiJa5KEOATpfpmwUt6O/XgJbQ
YcSu2FUe4D30Wm3/vRCtiuuLUTA3VI7riqms7z0xzBmdTxwDMnO0Hr89SMVaO6poDUfo5B8nvw/w
slGHz2fc08crXnEbauAFYylu+Fyp10m5ygVj9xbWbXK48AdGbkbTRVQFi9CP0rIQyWC1PU5hsSDO
1fXkCS30Z5K1i3cuSYKXPpHLgdQ57U1X6vlGxvfJkG1PItK6C2fEG0bxN91Ox/tvMPIfE+uJDr2G
dRIaxgjNyn5M6yhCpNBEtPxjYJsCNVInHwVd/9zO9/S5S8R2+XtrqRVDXAswLYNwfOy5ua9AcIVI
K8HzvJvQy4Y+XEVl4/Jmt/NMgKM1f29F3UNzOZURibpo+O2cilIsGXnvyi0ZPiVXk6nQZV458P2A
TJ4DIfZ3Ow2yHsWHVrcf+DX1ODGJU+jCOQXMF+nhpvVGu0POu+Tqm3C8qC7MhmwOy8R/2SHc+vb1
RxMEdKfYYewIJFQaU3Lqtdg74U9Kgb/m8ciJ598Z30dqiAAK8YHk1XI5cUgtnKEZOo+QYohYB3vw
oiZc69B+T0d9fCevGXxAyj+rcliUtMXEMk0M/+J7aFHrblh4QsdFd0ooGmNAPjoGBo3d4hRuyU87
g1cepNG5uPXBtg+JkdXiPsTCFZpwjfeaeIevnfHAu7npOXdaEFylgSlQAzVX08k+GBtCzaLlDqXZ
Yu4eu7VPeS1ItnOjGr3Gc0XPwpM9CFdFUkJEu2DW/zKc5CXyCr8KhbqVF72H75r06aMTjR1iHCy0
DaINxNMXCjra1zLeui77GgFSwrX1x/77Qf5OPIAaBCMbTleo4rCezrOnY06BrggyIkQS3MDvAiwh
jFO/tAIYimnOtbd7+WfxHmj/2B5YnQXjd4QoWiU+MI68R+5mK9xKEy99V2b6pBpjMzvQ9fs3hTzg
qN4MyTiSwJtK99Vw+yRjJhA8OdqmyL07OI3qklBKE6VUq3DXiEkbcQv53sRbLP4p8w0E2pV6f7xz
jlmVyoiQtg8v/sTuj5HOTu9VCIPuNOmqLYBGZ/vT3Rpi8aWK1Q03+eVgmrIUdNOhO9Rbxs0Fsu7L
XMIhhzjSFIQZeaMpexa9NWvCrTukLa3nXikxRIgwwfOKE+acXcME4uJC5VArtdTqbLtpuXw3JJRO
WWdlJA1cFgwD4M9W0GzG3sHgS33Ulq+qYX5GRiD3pN63u+OJLkDWEKwJFfIig4rMZ/dl0J2PynIG
7vV84wDRyx5QMXD4HJ0f2qcCLgVFJNU36Af2k01utgmRA/0PyCj6IpSn735kt9zrWh/xDKH8xecJ
AHj6HM6vS19gKzWi6lhoukY5j/IIAF64zh7pBaAbLjAWNnRljRz83TRJdk7Ox19qZtVgz25WWAAc
Z3pHM0IyGtvdWPPd9WtZ8XcSZ7vog26JYqM9RWFE7pgWn3/7FUeOtV3QwHlYDIThJuh/z2j5SFAz
Pz80HCapqZn21AIs6mSnrrKGKQHRV4UX8JJ3No8v5vwacIGftJ4/TxHEwE8TYdoigIIVnum+bLdV
Z53L2JhnOVaiaDs7OoJuzTv0ZGFdgCPHW81GHGIh6f/mkjkiLF2jOgFHvD9XQ4BH7hgk/Zp/IUZi
RxsxycoWDl44pm+aB72tGrB9PCch5U8GaFhLetO041wRcQ+y3neHQ5bAkLiP6yscEidsoXbv3eEW
rk2vjAhzu9DlCYis/mDdxT2zLAz5gYpQoY7NxLnDEN/uGNpt+blTswHSMczjb34IN+XZOL2atUsY
h+3OvFkLKmkTh8GdAVuTOLcCvsCnZATyzJ211VtMpqzLxUvNGrR2DZQTRTSnKCu2Nu/gL+mjkgol
x2JtmeVwALdwY9kQcHAK/u333ujcAVyzz4uedh5qbbwXLegcPW6yBJT69GcdB6TgTlIco1AU5OyD
i/p37m+3OaKZUTVlwGYExmxPdLWEqW+e2e996awJFyVZbOYPtFgQ49hbMBXMQUlGuGjESXXsRLTc
IkihtIOwOiTc62hUKzU2Z/9/EIHmE59oV3LiaWwpH5UEkUIrpyAK1da+q81HHMU46A4faf7/QR5V
5eDNdkGMlZLu3/tbLxQo64CoTn9zu3OKZmvK7Nl5qkB25cd4f8s4IzyuX8ytSqFnK/zhixZvcF/E
cmn+Wdzc8EPeBBTN7ucHaOPCAMNyfjd08QutKbsrwnNvWmG4zpDADT5i5m4FnLMGVYjA3qEWwbVK
TK/wrhLQL0MkkWdx7Zwxjm+C+nr+3TMA1fYpKYURXErfvt90KiTUj3D0CctclyJ7M0R1ylSia+7y
UtTxTHHEDcykgWerBGHCFOYda4zqCyUm7kQ3Q91vydZG4Ccpe3jh7bLjjEMXCxS1/JxlcLQXTN9d
IyZcdk8aBiYXUGMnRAXQrrxh0+7p8V9Rq8gXe0oV1uf59oViAq8iVNyBeOI/PqMc9nChfVggpDgR
jHXj/QpZNrDLuHnZFnqGDevkJ7K8I6mF7wIxKuFuM58tK5KqXOHojJSu4NvRmrB8Uok+QHKVskZK
skMMmn/m2SA2jaJtJMf4lizey48VzdmMOQMwp+pkWXDviiDJqyX3tHBpUsj+GhSLMvpGs4ZC7HtK
6jschFtLNBr06E/8nxlKLmjZCbTt+7XtJpcLPXU349mvVp1HZqSYYuApu7itOHy3lDV3MjdlybE5
IWS4XvhUjxmdqlRP7Q/PMzVvkKvFIlNpkQbRkHKaqCS/1bFwpiotpJgnwbRjDPQ6PUle7P2OTAEu
WqVnRLt+sFaDFiLLg1kdNITNM/Gla71h6yn2M9ZCbl20dfv/V+9qldUBUQUWYDuzkBl3GuMnsBsw
BI9+YQNGP8sXonhTDl1SxJPlk6dIkud3oPEmidmu+DtCQehnE+vnYBtfHY53BkOT46aKd9F7GOiw
1rjikoMop8h5JQFkGoqKqsc7rDa7FB77W6n/z0xwX6OMgseYAefS+BI+heAjwsnYQjUyB/NfW2pv
l9/09zioP286xjTdLpQKuOKnZ9ErRku9LnvB2aBrUjXIxva91DOWhezqn4A5SUzMtJIVjdKSbJHo
87Q+lluatcq/GD1rqyq4qNgWoUF8Fd94l8OMmtq/r65tWt7xRjHhPyb3Qv3N62QpTJokWguXgl6a
UYKSKIN0pPK9fNCL37lvUtsOLjSHd4Gm2nXtE5IW7m5DRO0OSaVoLEGxISywoKpNLdGKYFoVeGHx
lhHOOQFNwb7mZvczBWIZdG/eMQ5gr4eYyfYnsXdgC6o6pdZYvSHRu2lpo3IDXXFrgyNAVWJDXjTq
16RExctqD99YRe8GTUVqFKtcexpcJgJQJcv0okl4tI8OBEpqB/r545f7fiudlKfSU9vFYCiw1Kdv
i434eXq4JMvVEi5GHWbNfZgn7OCxlpELrWHmnq05vRzSatW3x3G9a+9REB7WP90xLvPosAJmuPSh
zdzwYMuNvaaM+WM0RvXMunEtOjUAJ5xkEfFxT0uEls8zfH9G3a77n74XhYt0KgCqF8g9Mk3NG8s7
1ruJBa9WgcLHfkeiYYvJNumqhVrpLH289GFNqwbipIhqjNtwn7yrdKqQqioBzRDMk6cVsiZYPFju
x7/AAIXPx505PCLAvraabzC53Ar4VNPhtQJPwWvoQGX1uFTYWEqrwk4ftBE0vQ2TzOeVc3t+uJV4
ZYghemLEtx78Y3kP3lx5pjMvZ3ft76FX5HU71MltM45bKr9GOBPZdlK+PqlYGGJpjEsAtF7RJq0o
udnESKlE80Xe/sS97/ZltpnaXSNA025+z9uJhHCsfqHFqu9WH/1+o4V0MO0LAeGlZDymjJ9AT+VR
eMNW9x8uJJS0G9aW70fOC6AU7Ou1peOUK4DnniYO3vZ4ueXKo5HOSQUGu8jNWWGBIW1KwYtz4nxb
Lw5mUQ4iyYnxpDSVbtSs3YJoYRkTfDLW1LzheHYdPZSKBbbpbilRcN6Mi98EV61MnMR0XNhLPAM2
5fhmDfLEjywLRow2Q940CGfT/GYZbJc4Y91XVTyB68/N4/sHfFM6SGEB/UajCYMq+T3IFa9sPGTE
cLd27impEv4OHW6INsL0Neyz35eRHJgSwal+zQveFOgGfIwsYIfDtM5nFgjeE3pgK8RoPI313e1N
49tmOg170VMOxlM8mZ/bd84KEsWh3n2VSsW6Gk/s6B3/vTA1KkVWQpHFlB31b3awBlJ7e/RYHiWC
72h+DRFLjgJirA+YWgcUR+JHginvgfUZT6eK44t66uGUJjhMKqyjP/ouVvp7nP3VzWA4S7uE04Bq
mVgiMkdxzkanIjRAYu9Fvc1kJVKAPvlXaPf7RIfvzQoEsfNT0w/I2TA+XwIlxChJQAEA8STQL6wx
F4pb9neK9YCKlnRxGAtr7c6xU9Xg0r+8hLtqzIdHI11O3w1mPTHq1Mb8h6LowkyhireMyPnFYwcd
NxxxEVEzE7Pl+s1ODEUu2762zhi2ol99rxJ6IDDzuJ1GFwdmKFE9f4V7IfMT9k7VMginUDF1mZ+6
JJ6DyevPJVFRlU4SGpcRkHLdVkueYxsxIDz0dYyAK+1TxPmd9n8JEsyDR1Z0QWyL6rZ1+V+GpzGk
HgBMV99RfAz/J1Vf7Ymm6cOyKVhnUYfdj+9NUfHk70IKgJeUK9ScHDhlO0yF5Ks/K3V+L5gIwXQs
Ru7SKQfw9HY8HwKfxpygOP6QFj3KArUtgJyVDTkWMnTMsHCrV3l2pXV2I+Vkx5bKLguewJsGGk9l
hJWCRGTvorLBeXsMWiC+aqUT8IBpLfM2UkzAlni+1IRjIakuLzWoDT4LqcPaX5m5+ysoAAAiOlDd
cUiKY3PMMPVtcywceZg/8BVq5ERAz8KORC2m/OceIwG+iKTYS3IJBaebeHfchfppQaS6dWgT/RZz
Bkqj6vHwuSB14Lck/PKhqOpMBfqyCm1qlSU1ClvAsxJEOzRXF1PRb8DVBUwxVdZ6pl8jrPZjeI6+
LtsC/ZuGVSAtUs53jACqWnhbkKme1F2mOqTEOzlqL/Cstx6i9AftcUKg6tsT0jcdt9af+aLMLALn
N9PGwayqQisqFdM4Y1o6W4d8vhYt5jqJAwEM7mvVQzt1QFKwEluBv7/qN8syJTpcOGGqLDaFPelt
CRVcf6OPWREWAm3gYLIy6Clc3nsjr8gRTQFwgpvukCI+Jqbl2j4I2I/8my40Lz3MRigqGEKBvfsa
IDs9IjAZJkfLAC4tmiggqZSWFGIMjgjJHJ+T7fF1McItoaQj3vsv5Kc0U87WZp/fFAUI3xuuIv0S
tACrILuGIJy9JpjwfiXGpceeLQAtNI3j2PQdDUKx+uCD0VxeiZRDLn8ZPDPjJzo0zaW/LSyCo+Uj
/VdFIvIaaOyjfK1TXgYTOk5kYGM6g4oPNLTWkKHVEY1StP8CUchv/A0+NeTEGQXp1ULUFmCtTkYn
JXqqtNQGxpZ6+qnAsBVeyQarOaNZVxxs7Rg71nNJxJugsfYySbcWs2rvjrgnfgAM0fAxAFpggjkB
PGxiV1l0HXNukomHZxqPczhRy6OSNcocROQ/nZY8vgRfBnbGZQp9Ll9VOzJlbQohWx5scT2IWTrB
m86dLnJxdwWhXQ9VlCoXDNZHeFQGx3G5bkDAoVTeen2I7f2uDKFO5EZcwWKofRzoL2relxTo8xnN
yn6NX/FWKiT0HawskrevItS09VFOHwVYBmjQEK2TNbGB0+uoGMMIP3oDBm0/7KhXToZACbUlNpvL
dkpylFXJdbPx7w77Dl+a3AkXexim3C2ggzrPtazuYCNjOIeYfzvfzYUCBcrxhPAjpKkQENLq6VhR
OMAkxxlAd/4nR0yJaJcsFEAutOQMiA82RZ+PvsOqugQyzC3UAzRsAuXkQ5la9cXulbUWR2L2jL4C
akUU1iR+NMyRtD4sJX5dWjVlVTfXnYJn6++o1svzdC5x8/+dbf95NEH56v3Kf4hvCVQESr35SySb
KeO/gjA/zMTS6icrHBgSupD2KFxqKZvzbEgLqga3cVX+QMzWHLGXmxwfSN8EfDI/bjXraXv4t7KZ
WbD4WnxJEvN9juIQPaXv3Z2CSxd6c3MnMMOmdFemNzdEfKJjbLFBmAgDbn6UYytdmrGew23L6H27
QGT43nDC8vDJNtFlvdusHsSU3T3n5QrcbFiNli5Ws1tl442gEq7vO4EglC3xspTlmkcMvmRw5Gqa
NIFS5X3yAItuXiYzdeJRZcpwPad6iXe8gNRCw9sNlb70CKrYcYef+oa50dHnkvaah1i2RO/5CVwA
TpjlACvKkXACN66ulzrS3updeLz59OVybGVEzZnTn5LfV92sQSwv5jyrn8YkjmhHX5KzU/VDR5aR
HpXH9uiAywpm8RxWzJLW/R7k+sSgeepLtdd/O8POW7AwHk8COA49lnvCd9mpBrYaqFZPW4DOScZ+
MFsMuPpMeJaBScqbCDFUKISV8XcUU+EovfUQHMcc6Oh5qpvcxQ1tc7LnLnYyc9uE672n2/Fd+h2E
9Oj0xkJDPZKL3aRVMbBvUnTvsxEgWIdvnR9svGbpsVK5xVQcTTDfPpiRYHz9dsgPPQ9fW5wCP+Tu
gyYid6KMib1fsgJBa+OqmQNQR4+skmFUbk8Clvk8m5UBBCwbqwQs6DzS8zppXDR4ZMrosrWSmrs5
wozbubWfRJ/ljsNuQUtxUOhhz1qMIN817Ab1LPFmHJs5ASnjZjhBIcYMOxnens7PPa/KwmoF1qS9
e6e2trerfNWHLaI1P3dp28qvjgwJttewhmZxj1kV0/TdCYwSI9ihc3l6YPqRPLyRqGRvznbU4k4q
5vnHKwlRjTqlmq3pqDhwzkSL8nJZ+7PpKvFUTnpcS7wypt9+x5cHApUCNLo6rZ2WOF4bnxr4IJ/W
LlDGcsUqRMs2aLz8hWOB4CVcXM4/SIc94EuLV3Ymoi5bImArwfrAS6heNKyB23hQM1Zebr13u4zi
myDNFMn3vif1jnmwz4E/SAMZfkE/MXkJdg9wV+Gu24r///m569oryAmaDYdJUJPK+325cLHgAI+o
cQZeKRPH/e1+FSCZQmNsFOFBTNm1K3YMIdZ4mE5G4hZLQby4aUQSTOufmD4tT5vibHCa+UHLW7s9
PMi7I8uM4AHxzkQCtTa+fQRHRLvvAfCx0mmPgnIeNHwJu0BotfucIox+pULret5SWS3I0UN8un5S
TP93XXsmjQMC02YdeBXPk9nYkb8+TLKzjqihqTa2Wdt/PUOt8J/thyCYqJXa+LVyH9oXenCqc86e
RfZnyYw00SviEb/rbqTi2wkUD6wBBOUULaN8KwvDf2cndr286vQ6tZtgQamSUE7W89BcEkwGtce+
urW1q3BGt++5IsBrgmPeDhpQx4XQtavd+uTDJ3sUhp8DSzqA1qMY/C5YLO6HOUfUa339uOqMl472
WN5+JdKG8d0Usn1H68IqCZB3Xnzh9gCsNHUirhu/Amch3e79op0roZkB5vGL7/X0Xbv2ZZOZmuAN
LCyhO63WJAoFyca8FyBztOIWY215KhcQq5t9XRCvcN/EvJOOtHK0jIWNIo57J10XFDNdqDO88cpz
+FJMJJugUTX0VD859VXiEuN1OOacSlYMSSvpgO623PtqK2B6QDLQZNJuItnyrXGrZdVGKubL+8ix
+p4wXnmCVRR5vgqYzsoHJDbi8LtBd0FcQtrC7emEon2rcgMX15N8lIvwVcI2HEiXS67zI62Msnxi
qTd0Ibe0PxvF12Ea1Q4j8WHZBfgCKFHajDl8fBNrOQVFR+u0amD6dJwwgqk7CeDhFpD4V7ns3aAV
i1IM27yzqwOtXFQ5gGLLlWqed95fV0cgH324/r94Nai48hKT7KqtLynbBhe3uTF4LWL3K+xYm70J
bzZpxgW34AMQTMvCuJB+MvUf+p4zO3zAJWt3SFE8sFywK9ZBQ304FGJSYQlJCgPbDp5rcQ4XOOnH
KVywoKryQTUCBctW1JQMnhTLXY5g122tL1TvnhFZAro2diE00oDcWR5Mxl/5R/QtZRbUlKhVs4wp
b4IkYqSU+7RzJnw2T8CWavVETgZT3QmJEi8Z45UoCtS+PaZ/yfdBTpbrVM9MJtjO5Z1M/2pUWkLz
nRtT+6T3iHwV8l78c8Zt15/FJwT999XOyimuFSu4IXgf2p6yLK4C5kKp5VrTYsME9WRGWrmB8NKx
RdNOGiA1fXUXEwma/+Sz8sApG6w+xhIgYMM1JkXt+jRhSjZ/q11gpLtRexMjJklxjMNMesvkC0n4
RbK3uBtRUyCWHLgOlMiA+Ait7Rnk+NzLogLG9KEDiS2OtYq2RTDlFx1jNOWpDQ9cjDudeAC4XnQn
cIBZDteMDGD8vsv3eDGKoLSe3d8YP1QtU1tX6vj/+rf5BvGfBZHiwo9bc6dE0YCzlWE8kIzyCpAz
djssw8O+64aAuMyPBZacTT/tN4JFBWD0UpYSPpd4y0GzwLWaH+BfjnPJkG2RrOrFdPfS8HVbG7wf
E8Sj0hTv9TvUhbqew4rwGMkzV324z9ixT+5NGVEnAPgib4hrcC4a+DnH3B79bG6wo96B1DGrXgXn
aQU+9RMdH7OhOTsxY3R9HMxaISOAiYoYd1ORgU2fODgIABbVyGo3hIWaIraNHkcgF+n3I1lnFG41
tClfxYa8LJOB+2/Qp99bBrl1tiVzn418/AsPGVD8lLs3nIrT6SkBq888Td1zJWBu/9/mv+vOYm9H
ceynbZmOwdXoLL6mKqMKWqiEJwX6BwtXYSGCIVD/lFmLHybsBer2uhh77JHFTfMCKKAgzLaq/O5Q
RnNYlE4mOtNI7HWYauG/NkMK5W4xdpiS0H39qb/0Rh3Qfdl6esIrboN3vtCzNHotVOGtJOIp4bg0
W1W+0oY/XfmtyML1WcW6LIANwLjbhMMm1POKvUGXEkSpwmDNwO+PXt6ojRvsHQGjaQDNBFB+sWKD
Wu8Um8qdI1Ow2mFf75LZfxGJ+sA7OIJaD3cQLNJ26HkuooDIk/r4IiCt0ktN62C8Mr2GmuK9cWf2
I8EgptxM6VlN07AY2Yp/SY+YU20kKDgYNzMxz85JYCN1bYwV3IEVSM3rqAbG4rJUmmYo9WcGDAJ+
glXZAys9rVZmHtUI6lCIKAqaxFGJOKlqV+Q21I0N2G8yKAzsnD2wyj1OKJmCy8KLNz/zF15NNkwT
l0R13FzdkVVlMs+WO8ieNaOE7BlmRajyFk6QCUUSLuRlr8IsHSHTCHOYn6ytgfWLDurZWaWZ1pX4
Bmn2132D5xyaDojf1na6ncZi+XtHrfk6uqlRj0WNv6NTBQkYptN0Am7EWkL0JB88nSIEkCwc/GtS
ZU058y2HFoHvIcQAANBwI5aQz7tJV7kZqG/9bObKzD8elJyWXbakgDJcPkIutt3RTVFRlHLAlofe
akIP0P8S3cQndC6S65Jhb/3wXEivbJE0P3s3Nu4NsIv2gDP4CPf7279hT6eW0/Y74ffFplw9JHUV
9UMyqJK7z2n/UYNBgEeEPXwtF9sSr9a9DwPI8BcbyCe4/SzfJActdQ+FEB04mSiDhtH8Sy6eQS+N
2nn/n8kLPrYE5eff0gWwsoqYwSvYxAGAQTYxSKP9QqmkC0vdenU8+gYlDIc7P2NTd2g5VFcheVOz
SHQ/PPyEUNi5f/gggV/3oS9N/c3CKUJJ1jgiDP1ksi/ebLph8PQ+7zTVo25WVyJx6M0kYLyEFe1u
tJCnJSpGS0qjr0IW0UMnSwI6BmGCwAOP99qGj58dZPsezGUiPT31ohTaemvzF44ObMDiksIZN0Bm
o+/jW81VdoY+mb8FAhuHzz16X2TXPAd8DAhNXbrrKDJgaDoc4Q5Yy+kfptCjpPIwDwHr+ZtTqSyv
ATv3H4U8UaYxfF3Q/C50JQs4k0Ywx5QfueduIV/+gP+8Z4572vPvHqmH6ufGPcmKfzoeOTRlulDQ
NRTzCASEfGrW97FYHJDjFt2z4Czby2nnilKeai7GxfmCBRqgMafpJVQxZxDFG6i9eIt7RvPyR/fG
iFuc/4dzFBLLLyyCuZ4UVHtcPE41Aki0U3Pzss4orCqRIsIF1ItM9LbsMMv/334xoBvrFe20iUxs
nZeePGKgSyobKyZ3UDwvOPG3lufrzhs/GakqqHt+M9E8Vp0IanT5kde2WwBSgje/2vhJLGym14YL
Y9oxQkb7n1eDvEGDg5y6k7FVkqiiZ0j9lc3JukGWa8pk6bpet3X4UG7Wva5bh9CW5xKjH5uSSlba
oj95adsY9LcEHQXpG68OcWtR/cVT1TbzGfuRhuTO7STQ/fxYUOMzU6v9zm8V1tY08dFiqOeuPhxh
/VWjMZXwDcbogjyqbLQbxqpGLwyuSZoBVMUZ5B9Dps8YOFulDllI2+VdoP4XifAHe032SpkgLZWs
hmiGXoiFstL0pabO6g+4uNY98IqGz5Vi0QukC+XGXMyLpQqYEgMScuN0dYtYi78Fz6eHPOFi+I4D
ctihhEBS0tOQWpqnJ25Yzt5VsDI7y/6souMRmZvIEmuIF1ikOlafPWmzt7Uz48wbxLk3OKKU+UHt
dKxU43BGxVSahfBFe9wmzPTB0Q85psYM4X+8g2WJuY69NofbiJzyaTHAnwRLjYeeJIOCX8f0EkUh
Sh5zwGfywHx7rPDeg/VIxUvOmXN+A48wL1fQvdG0tHz0NkKwqqgTTjkUYxF4KQPc0Dk6D37ZwbBE
1wfMTt3F6sk1CduN3vTA62EPwi9asit6FBDZbhwhWOfWwQJu+cu8jj/W5fEIjl3WG699hNVYOx9P
qRweaR9a1PKbcsNN0gvRl4LQIm/X04zHPfFOD0E3nOYjvKLliR6XHASsdD9BNI38xulI5Fp6UPKM
v/ETsYuwNc3cgto8UQOQskHmgwayfVw/PTN7i7WSAaUtUpBf5JzYG4/i4OVS91DcIScoA7qsfVoX
oMy4559HP2uY/CB6PRtrffFu4kWzXaDuuwZjwHcg8F0rkfDt8thBCrztGDuJ2BbbfChnybItDNah
TSdMGEQrlYbVRq9puVKLeFQUa8pa7QpECdiBa5U1nlkHZvfEgrcP2BSmgsoFbbIOkUMXMFSutJDJ
scjwC4TdpP3MKHqR5BzP02DqvmRgOkWJJhtPWCNkO2iifvgi0k8p7vlRcgx0q5ZwRjXfIlFaWdDW
BiC6lIOldv/apthZCLU3vF2KPmQA2Ah3KrAMHFlcho+wcdoao605jBTzhnMUq65E3qyPkBX+VbM2
JEdqtRfThcuHsbWZhzBEAuFzvuvEMa60uq/tqGGyS6MO5N9/FI5UYTC1lkulE43YvqyqNGc4tf7L
GpCfsjMMVbwDW/LmXHxz7l28grp8JqH7qAAPFy75iTVFvesyxp1D3Kjm678gm4rU+KeloNUrbvEC
7ydPNqSRL88q2ZRuxP4LiQy9wFNC0CTrUfcK9rt207jlheNznb/xCf+CjuEadqRyOhqH7xNEK9dd
oAR5S27eosGsm/AvDjZEmRDHmCrDfvDr2hQ1boMfkdZ3UQ5kQXnxEvICUNOaw0zb0Y3viHDPlhQO
rCfCoytQWzwlrFQa5OH2W+yeVY+xQ1BZAFa58Dd1KpT2SlIYdIgclBl5QYxGQpxZ3NnIvv2IMoMn
bhx7omvJHWpKKHA7MlSUtBcWVX934SHEGoeXyiSH25baOcAj6tgTkk2978lz4G7eUaxVv9OtLBIO
tohYuQObh2gRcxbngxqCbn2fabctXupHIjveHgqcLdffnblpbcrA99IIgutYs7McjisbMXdHz7ro
PVIzHJG0wI2n2rqJ2PdQrb2cYgCD6FcrNWpfoarIzqi/4OIGuKfibZnpr36gGZmGqh5phjPYX52j
lxbeTLw3q7gun6CQiA0rxPjjAg6Z7Yz7JeQd0V3NqAeid8lB7FYccvTaS5sqgFEX8p8zaIGGW6Kg
SIk14TouMloSjixYqSBmcRGVQU/288ZZn9o4P1wO9ULdtGtEnEz5xX7l90aHxsNQ/6nAqim13qlP
FCS2GQ8SA4Zd+lo9fw8cxo7Glb336/GMmBJgY1sqiltEM/ZCZbJxZjkMhg5MTJ/Hz9IP0xh19dmw
lvsQdz4SdP78kZeN2VE7Te1kZXNMmfC+bMwg7/PoH69mWfFuEHlzg5grNIa6jQnR+KNUDwoEaUPM
2CasRWzvTrHQQ+96jAL02C1vFGAHImfTWGll2aBgk9chRUvaZokOkUPKTXYq1en3DCubIEOZ1eeY
wErHhDmPCLC5W+6b7rYSP+Lp1cU50FxZzQlP2VWJufQS9PUGCLNKMBUB/qJBDBSxRpLAsa1StVcA
fdtcyuLFzhyFzusgQ/BPf6gjbbfThAOqJv3j7dhJFc6EbxEaOyaFuBeQdU7ZY5SybYI6oN3fJE+M
4TACI89rnFuFBb1yUAJYxnetgu8NoEBzlN6UTKx9Z1ET/s2U22NhPlc453kW/0001xV5JVPNJ4hG
f0xXyAoVPreiQtarbbM0hyDEwVnmOy9spfY/MXjcw55s81xRMhwzaBl0u5FTA6Ah9YolQqs1YbGt
5Dt8rGTN7isdPiKJEgTwTiI0ud2lDC23txbzPiZX8GC9fZ1ohwQmPPIoJF6eXLnQ6InpS6m4XHA3
xdc3geSCUvwiNLXrdT7gFORfV2N16feybAWUWcxSdCbvgZT0h8DXqPYLLfVMaxfVO2JL1sQUtyVj
YKoVcie7eXzQcnKqEZo4UH1Np/FfmFhqkMCwMULuM3URjaZhblgQjPAhlPM0nwP8e8EqQSurVzPg
drqqg40GLFOd1JD9XBrOcyBWzuEBiKW1u9X7X/FfOqAsIXKBBq0fxhxzX7l0okJC0HaLtHZq7G7X
KCx9msvWPgYESihyPxiHiPqdR5kuDCkZyhcigxfN+mdLBM2Xd6Lweu9wLdvVmzLX0QAOsjCXC6oj
rv50QT2r8WDzGmcqR5uKS+hUJU3qkg4zS2jXX8V1wpcVwktj01nkTPrGNO7z806Dx+z6UyHKZ+lw
ZiIkqlC+SG870xSvB+ymMyBskbe6TR5w3eyWPXBBo0nMZxOxYWVP2u//y5JmUdLE+2D4fnZoL0q1
7iN0cuXILDznOe/qpfvXXL4TKCq4sURTWUr9qgJFeIVUnBNqIpZvXKHZkUCk7Xf/AuMnSZ/NPYVf
im6QB3mbTgz7rhwUML0dceaQcv5qg+ksKQsBm6g2nS6OSebZ1zUiPDkmebvYIknRELYKx/g+PLIQ
y0kcs8JVO7/Jm2MW3HdMglAUQJrBpN0asO0zdVWAydX3Gdu9rmtgwYCYj/Agq8w9+MhZeZkiOF5B
cY+6oZxg17dfZx61WRvJQHwspQgTUnDhhAfMLExQnFxh/BO+8Yg0HqAHG195CiGXyGT7QTQfgg/V
OU3c/Zoh44WB+/+msFbDU4A52CE+1fny0doZjp27SxVA9ZFv2ssglbgPD46GdPH4Z7n7cElEa3kA
akiwqGnrsVTYFdKH/70onlJhD8vzFEs4z3AQwksvjluqX+KyLKW88QXI94hXE0KL7/9NCVkb5pOr
3oobZWQNZCUYgjvbdF8x5Fj6hfBEZI7M0jSp9vjggqBlIQlDuCpTUCMixbF7EGEV42TUpnwOK9Bk
lU6GvY5FTTrPc5h1WAFN34RJRkaNSh4a8LP6Z4yp1qF8ks7NnDz+lVE6hNHYjpbRf+jGaYyuKAIg
yAhY29dxkhJNcVKcxug7B0JEwJ5B7RK3PEI2HIxBN5Vay4W52vvHV+AFMrRVRX1VmDflivpInPJ7
4P6u6yX2NKJhAKTsH99w7cDR/A22fnOp7fFsOd5dnwaHUarcvrbsyd57hDoc2kP9YGby4v3U3+Aa
yz9AMFIykx//ZFJRuyQGvXwU9oG5u9X9zm3592gFT09SYynxgwNJz/pVrpvzR4hfxcA1CitETkeN
LEn+eRFJK2h2LgZKY3xGLwhEtsQGreezh4cBEl7wadIBuiv01ZLf+Epk0snCSwCWjbXd7d9xJX1s
Q2WO4UbieMF7u4uKfNiOH4ol655+Xk0lt1u/I9ArkdC5ri0Qu8l1ingBGQc021U4F2Y2nRgBX8YS
o6P4SkIaVuz04hIlOT5ZvECuqTAjiHg5O4XEGjYt4jsGcHkHoa4Iij1aAhPEdurDlYwe8yLO08DM
kmsdcs7btZZVYz8XCKi3wsea1vtaETiEZer26uZjsVHasFO4enhB8cNR/f9ew7tePtetbVwYrUzP
hnO1VyOyXizLHhzzN+Pi+zludjg3kYn5NYeIWiC1C4h/agBFgUh8p8ZtdZ18O0e0WU1AvCco62im
hnptxkRYA3sVfllv/QxgAcF5MXllJ0UfvYbjOT/kECDsSR7Je6wfZvu/GCUNy+YpZJ/G5tCf8/u0
DgonlMtACr59rxXjBIN0pJ30dlE1bpo/pJr+2n4/uB/o9QDw8GoZ0eI8hzAq9Ws+WGD6J/fJcWLC
n8SUDlklYw==
`protect end_protected
