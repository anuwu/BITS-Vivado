`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HPMPLvpmoX7LOmPj78BMT9X1rCnPz6PdhVGZQ307N9haGfAdMGVirvGR3e0Glyn2ieoWqXA6qOQL
t0xn28+h0g==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nxv/BnutRgdmHnLyK7kvDGjm7WGfFKW2mxQ6xUKF14zS4ziz5pSV0ueW4VqAzUyEPsErIAEuyV6F
m5KCqRBB197Q2NbZa7O7tdAqboX6tPAJzbB6u4U/MmNS1AQcSgtfj5srMbdBzDa5pR4V3HrI0MRj
0xhV1BWf725FYPP4av0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F5KGJgEDQsX2btdjtRUlSmNtuyodIhGXEa3/AXv1Y7qgSO8gknBfiqj5HcIaVA9b4npQpDnNcmq+
1ONAqLeLhdOm9TES+GsTAkh/lClvl89bzfqgOV33iqwQHYIHwSsWMRXT9JSUx+YWu+g6xKpT1Ycn
8BCPsq4QUJIqL6W16fheEHB/lkMgnespIWEYJJG6R6zvv2zG8GiU6cG8zHrRjdvAj8kOkhmiMvSd
YjGXJSMfjw7ojCPSUF+nb6WWhUEmoMA/6lgSVaXRm00YHSZ09k7rKTJWSXFSpTmkL2WOsQhNS0ek
jdTK2KF5K6z2YOK4zkfHgZ+fB0KJyANaLLJH/Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lFuQXeJ0hi7qnIKAR+37XCSOwp8bGLukonngcICceOVpL87+rxvhP5TyNJ/zXpAWDF0BaRYlGr7d
isPiUStrvUthNyOqCr4vFZyhCdY8n+Mrv3OCvLoLQSarxVXbaKbXb0tPsXJCUdXTrCt9mr5x0Nda
6DAI8FBPlFMAiqnFXnYMwlUiSlkNWUpInuNw7+1eD8kUdckEUV1PDwZ0yjpFqMokMH9oJjN6z0Yy
65D8Tqo288ZMfZQuIimjski+X6EK157XbpyuoZIuYLJ7j6oaATdintgfZpgGzVvhCZtMbx6/SJtR
efW5vLBGiGs7rPBPE2T8fosHGOvmeC9QBSj8Ww==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q8VVvHzTNgU3tZr4+8ia7ylST+kbNPWskONHDOT1dTkB7cHZIAWyzXpQZPuEgk2wJq21PoqmVlG9
t08IYzkfC8vYQ2LRf2Co3SXc7p3gF2OFMC68J9Nf9D+/PXJCJy3QO4H8oO39l6bn8c56K2ARnK0R
mMIALbCWSBDGCWGQmXWZJ+xmDGs1KgTeiSW3bZRftWJ6K8l8BhMit8BLOY2Mi3jJ0WRhN8kKd6JT
D4NU1jTZT6jEtmI7Gnj/AXG6auTqDPHsVQzf+ZzBsLTfw83CFoO70xM997L5cZXlqz8fEDmxezkr
wWxPwJbJeVkRV3tUxlo2Bs2x1uVkXQeNVMI8jg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oUeTLA0HA2uKORUHo1HidNC3lw54gxwlLUkv28qRPv1pz7AEVUbIJ7wsyu2Scju+EkC2Ivi8HbBn
jxkeqRDTAwAbAqIKnY3AdyfojN9Hb8SMLcLnpWLLCpb6E0vwA09r7uqKRZ8wYAgT9CPFvzpQ3zKt
9DTLgQ3rZtFxx2nfCug=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fayrlym1l14Y48yZ195XboT9ZQmp/mAzUyHby3Y9qJTzDF+m6mRQ/ZbebObo8bu4VAm45JeETPx1
YI4UZNOK4IqKv0BZsAlzUfAYAmqmkmIJYbn2gWUCwXyKX5AoA4ONnlxEHxzZhqtsmEXvxwTEs25/
R7iLzeoMfmwwNHgPNQkteiR4zDlB76CYmgu6EOSUX5Nnitq1oh7qRuU8WqWN7lLfgIC6T7qNHwGD
RPze2yiP06fSG45jPrOn2fvBX9SRbUXjNtiFgmqim4anwJU46v7y3ubit/I6giZhz5PJMZfkDaFX
ag+uCMq4Q8ZEolqMBmjUjat86BdVd4Nmr0yUaA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kIpxh3qIIkWUg8aLJSPKvKhKTPFH7T8fisti5RtNaftS7xh3KDsGLYnF1lYhH2RVXgzbdaVqvtED
5QJazVo6wUFI91xgFeOR5jX+Ny5UBUX2MngsK+UZyZg5+EdtSiDtiJNtQqgjq1Rn+XQCGF3xP80n
7YvuVMbgRHCAfWrWw7ZJ7Y3raRzeIkx+koPFio7XnC+QdRJ0ItO1YtQgF4Sg1Ihr5TH8/RrNn903
kPa+anH9spo3SFCf2Ts11UXAGLdIBmOLMtEAKjjCUbtmjGSeSc0gn2q2I+xRTFcegLevlr/iuLTw
3lFndBAoW40xOiCDjWZ6Rz7J+jZhsRl3D0Bhwg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967968)
`protect data_block
veEEpIRLE4L2ZtflLmLyyYEUhPGOQikg+6z1Yz0UBd19Vc6FcDcPjC4ImNHzrHzTZwBAqfgKLP7m
ljrc2Tsg62nnj/jpbIQeFEqd/VjYTogkGyOlZhWjx7jKM0/1zQ1R1p8nY32qufTFQPqVnEsuJIkf
0Ogt0Bb/8RAyNHFNsnCBypaRB6tUSNBXXIm3F0XClKcTmDGKvS6HjG//j42QJuQ09PNJoJvU9SfY
JqxvM5aa+hbC5hZ8uMfAmRJbbV7qeHyFIDet7wSblJBuE192ZY7vBfYmIuzph3giLIwL3c8k+s8o
vyPzDmrcRp8HHeatCdSfHto227TPaHTW3W5UL6tsf9QbpRp+CCsvRu/EAj/W0sGgdOeV3Todm8I9
7DQJ4TmI6tyxVNjfcoLHLtr/L4AahUer1jAq4vdHev7M6sPSQR9B1MomX1LK9oV6PB2QMicweSZt
dPtLJAvDy211IFYd3nGRBS8cXkROV0uvT2oh2KQk54VDyBS03t0uwmzhmvTL51CEyQ/7tQJ4fXUu
KsTbUBx3Y+3x608PIeD2VDCTBmnCnaZlVYeOPwLVQn4m9aECWkgqtp5g62yH7xU4BkUJuKqRFVY9
bdIgiZApjKWO8jVxFmWWq3yVoni8+VXfWVAob4I687JxFJXRmYcqktl9TadsEyb3pzVNjvePcJuJ
/XFJA9SLyswW0LOq8bndd/RgDfEyN4lnN+IZpn/VLlELqMqOzBHBQhygqCyWNRnxZXvkFq0pL86a
FjNHE7kfxovE8a37sK22rpcqt0NFRzmsm6eYs1CXTFj9/hy7FqtRd0SzixqCoyFjkMrrwCKSzvOq
dYwZ9rG3vNKwRF5HIirmsejDAlBe3AdLn3MRXSCjWWFfgOZgHyNm4SPkFJfuhRDMrOKOsYUNpWzt
YMMvUYaC6ymQeyMcU9PCzxESzB6+BYdgpY0BpVNvhLj8R7kBjhVNt7sIuG2LjhQYkzTmF0Ucne71
Enzp+yzL95QvPVzA1mB3m3dy2XVBQJS+igHG7GPfbd3gX27PzMuwKVtVlAKV28XTCET5T/IC6Fgk
qhG4Sfp7v3uvZAWqrYj1M3kI5wZu5IrMa/z0Y7Bppf86sG5H4G3ruHyikM017VXIGXgb7SJF825i
3yVh/SOcXm3YbvfIIxy/gNPBsvVFqN3LuGS0vFjIHjUvCPArr2vp19i7YFaAdLB4jnOdO3chgHin
5mlLHGL4CAih6iOXScdNABBKOJOnnx46ajLK24915F/TYzNVKEAKfCnvIR4or2q8bOdnFwYiRfVP
jfiWw0X561vcmmyuolFvTWzrBIVGaCNBNbNcRIJp7UCwm4stkggC4Rk9DX5vkmSGuzGKVKuEwPJV
s71F2JhMuetOXa40UICB6Kgu9Tmk0tu0rPF7BJNu7qz8gcDsjHyCzRqVkO0PZBDs0TehpK/cCTxR
jVjbwkRJTOYznkB1rFaFfLjS89nptaM1sx+JJVHtvzdZq7NODa8NIWDQp5Z6LZad6uTwZ432K9p4
miSq1dzTWn/TZQFJDUFAsU5RzVA3G5hI/aUefa0cMNQrVGIUl5rUoIjWw+RUqW/tYrIL4PjL/D0H
OtrkTUzDQNMpH74EcfImq93KMCz4yS9HeH93B3K3o1yZSiiKAklKG4yShuFYmP7Oy0Bv7s2+CzG2
KZxDjUz/UZ4MOZAUOE9v89lfhDaW/QZdQcwYdBaW3SAaZRjBcOo2h7zc8oGRvBca70OlajmUnXz4
VRMhxIfIfzteZj9dQX9VjPOvymAuF44MyZPUmV71DAHhZUnC6GGSafMMEwp1uYZGBwnbgJzV2Gua
nf7yhLLQHG76HqGFH0niygx9LKhNSRMtyq0FeuOVsl8agt7XSxglVyCkQL7XTKTC+rgb+XFMNj/i
uP5pG4EZ7zDGKXxcCldWmTwE9PLXGb4d2FbP0HzytZM9HsXI/z4dKU3i/VrB8LM25Mm+HNuk6vMn
NCRmT0CPQjbHL8qsZfSihssRbdGET46YvWd+EP8VOqJiTWHh1JPFlQmFwzfr1FmMSV48MvYdCST6
RqGiU+FjZvb7rVquPL6Z8MGJJ/i8fOHTW2k5e548HgFmFpdeNqDv2K/N+iIdFDXjLUecNa9VIXeV
zfSOZJBJqy4StN6JD6Ll+K6OBc8dS37odlmwaVE5eIea546KMtRNTGZMSDh72bbHdX91HGM/Iux/
j1nVtl+YHCigVoz/qBonE1UwtIokQtY22mfAl+uCOzd8a+aE+sMA5+xZkZx1/tl6wc9d2AKKprjL
3nPlFXdtzfPiWGB54F4jDiYcsA2001OXTlAbgrVdLm3Zt8vrw3hYmtLl+l6NomOsFkX5+vqINxrC
f99kSl5qccvJveQ8PM+mGYhnSHiSH2/dzbmth/h/Ktug3+L3ok7bxFGS3isJCz6aW29AWL0WePSP
+u2F/DSQ3Itk+bpWzUc2wBDGS4Stv4OQ8u0VzIA+herUcpEw+FVrDbIBEBRcasqlzoVyqkCpMkOM
3MzFcPqEzDsx29q0Gh9CjZz0mYPx2f0lJyzGt7cjUIQFISiocIX1YkmvZmPc88Q3ZfWTnd6lXdyw
4IX+QtKzKT5/QWeFDDWtCU1iYl5ffvNs5pkhX37sC3YX6thaIvvhYYo8RToozGHDRXA7HbI+ayW2
M1LcToX1rAoZ0O+qInhsGGWdptz5fWseDVbpm+IrOpCLXUroadDlamMdqJpJfDlDG1JlUD12ZZI4
7SE1IDC4Vs6Te0RH0ZRj10rj50ICFOHvi6eDdX9YmMymIPITrHtAbtqtoNAKcK/uyEMvwxqy3R/I
VmF4YnRvEM/oc7U3xXxL3vyjHDtjVjl9CR/kXa1HH8vNVs6WL+0qRINOVrmLtiX2r7PPRVTHMjL/
0mlM/pDf9vTFQglQ5/8Pv/ULF6M148QCjTShlAxCS5LM31yaRt3bxsjmMDAWI3vVnyeqsKnL/XPC
bIcFuYV+PkwYYWtYkL4fyM58A6Sg0/7IJrv6Oq7q+xZCHeqor688CPMvsvJUIZmX+yUMGa+dVWhQ
LeCt1Lbj/EXJ4gI1XCDmUWsBmo7ls1uW7g6r+jMPYASVNDKszFH6xwxuDg+8WXbQmtgwc5NZ9jIp
N6lagfRo6yzKkYMHRr43aAKxGQ2oCwv20P3ppwKSyJ8Po3+BcoAfc1aB7YbAANfzM4iG+6q4rTCG
unil1sRkQfHrUlsuwFlVWGPJax5I9LfJzxNe9gGxgEfrP8m2bndSbzdEexvs5a0uHVNLDCEUJ51f
ELVULf7oxTz9QhEK8cJCtlrGgelu7u67EGjpGrIvqkMxL8aH5l9tnheUpgSadtrMZyk2pS2NPwMU
mD615oUOaXlsNAcGzV0tnQ59WuLsUW2oe1/4CTWp++40NLx79hC+bl9IRjkMzIv2l++aNO9lRyF6
aLnDu3ugvuYSiimmYkIyxZDxqZuyfhfjX9eydUj5iDufQzzoCFyvmOfTDICqTDObhq1SY7sGZWi2
vApzsn+rtmmoqj7mBN1yuZJNjiqUwmAWyxrLw4xhHWaRkxv5ggD7jn+cdDicjHQ1YKY8laxkpk7S
V+AvfFnCXpyge2F8AHchKeRRxGc6EfDW+pR8NeUGGzfD9zR7REQ7aR9SF2UHA7yEOliLKSRjPf9t
hCP0hShaYUt81bSG1eDtBJhnSpuVpME31krKpk1IvwUrO7vyN1eDal1o/M6b2s6c8Yaikgx3wwzZ
6eRJvKQ+Dwi9EQSLWkLqZUXYgqNypyMpUITWGdN/BQyz3YWTz5aShmXAV6AvrxuQlAhFH6BBcuSl
OuJEh65Oo0G+n8bOtbyhMLooDyfwec7swckTplYBoEL7GjXVfLxe8fCiB9gR/XyGYL22kL3Z0Gnp
CVUSftHA4wFez/4pMsekRSFUaOyjxwN/eOlBLlUpjnsO93NZXnfBG5lG0rE62ELGY4/4kvHLiIPA
UR7fQV5hXfMhk3bxLZo8E17RKsbTB5oRfYUZI1P5/OgGlCYJchBnc1uZ2mQDZfRdnt165Lvztl10
PQ4SpcThFDNOLAGczF5Ry0oYsdbFolMeb1Xy+2zYE/u3PiNxDZlCn80EzFwADVqsX5FENDEz9o2m
vLDRihi5ZyzIU1wu9Q3cCoUMtmKuzvMlu7iHBauzsR0oga1v7GX4u6wrWL9pcMhyE3sjLgfPgaQC
iEpH6WxdJ59HpD7ddAXXJG07pDze+cbpIBmgr75r1FsU2zbjXuYhnxPDYMRKGsTbJfpssijX5zwx
ToByB/w9PzGETubgh8qmE6l21ECYVIQk1vwApYu9hbSiGslIx96Y92KYinu0/P/r3l3cXnlrwISQ
s/BQr851VAf35c1nr7H6jIk2EfCLYnWRmMC7D9PEqTNfICZqBSotzp/ykEdYythRP9LuWMDfZuz+
93coCQH9nZ+ud7dS/lVO2TJp0TjTWBFmJTojvvAFJ6TJsGTDqNG4NYb1OLU2qhXEpRgvQegB+cZs
4Ae0GqBrKx4Bot146erW1lZK1ew2uNltLfK8sX8JCLfMJ0ViDWB7C3eq6UJjJjTK/eldZh4lfCK9
r70/A6jykKIDhfuecR2RFBspG0dP7RrAekP8pmUEYZPSfLnvtmFfgnNtvDgIVLKNS7KmSf+qq9cW
WA7vRSGWBq7GoSFqO07VwzQDx8QN+7IR/qoRmzPT6I2Ws97ihA5MqDtTndCFmSGA+ErOA0orJGhB
4RibNtgjq8ZDla1+v/TRjvO1drXUQFuk1Uqv6YaJSgYOFQUjq/cND8NtOyJkE0ZqzO01b5Uqvx3G
5GqyOi7a2rVVXZp88DxwRFOxXmkslSuMxrEqiNnrw04t/9B+rF2TGtFqdqs4+jYVBIjun1KJVHKP
vrCgo9L8TE4WaL/CXeW412+dMIhG8dUxY8BlOMmXNqdaqLwvO7Kfzn/vu/ch2dakrKYqETMoXuW9
x63tqjaz9cUrsZaEoEkbxnvMXLNE8PRd4oHKItstpjyqxdDxGdwwzcen/OPad+txYz4xxSRfWkPW
N8ISsMcavevgmLqT796naaj+bZRNTkTUlJ2KUdnmpp+oBfsalMQ6ec770WB/UlZR7Im821tsEyRt
nzfVBEW/BnsJxrVu+cppy+JIubp5iGixJuTRJTwnnNbYiv8Jpy9p4XuVJPYfLnJYn6wNNhoHLgm1
yWtgzeouZGASNXOxIzcJApHeSpZoruf/yAwLsK4Wi+1km8VhFQzhHBEcE0QCvUMjlE8gYG7DXp4c
BrlcOSsGIhEBJs8WyDCE5dFWBQK9i2l77iEDjCR3bbu8G7pE6GxTIefB1fTuvfa0oQ6SZTWmEgN1
632RxQrJm8hq8ACsfpFG+sXIMLr7kkmN79X43i5E33WHbHxSueclUXso1GhK924VtFaJDqOd9ALM
laIoHv5ZREmoEEG9b7kkFaYWaH4Rhts+kkcAXvwkSR8qb2ylt62TJfZsEZukNwNE3P5f1WUB7qx5
tzvW3/MzrBV3g2YZNyOgbA3R8cmYWJNL+pCKCnZ2WONO/MQFCdA/M64d75FiCNcCdt8tpOuSHpzd
vokMWKrNmAB1zcNCnkaFwCFo7/Sh7qQEvLyN6TxiJGi5ge+jCwVRVKPM5MlBORh99LNJS+3FLnWv
NFJ1sQ9nq2ddGQbpGn9D89tyNUgkDbNzZc+O0GVt44QoafFIeoHuJF4XgIQQ2i6/ig+i+xC2frAn
AXe8cGVlsxiBjICUePGWghKKAiHCBVRbMGS+zEfEhe5U10y2Jg68ahAHjUB71aFvWna9YO+MPkWY
bQdksJTAmuhvBkahOC1YV0UPPkgxmiTo/kXQ0sZ0T+pyfrMkf+8wQlr20o1dhVdeSz92Jci/Lj+U
CTTG5hnciu8W9BN5/hB+4/yXCSy8ugXCJw1+tLROAnVpXbvnmqh7EkdrHqf9WuNbjWKcuaclwFAS
XQDEG1BS5DSooboxTQJTvysFB2vt73HmTbq6df16t30qIKWr73WT3JZNp77H6aGk4sGLQTZRaHJv
bu4roRzucM8g3qCwGhYJQt5rKTp4KginkUGsOauIcczad8DlCu7zVg59tRDl8KioGs3pSOz2Y5XN
CSCx9CynGCb2/WZ0PSDc2CtvlO6W2OOKMhzBG0s6F4CSKyC72bfZI1tEHZcChetJojkaptS0TnNY
IuRbwyNLiggGtmOrhdGuljm34Kxgw0QeL5ivR+uzxU3n3HD2RlbR5w1Mr+OsvnQ8CDIEmoXiu0Zm
k7FWH6gHjVZI21iO1kLGWvoM7p51rVQnphE9HaOWbwziO0ropS0JT0U51HNQIrEY46EbYUhiX1qX
+jxepr6/gir2sMmo1dMICMBxtbZzT0b37/2oRhZ2whoZXknLTJkVoA6/8F7gEu/MShYS8sIq33xF
B+v/bcKurRg4pSBacWd4ORWQPGbu4/irsYzrmHcu3nxKKGUTnTsl6SyKiPardx91T+4c+HZPpuYG
5gNokNueAnDv7H5BZBbDyZizsms0xZr80xV3qLwhZbunJbUb0D5bLKiw5xp8QlEGnhyBDqEELXzN
uSnjZcaA9MzxhhnxwGxY3EipvNyTKpODzuHam4ZhEsryJWoMyyCfjpkxAD8paP0ok16IJ+nkumy4
iwxvLB3gdfMznZrzF9O5uagM1MSe/0ghWB2qj6WoHNaj2SFGEaJcusBKrwfb1FtH11wqB51WDW+E
prQoSCiPvMtlkzSDV/ksUgYVfQ/G8M3WCdgQICaOd3AtD74KvpHnfJIhB/boWuZF6yMceXyLGvWR
eCC2jmMCbS6StJW7jFs13CleZLyq7p24FcCgY0h1P84f1pr4CfVH7PK+Rl0MCoS3Epgt2+ugRHDg
Eyd/A+pLpA0u2Yh/PL0Q7xMsRES+ONAnXyTBkn4mZD6esWzQizdz8mOwpFjdVuMkS/0JW9xBYQDh
Bas0gzOOA78NPS0qeUXZIBUoebnt93LFQqBB+SifKKUbbwSBYmL0pAGzc8f2h5+NCQdK8JNf7BGG
RHeHuaFNoJKStCu087kLHaYWK1GTaNSlCZ+0YOvkwaW3iPAv+op4DtmJ6wh7jlSwFy5vZ6Gy9eqa
ar7x2FhHMGMOPeMv2KlU8LPl7NWHrxIxhPHYhYP+cpTnMdWDXCbM3fopRWvixkMMImxoWqszyLtn
3muWbxP3hUKCF/q5D70ZgynSUvnvB1/5xccQH5GKVdYmVZ+YLHDrNNQLFWTWOkYx1peVkgRFaKMa
PqXBxRATvQ7X01asxKttrzEUXILpK0w3vInEl+202hFYPVSgtHzuW7nj2VZvykKOpp1UAT0v1cOt
0O+IuFLhiTo93PUtt8VCobFBhFa8w14xGObt8kuwjDWdSfstYErI/Z7Fch6aupU6z/sbU8X9n+x2
3K03HFv9DydWfVXObUu4AB+/IlbVJpYjsqipC2tWJKpTV726NP7dwEIVKhkec4RlA4UpWfgd7ZRP
LjDjMzBB6BRn9Zfihjc6PtV+65WcqoqLmw5QeX42HyppPhaf51qX3jXPeG0Cq8E0a5A/dB6RMdcV
47Ewuq/p5ANokXRVQMF1Rw/+vlK243d5g9vUwub4/Wv03pOG1u031+Rw5UlKad7fa5RmKRtV6arY
7PeXpeCUgmC34DTVuvf25+eNJXsuEedlKwOzw6Dzndpxt5aqEFOq6M7GsbdSMVs7pE2JXiB+JCZT
sG7SjLM1H31HSvxuzPN7CJvh59MOT77Q2wXGYXXNJc7/IAN3zY94WabvD2eFgGSuyIsRXz9Nbr8K
TGZKNv7+LctFWCPPFLRqDVr8x3iD3dAddUadEkTDisN3qMA1L1AY4Saxb5s8qStrQA12HJqgGEqS
GjZb8izXDq2uviCtAKq3bSuqp19hIWu6SDov0DV0eBm75dOuYGK1tSBDOHafYfGMdixyWV3WUM25
RCgruHOA3i01Qvp3C5VdXN61QFztF+g7x1NcmFtz0g/sQwk5hg2ThTMPPV0Pm66p6M5oQvizeXIQ
Pk9ra7J+wNrTue7QmAqKgmejazr2Bh2aGeTK+L4nOATzn/l16J5cf0xxLUcB3765ut49ms8v3GSv
bD3/MPBBOaMGQzWVQMGOgFcF64OaS/zSNXcs5w2cz9jWzxLYHCo1teQ6xsEJxdaL+EtIkmzEetps
tsbtkYsSpB46FTt+C5Kd1mb+bzaIX2C5bLavOEB9x9lgACEl1heZJfK5qZFcOFNwNgbRZtmRPoRq
k8NBqj5xQ3hUMJ8GygW41r01pa0zeCRDfXFrr1Tq5K20H7GZvc2J9Mda9X4IJroGDZ4QCska3pBD
xyuDS2LHKtPaAZlSNJAAPVCIMnU1SRalOgnQX202n0F2oBSXDnAWu47WmL6Gv8KrxfJHM14cQ8kx
6xwIiLI141+McDv4n/usBFTThw+/9sxvWUaOXqhTnrW7BxeR/zVdibtXWrWzkDVHdSsOxFuJrjyo
jTXYXAhSmkbarjF9iLXu8smACeLwj7XvtTyg+HfFye8UpcIGsJqrQ3iKwVqi46JkAHLMgFCBwvFk
bUZSM4L6EHQGSHL9WnSNpwKPXB19nGvjAIjDjLlHNn1A3tdJkgV2Dv8LjVcECcGgpbJAWG+UEx2e
pneRHLcycXlT5MN9fXFIxDjkxzhDdcWZgRvFIz43hre/YXWusKK7lcXyDw4tnHB/noupYw1+UvoF
/HubhjmW39z1txvwvgEZijwDw16fX6F7bC61dkE0dl6cE0mYuCQ1PpOp66L+yS+YJzdJytXKM2M5
Ns4maDpPV6z8MZKTyXifPgfc8k4IUSCjo/75556L4cpXHxADh5rHD82NqRNZ582Q4dgwPgdTvWYB
TmUbjX7t5oZX8MG2xe0NVo0LbQ4L5wvDVV4BUIX9HQCY01vM1KD1zMmRk98FxDOKSvBS6hRZkUNk
8W9sxL5j8b0zjG7omehVAnI0+OC5z528cwUWqBV+kYJbssLpaMOwFKYEvi5xi7JOqtRvtfiUe2PQ
ZCxhXwVZaGl27nMx5GoESju/TfH4IPQEBVIIwNtZCI94a14Jt73rbQ7i/aczGeVdT3M6R2/oWq8g
lEXoK8Y9I2f8gWVnZD4MZbaI1KSiy9vWoX5myFss+OJKKTdijzuo+eUapC0YhpO9ChGpII39oTJU
1t67o6DnpoUoNNyLdBI09XNj3gcMgttJZWT6aaTsGP28pEdCW+BkzW4X7JKjW+eUKO2k56oNOn1g
T4jQruX7ZBuSff1wJeZBfIpvF2U0Aa/u12fGWCuxgwxeSyuNDsRtwjtgejwoQ1b+nR6xkVWdnFkc
mYhxVdEldxPAgQM97YxW1eIi/ZI+iai3GO+kwe0SGGsqBHxUgDlzQ3fJLhwit+nui8aHzqlDF9Bi
7EPXUETHtAb5zYK8H87Q7VD2UapmXL8s4v06x78WEx3Zuf9VFCHviV0MeHT5HZ2y86/zFRN6mZo+
igv5JRvVmRAjhpNlIa358t0U+D1nbRZi2AkILBovFkNeBq1xOSE0MU+4DhlX7y8B0cC8I+0ZweRh
8SVva2GTo6sozK/agVznGaaR925pU4mH/gNq+6yOge1PXVQQ6+8eKSKgF4yEv7j4x04ryYIkD4Z1
4cDOcy4qQYPcAqNUZZtwn03IFRdaxCvg91iWehD7UX+kDHLmxqvuvx1fWIBh+44XKvTzecS7dgyU
ZPCFmv8qT9TUJQ06Ag42GEubFQq3R4Hz+q3CZTkhuibZbLzTmSqs73WDKncTwIhLoUzxGZzN8Ii7
VIE627H8y7pkEaHh3QgzEcExZzxljLYkWLwonM4nvmh3UAdXDXSORpvA7wJ6vYn3SQsa6cORgNAL
quy+d0rzKDvnatxx+pwF68u5ThUHGpy3hb9wG5eWqjogTYvngi6HsIqUuGE5tXB0oDhNTxawVrYx
v91eWTgSykYbVS1RIQ8wvH+HT1KFz5ZUwep3avtXZb7ajFh7hKj5k/oU8DsIFyqEoW9WhBqVRLfg
mJUe3YKA6geR2bWegJMkwGiDeFcvIl0VAzvt/xxbpIw5/6CyXw6xESR9vH103NCuzCJ3AOyIEQjQ
cspA8z03Knyls1m/f+EG+gHGzMrOwzLq4IEt4hrtca7di3hc8+nJkt1AT2WPSBdWsc2cW/kckdpD
aTfH5SCUfwppEZjYpFN6sZ2JvV4W0YZy7U1Yd2myD+gpVcMYr1Z40z8s3+vAaWGPV+2/i9w24X37
6HDjy1ECapsyaItP8imagG23A1AJ1FDM1b95qMSKAXTMeQ7xLYKFM7Tfgt2+6fflWK3a5IPISWlB
kCQLWrUKGjRyetbkYIwxXrrxz9EF55geg6tvB+t645xjlvV272sH/A4Np4qJ4UpiruSBw5xGnAJC
AzKysCTJOXC3P4vblbmVwr6ZWmqY5KRfyzKPUOlDq8wrgUIbLAEc/UWgL8zccXosn9AttElPONo8
swXvvj5SarCzT3NTT/YWWEuklp3QExIpCRuW/r9omVtdiCazCraaFg61wupRmP+5P6TdKq271SAl
+icjLlC6jFet/wqkx6kAaoBqjSV2JcZRLGX33ssbWayxRQ1Hz9M9s6AErQcCUW6JZQkNLTVPO8p7
FMEMzTP7D/Bne7rNM5OyGDlPMO17N7ZlazQnOIon5dyB/AduNmnYrce9V8Cn5VZhd4ZmBUwdtDAa
fQj8iBoNRR9Vtp7YSNB7Gy64MzP/R+zvSiJitg1/Opj/Xx2C1oAKfMMuxtneZogxjZm0geItujjX
z1rBqotR0dU/I4fu/EO7uW6ih2g9OC1pspeNCZZBMYeQG8fkn4uQ8C3xLrcpEIghS6PD0NJWz9m0
AJxNF/Ci51Y60HPGo3EDrZJiCQ7KPgm4UrnlSs5vtggTrnppI8IpRv3xGq6HBmDwAe9Ec7jt9lTh
OpIKgDcmfMO5PExs2dB2Mr9LadxUeTI6cuX0dXDxILbTXrTxoHAG45B2l852GmZ3PmPuGEooZeBO
zo+t03QBOQqzZv2vf/ic28LCll+nnyko3IK6Szts6TVwu69MSaEE2pJiotsXkskwWNsovO68SjmS
NAHJpDMyYCXtYTzsRx4kUwT7mx8tTp7PYgQ7KYcmvqo2eo/zV2awAfumjrHBHRkWVXYaHes/c/26
ZiVYC+NBJlMUJdaZP4vD5b69XpNwVUsRpfoeUB840hwwabRd8dJg4GH4cSXM4pLVF4pfjCYOAdeP
HD8a89wl5z1dwHF1cxA8IqS8aX0HE5G1QMdePBTzAFl1zl7iW6rud417XWQKq/Djf4fGxx+/SZ57
B5WEhT3HiiTWbF98n2EeOJHGHEbLbSUkukxDOOHC+OmkoVo2VtYBAsi/lLhXURZ8ckhzKobP0Fwy
kt36iRIx5MNA5smSUgnXI0bVkoKBGru6ySRQorLxPszH7u6xqnQ9E267TZVIi99kh9QpvY8P0vKF
6j3AKWUwLhSXdvJvEPdj7VvXjXEupjE1NSVeCByamL9G+MAzu/8WA/yyL19YcQEPCt98NngnM23+
rXB2QerB3H1in1hJZl/+yRHQjZ8X/oMuQIA/++HJCc9vIfGJ4+tk7J9f2aw0xZsw4Q6IMyO5CYAZ
YCIhnVsHXizYtK+bnUBZbHDateyl/nCeT3Bcx2qmarO0tUVXQrJH25Hcr/Sya20C62qsCeRAsFG/
JfFTTbnUBId2hG8GPM/kThQpNw6sIIjZqOb1itxfH8qSDLMQEV89Y/Xq6pzHFzDHj1g0zc0nNjeX
d72pTX9n1indJOklopEKrQnGwL5TPrcZyK/Df4zLebOrTsqJPJxSkJreeXWrdJPrUy5NXUGu+0bS
1ee6I3B/P52LCl4PMfy+/GqSHqhd0uwozX5C7B1QVLCaZRG5CknJo0+ngjGTPmrHDsMMKPjJigRI
dEpLQNsHFFoyBIBoh3id3vOeWAgYtao6IjpJMYQqoMNEowzWxzvYHCz1ssKYgkTRSVOxn2huMY5W
fKK+uNCm1qo7Po8xQf+ksG1+PgoidyKY5vsu/MS7AdhguSopYjVUfve2y2EgfOwKJ/lI2/D+6uUY
qD57UogJEp92BS7qMyJhb9uXDOrIauxWEhYuMnRc9S6n4IPnGWPEYZ6aWKzy/8tQkWmd/BTcpRLq
I8THYUzXlsJkbcJoyloWX4YdJAXPdc8499GJtLt8KnPJ8vN7VK2OTgY8zXxMBldYEF8M/A5GtHWY
rNUTq4Y42zWejIAz8J95THkM7rPEvhZ10PguPP0cL8siBfjbuS7dV8bdt9y1H6xNbjZrj9Tzmdd7
9WTF7OtRbTH8/AWJ2aK0Ss1f9025hTjWPfKFPxrlCM0gBjzqmfdb0JY75jkbYWEnMSqtPv1O6PuM
rJzQFyblvfSOxLJ3ptmuq8g+FGF9YvXWuMiCnltBhTYq+yNt0jLovn3CA/g8TszTmWa7tZeVAhZr
JnqXQysbAbrrAvl8cpmkXlD3xDOSojkybLmkxckbJHCj1YSE6Tl1BJW9WWiD3XxOO5vGhmKYmHF3
6ez/qjSqxVxCoXxa43W6a1YUP262jmigKg0gBtM14Tv1xO4K2Pisoso3MtyPIty/BpkyaIvyqWP8
YUZU5Dgc3KLTn55sUxMLeBBiBg8GtMao7T4WorztiO/GVJ7HwR2hcBU8Cz33q7SoxN/YZvhjGA1w
Qj5p6vU+gLBVWb5QLRm5wsZLhy+yESylEUuq4904EWioT/zQvDSvvaroKj7muE6K0BM0usNwVmWl
31/ZlicX28Q5yABCOrnCgJHJH5OJHM04g2LIkJhPm03x5KrKUq2NSxgd0s0/G1LWiNOuO7NXorTH
EOReQz7PyGBLTJoE3JnMBio0tPQRU7Gf6+1/ZFGDaiw6gMQdJMhvi5fFkWKEXeM+mG7NybriP+1k
NeQjtwEVRR3JRz+0zwqI3sQizM5CnS8DvtOg1qvLELg1cnPikb6DuCa+RsoHqRYdPWQn+2QMoooz
4L4mlg1jo+CwJT5f8F27UHlHfWjro0SIqEC6++f0HoYZkqf2r5h7jwBISnuLoFpDUY3nJy5wU7Aj
eAyuStQ8YOU/yb5oD507kU+QeND/ey0kNb7RY86Rlgl1++DIZAbZTxM1L6TILm7yUlzZ2u29bomU
+Qqlr1z3zo8oh6uJCKVgEhX//gFHOQFtBW1yjG9rxs7sBBtqEaZVK1kBRTZPY6lurfURKpSbTICd
QPDnBvg1Z99lRODmRbmPryap3LFjyfYq3goQav0TT2bqp/tSjQsBWxAUF1g3RGMCY1J9QsFiuj/x
8YX8RpHxEXypb6ewJMIEsyGIFYeznO1ZDyU9c/asqtHpV6E3BePE70uq76jYzcOAzk1wltwXiLm6
z4aNvY+STluRRGuOFXZY8CllfypRZlNLezHiwTUfWSoc1TiwjxBUcBMmAyVjvRKkFAB9nXYnXMcj
Oj0mF5RB8C9y97iBGCPw6j+Xruq541fp3oj04zdnISm+fsnQ4mDFk6R3mguRI6oekmvk1w8SyLpI
bG1hsluOj+0H/45PeQ6toyFw8KDZlM6QhWLhEeZMBS9hx9UYJCfqKeG5BXY1OjiKnf+/X/dFwuHe
3o6Q99DK9/wI9sjBsXgWDV5/Qa0OesDFPShmAadWv325oRh6iu1uvRozJAKA5ws/26b04OY2zGvX
yh+g06YguLRkqZtPcRc48aba5OZVcQ4mmKBNw5QEHKcO8zN500LkSgGWD6+eBK56esli6KV+KnLV
OTyhq9h/8Qlo7oMGN1ayXvd30uU1K/drlMpKvBngv26yGyJAvEgP4YG9TOuR6q1iDVW8fv3D/dPl
8yca3kdB1RnYsvPRHIL8MQahcW7M1/j9lthA9way2+DhwAXMllwKMmiA97aMg33qDIqlhQvAgL4m
S1TPmLsWqy8XojwZl9ORrhbUrfY3VUwjtr+dGaJDMR73o0QvWBigauK8CcKkaU9uLCTpbuUEYU9d
LxiLge8UQ5lWC27lsUCtepcjnkv51ZFejGvcaYRZegNo9uzwLH0TRh548bmXwYhJU5/UDtVIuwtT
jT+mJ4emiBtQoMG9LpCa9O334M6Sy9C2j/9z5X4nua8XuvVFmB00qGPebvPV0+Ql6DMy4WktZI0F
DghKwgHDhUYGbhWqM7TIgXdbMeJXPRswu2zIgNyxKcN+UB6yEhaKX23iCtwNWY1pLFuY+n+c8OVq
4Dl4/qWfYJuxxDmqCPwnAJYaQ/VBhX3puxQQfTk8INaehDmmP/ZJA+pvPwm6S5TdCz/2Y4Y0zGml
/Xg9C3H29SNZyV4R1xeUIFurTxN+ajpDA8u8F4YtfkXYtvD5xXDVje5ZI29UmPJWeqQWpdNQ8r/P
8C/mhBcWEL1wlqcU16xH+RlSaKjGnVb5K6H80XlVlNZpCEN/vv7jCzroug4Z3tWmtmDdcx3xGcaN
gYXBEYx2k2jBROQEqzkfGXgozrxtdWNAqeXMZapNUqHrDqFYMskE91FuzBeEVvT3YRows6boT1g1
5R8ol5t6JH5fUhYgKqsDVzzJiG4aIlpudEeMvRpOvnqXcMq441xU0LUuXalWmwgIDvdchey1LHyD
r6RSchdkDkmTPmA/BrB3mrGhZb1IXOaWcaRyeHoZp9ieTLbm0pTiSr28hP6zQhjLqA+3h9HLn8HC
UsNgjZQamZWR+qB1gGipV65NGY7DQRWIX8WxXKuF26jFBjaSbTeAInIsIhx9z4qqNzmhVy1FPIjA
eI1eJB81yfqfLaj+OswGQEbqM84uWXJn2HOJIgdXawxpODiEazuYRYQKmwECZEP7Q3JczSlLKVsF
lJ40OK+iHQ5GlpGZlVfB07tIss3onWJImWuXsQ45O/KCHipO7NTs8/JcWm43SZaAEA1Ey6sG5WeI
osUSbKNmskiJECz1hYn+v1Iq05CnzteE3FN084xp5Uh1sL3PaimcNrh7GkFD1mOjD/42NB0ErFHm
emHPatcd1DcC0OpI0mKnV8fMFRw2zD5E0TOz8ji/3sWQmPVjvbzmy3op+YFqFTTY6FjBehmM93jp
A90Rn2G6FNL1jNgB9d5nEDn9zLywcw5actHIrAjnfN7XBldNWk2u0c8rYWQfqdRyyxt9QQvV5CC9
2XrmuY0YpxkdNZ90dp5HrTeQa6i6RcduKyRW1nNgACNKIuxE4yH6afWfB+kzWGV0sQmkIHHmafw3
SlZCC9fQqDY5i1MxTzF1ajxNPkXUfabckJ8vP+S5xsjG7lYZypmcbS3+daAQ6kz7b+GranCudevZ
c0iNZ4+cKHghWnw5qkDPbYppES8Qaz5bq4qUKxeWVEjUA+8OcVqxe1SjRTUVfO/pxHXsNi2Yp5ju
Ea8pnqIFLKJqczdl+ZCIq3CM++IUVOyG5T5vjYikQQXM+3o9t3WGRDZFcG6z4bRKClg0cNtXPVU4
GMiZ9OzIy+06BhrEG9HivMLvKaxkXK99YDmytoenB3v88rAj7yQwjCjO3pIuH4cv6skgHX+BIYVK
v4UPWEy6CrwB41X8J6ZMgUcvIVMfeHHl0K45wbC/WJWvLADv4c85CpPCazkHgY+N2AnUdjsYOtU7
yhR03zlSq+nSS87rMTiJoFS3rGNgXYbplJKgL2xWFDglmYAxqNAtZp2pgjOrPNJcko1q1zXgZ16W
ry+9ihRcsEzMkEWCyg0P1BhLpqRJ9qNx66olZ2QENVPNKPvEotDiuOK+vn0wY/BD7ciJMafJJJY/
R9ubU9DECrJifMaF/XIHJLRjEwGHKAgNv9TZbBCIZtVfVSpfFsK6Aor0F8xJHX18oB314Xh3z3dQ
JnbSXht9MBebIpNfG89vK6od58MOkr72anJ2gqd9C/GQS3jf6/I0Z424jLcdOYKk989hVtwNIAkr
kLwjambGfB0E0VlQ8rK8jMIzqupgKBOMI7KOE/2tqYyPNfEalKzVL1qX1As+zoh2HNEaOxgYS6Ax
EItROZMixrWcIFNDCIOGIf/5yJDF5QdeQvsWns5YEhYL+bvvDSWmJLGQi3RnrEvsbR28QvyqvA1/
fvpxVJhvOjHS4INvL8//r7lMvxX2L8YD9VRytrvmIcGjP/PNojpuym36IAtwuGgd8POfh13dcj34
Fc8+qGZHVw/GKGVw2sQfHnxr4ocw8TBg5azJJRq+HqGLaMaxF9LmqdTD1jGB1ytLq716FrMA2DKK
FptqYffnoUMd/vnGeWHXvn7GQuiBK7nfGURTuvZo9ofsCryIOceVLtcIWH5yPpNtRLhmcRohLZaD
EI8DKfG/aJ6XMjNu4Qv7lap+v38IguSWM54/uzU29HVvNbAWqQIK4wIJpC1rwYAY0VfFopo8YgEs
7R/ueoJtl6uRnBd80n1gXwGwvbsaHc1jp1w6lSUS5RAiZOXH41BXn2+X9ZPHtS4MFfOPqlvguuoZ
R0vJP281YEBYpROin+EmuMqF6+WvMz0Hfbmg6iRaDwSkjBsWaORjtPURCYimsnIPzYsMy95B0Arx
5exdrKvlGeuhhSY3//9VB2cJmfpmYGD/WJcz8OZTtACfMk5NB7IUu5RD1bqebryuA2Og9GJQU+yl
lrP4l/VNdJ32GM8MfxvkITBhlGSUu5kPmejvR1VofxwRk4ckyzO+Xf6QpiYCMWLe+Ov18VK29PjY
V79d52iM32EvW47ej0YMLgayPRh8WKDhJrzzwKOc2yGJ+mt+ud02fUrwzucS3j1/d3n5Vmdg4AvF
y2TPVVUrk5i5gnTWC1NxUhfiQDrBkesxnC+lJa32diKjoFttDG0Ln7+SrVfTC5kOC7Fnfo1GDXVX
eSDppP1+1mFcvaYFpAEaeD1KmGFtC022DCjfbPvzCbYLc4nc/jycRdszi2JO/ME21E8I0TkNWisZ
YrvItcqJCfVeElSmuzq5byc/BwTKWH0VbAY4r41qzi2Ay0CFf0e0anF8DA6NBIZXOsgucHFi6xpX
PK7kk3MtcYZDRRTIDnUnitAW+YtRX80VmKMb5jJ6/cQ+mhzhmE7feF9KLXzEoFGhYILGf29UNxCf
TgszdZRpV67NyKCvm8vZZMpVmK8U1r+Di2u8VDpaEuexOPPTPckblWuyuwWHGA+n9V/9VexrL78w
B60K8WkWy4vaVjbeNPz44fzEd0Z2q/m3LmP+zI6qDEkxKc4BFdGh2R33GQnWk4gal/Swiu1dVHf4
pv+QtR/uEc2pM01NfzOGLR+Y9tyfaHU3jTGYUev1SEE3F2eMGVdHfguItxNROV3crEZfYk2rkCnG
wizkNhJJKLQsxpjd4q+BZagoLP6r0uFF3DpRSr8+9YO0XjqB1EoPepFaoBuwQ5jMA8acPin/4ILY
/mFfRH0t5Ooo4FF/kp/dbtnlR/KqSBXL1ugiE26HIGjYEUDx7GoR6kGebRv3aBE7mtRLSHI6+4wq
vMdyJls0Qzf6PiYMwbTmuwF2o38bw8d3aOV+syrIV+kBWY59eRc1gu3EwbJNWsE4uXImzOIQ7Rbg
9UBBMQdxwXthTjoX6//UV9ZTyVBTaeNJOOAeh/v5KeHlwRAcDcf3I/0rpHq9MkLEuflfaI1V/4mK
tXzPTfl7+8g1u7uySzMTOiNSEmXdVtXbmo2+HQk1ASuhxMBd7NO0OjSjw+RxnhjvTLGWourNJQTn
1v0A2z8mfon3ZtAhUfM4xl8TMUZ5V5PrfQq9L5m6TC8eDOqJvSznf5gPNxJgCb90QW+65BohxLw4
oNrf0DUBHvcDpPexbCDiTj9AygeRdhth/rFdknn7XRb+iEmek76BABV9SeGEgTDuVOPAyoXl64+k
RsHFITqD96rDWPcOGvZV+MWVDggFQNKF9MYsqPHpkEFZTHJHNcczraryiJdHe5aggvk0dE+UPp+k
Pfj4efgSH+XvhtP039H+erR9E5I7rTAVBeJqUSvy6DZgGTpEX3QID6uYeAJUCfueb/19bAPUwY+4
gb/WH0KLqLjo5lAjChOq25TT44UptA1l5F+lgEFzA4+7b518YBo7IuYhYvcNNNE/jSyVPpRSmZ07
8cFIaZBECQ6oMFXqBpimoROIhZ/rNkJbhCikyySIDBRm8Y1LmrqwihijBKL5qthQlvkFc5GjQpTL
tcOnUNZZ6xvVOGMDj7QpwNIxTDsHkJY0OM1sNpuvPdvuaTvwLPNEO4FISXYeuLSnx6lCUPAemViP
4A2fyfAtLgTyE4ERlT/baWO/w2MUpuoWGzQvuFyW4ao3ozx7mDPWtMmoAEIiMptxbjiqHYytp16u
6UppB/nHM58AfNiyNoVDs4qyOxTwT0EaGOIekEJRlmxpR0FEqiwfv3zWRZO9Mb/qhtv7vUSDC+bu
QN+HipE8H5mGbli7Imxnhbfr2gWAONCs0TtNtor/3mqHXIwF1Hm6N5sX+G8igbs45H2QxBp4Rhoy
aHmafFuKIpFVJZCFGy1ADQf+eeRdJW5uuQAHWEewV5k0Bdb7TmWrQq2ILkGr5Tuosde9g+5Ol8aA
vviooISoE8fdaBvuSb0Vmrp7arQtZA9c/CDHiXq5KGD5HB5fPhclcTNvrLLAC8GfNiaoUvqb4Syj
AyNrSorn/Ubxd390TgteJPOV+oxO7JVcd9au6noNKEn5G32klLsF77WkmHgaZKrya/bIJCKyKSYE
gRjhuAwfScfYqUlVRO6+cEraX8ra6EhraOpH+UfxBiPBJvmooohOUnd9+HLocRQzYIWCANiLCbT7
lPLNxBvEhhuONMaZimdU7jWAfVjqFyEHCkuBBaXtAcF7XbfBIJ5JlnCZKJ9kd26IhpBHMV46zIsW
Hgxt7H+loG5crGO3zel8mToeS7U5VnFc+q3tyx5KBG1bBa0R1yZgLoECEph7oEnlajw9gl6/+VOO
rUOc5CZpDmDbYXPHUOQhZqRJnfC4yvuIkKS98DZD/qSX4nzR2B2gXlppSk31Nnlj612cWM0n0Af6
gWTw3BESetjnuOKPktkz86jkLRBmtTpc6und1T/Roa3zhYzm4PM6bczQwBWYw0tW5blrK52vgDjD
dzEhA36yagpjcVLsWc64QR/lEPPSMPM4zRBiLwNlpW45S78ybfApRZNCx/lcQvsKrz8EDTJimCsz
r/zHtxlVql0/1ZGmmUzG5HnWgu9xQQzrqHLHEPys4vVcKGq4Qe6IX18SBG4zqMnCvYdchb7jysQn
HsNyDreJTCsyvsbXZ0rwnSRhpnblfu4fMWZ7t1SLVo6lygjQrv4Lj7tKDOnEscGUMs/Kcgp2LZBJ
zBqvyudYAl5pCP4COG19U/0mDqT3V0mBoKdrfroOFZOuuVmVSI2eBHx2Ba/SzX09aX8WthClZ/SJ
RLBr/H9lQ2ft5rQ2R0VhXJ9d1HFn1C+O0isX8CprrTK1hlHiR7CIPDTJYkuP1qpw+uAhwxuxRflm
0zELsr+xl/RPyrJ96TuULiyEDAkTGfJekFhfTq5RYyPq2UBthekxflk8+KIJsflTWSXRVivUW+n9
VwcgHBMz3zYDm9erweGlZ7fQZqUNpTixlKKI5wn/cKJSL8+12EJAMV15aC+d4HD1tmf5jGLaIISA
A5bmDCmbTi0+JaZ6UZO5FPLwdxl2OSbI3OreMuGNsZOfNQZV+gF7c5yBDPVSm8Z7W4wEjaa5RnPz
3SKf+qtWclwv3ulu5zRYyT8cdWiQcvjlHUk6ksEDYBWLBA/z2NFvkKDPfOlKNwcIN4vf5Ho22y5G
CRh3ElAg2lLtnrAsiaD/Y6pcpCX9LlHpQ5g+CKrqLadFe+fNjc4ktV7vb/ID+BiF9AIJ5FgP6q5Z
zaoddJMvxzm/G4M01UEbFwZ78/vg+olzsQMQel1Cv8IuafrUegJbrmMTEgIhEalUSC5otwnn+pJ4
UXE/F19pjBJ6XbiEjAgV/fhHg86dthmfNHiNG3THMvX4wPHmU+gH6sEaiRRgi/6XZhXpfSjZTr4o
u8dmnsqZkwyjMf0bgIKIfHzA7d16FWpZvXgCVBt2RjzQS/Bv+aPoN6oAaTNDgqeHWMPvMZBa0qFa
lCoKpwrRfQYBhcYRnvDnMIi+kG1/48rFMTCAUkM70qb4qIhVKMQV/N+5kx15pm2lJAeYupCA+S7d
ao+Bm3bsJVPa+QCVSWzDYyTP44FerofhV/YBILgyynQYXRaiMRgiuvnshAhMWuOs+pImJa6fFOVJ
2w8DT5+gE5AKbLA2uYlBr6zQFjNiFlEpgXFXaur712ZmXj024I2rjy42uICbW6Qvpylo4QDp1wf0
RX89hMuxwnuiIdLLvrNnE+2T1I8/+Hj7/V2Z5WnHdg63VVUnPNfAAbt/3YaT8O3U37xNVc0Ec3N3
BKFBygdzgE7VuF6HFWl7HlpxzhquPFu0GcvHYhD9fhKj51GQJMwbbAgTTlcNfWhzMdK56e3ey/zE
BS69t5dJ4nXtoOfKP0EG/Op0AIkSt689h9c2mlDWBJqKG2cz+RiFolPgPv/DkNsOop7JnGbLBHZO
GrmE6rkOJ3FM0c4+FibWjBb3zggIjVstF/glutfNO1lHm5Zh0vUC/HoTD2RHoWTiaZ1iRyvYBT96
AwaG1Vo8oCz0+ybWA0VnB4OSDVDDga2Juk5xdRIWGDJZZxOt+EPzN41IM2qWlGbCu2aE/Gm85foG
6d7CbDgVMQPuSiA4AHgWtriV2ZIrN+r/aAbhEUW9WEe8iTSe7kMGFb4LVpMrXO3g8jnmm/TomTY5
QkmQeg7GdkOEhRLRaU3KIVALi8gUQlF2gggjzKR4Id5ee3ROCfuuJyB6eXi5Rajp8STGfEbLLiqV
BhtCJrlN6bPBWMpmSfDCjz31zco0dXCxJnY5rV0L1f9I41I2/+kjiOEssU9x1piq5tn3Cpz8/VKh
PPlEqC2hq3BuOZFGykvku7PMZJSsYExZWwAeaumbHwWau/ZVZ/o4LiPWvySB9r8FjPV4A4xlLT9N
9jj9XV9Yp+vaEol3ewB0BCOudG+jeiPkSniZpw1z+twRW1EVrsgjj3ayrbS9SNXi1sOfdNTs6yi1
6fiuBzk43Pczn2AQ79idc7AgTouX7zV1go9qBIuWc677wFJas2PCxcNWvbIpoKdAe5CJnTdRRfpy
CLeoJPnkmCtBteatkDtOo63YWYWj9OriIwCKgdcGOnayjWOzuq/WaobpBWEbGfOWKsZh8GWbcK75
1h5mGDWoOTGlaE7mpgC2aAbj96Bw7eBstqHIsh+142elQ4jpEMlZWnuLTZmGt+e3CYwIHdbctb8g
puAz5pDBoTHY1ANK04C+QtZLFfY/B1016e96lZ/riMGfPgGiiNwvpFaQZ72KZZdQi11TJ8gYELEG
JJld6m+TtBL5s7+DRUFAorlg37GTXNWkCUmJJAJ8JafcoOaMSp/r2W4INCbd7hDyH475khMj8lDV
rsseC8hxLQHONY+9XyPy8Yn1Orh0OGs/I6pyXIL6XuCd6+RRfY7ywlW1Z1bNiWabRWXEzRNbHLUb
qaSZJHUg6gL52jkDEIGRiEy1FpfK8qps26lt1XrjmUiQA0++JYGvG+n2pGgII7JFnkqREXD7b4tu
k0H0U1bZ8txprbw599rYV9Lo7eB+KluZVfSgV0zXdd/GeVOhA4IKZ2C4dQMeaFCS2gyz6S7/Z4vF
l6t3K1jJzi2TQdvaJ7IbFUiP/Ps/FZuefYLiUEyM1B/9oxPScH/2HS/KRBjLUqY2/Z3b7CGFasGp
XU4YzvtqkyOFWeWYCNfs1+eTZA1ORhyGgrL14BFSGCzveLykc+hwT8BXVZ2LX8Ute1btblC9BvnP
MiInwf4vGX0cZ2IR8W7V0YVGh7f80UlTJNSbAd8lfT64m/xnlLLiI0uMQfiMw4DZIQseRQro6O48
J3Lsmu7+1wXsl8m7YPNLEQHk/mXbh1MWJDV6vsvBPqujGR3x8W7u7v5T+y3XBLXyZ9vQHKYkeY5A
zmWd6lrz1OaSEg1CVfTw2gLi1EheLyoj3VFS1sqUcax9QO28t1VOwab9RMvrEBGy1OG7zRu+EzrD
EmQxBe7+ipQREHz3vadveBPC3PFZEJaVchwjzoKp718jV1h3fGZFeyAUl+7nZDSYBuI5S4vyJeRL
kQoKZiAYafwEVncD23TUFAByUufktAKtMlbEq2mIjpG0QpTQG/8UN14t0CHfHdLbruBgBUXzbPJI
ZuhX9Q8S4eF0Y908qJZWnExTDHYTHv/p3twYCDWFSFfj6PoiH+ldpymmDB1coYFrGI1t3qJzl+5y
OEUrBy+J5C8C95F4DKXmaIY1tCa8d8AzBXHJRx4ZyFmKWRf7gITaN31wwT22/s9+2MR7mArsjtoh
LJSYay+N07SBheXAgCh3Bgj2NRAJXKPoJB4k5F1SDRrqgaZxEebkXnEe8pzQb5cAYnsfM/BRaB9m
lF+LAML5N+1lHJNd9doXkLMwvySP/TGoaftjVM2ykOo3a0Ln2esQdtH1fDvMODECnZ7/Mwi/SU1N
M450ESS4B59isaZITLnixBkaaKiVHpbg9YFloScPbkHX3Hu7hpptR287gvKhHCSahwa4HQ+qNbiB
6jjhY7CjSVVRGaJLxN5sMH+rQmz2jjG+4vcxpFlBAjn7n0AXXeUo3gN9qsWXMKs+GKYrpd3RxX/g
IWuLQ0Xb9PntWHW25MPGkX/c9VPF2I8Yx7sbMHmNiPQXD9O+LZO5nG3nEcmCX+GaZlP2XNbWMp6b
tSq3urP5ZrfY/n8ouUYk1YR9zJfRvan5TuOUWhf5QUDH5mS/u0U4/mW227hvNL5VFRjgBXtcUCGM
E/OYPQD/aYAO70zqZdGnwjHRY+CgBok27kF/A7coAnC4JeqdM/ZwGW3mHgiEpDdHOTvyRM7/StRx
d8OBQUZVBmKVV3Hcls66OCbSS+vfO3RFHLfCAyUgsCQIi8UbnsOOD/nM0K5d5MVHLHAmcg51I1bc
rbyLicCl+Odbncvz/ZkGF7h7ErSs4gCfPWaeB94gJtAVBTRwZMj5s9MXfwao/WxxgrG6yJB59T2a
spm4BMfO2x91hhcKebETG1tql0gBtw9hBCD3PGeBtw0I2jyP5JzEH0oeKVWekah2nfMqQyQaJRHA
GBSkb7Ubvsp00DAWWEpU4EWZy43kD5mia4X67NGJu3XUXIAwOeQg5B8tG/ZSiW/NNNe2YrzS8WTF
GPeQU120/8xS7e9/r6UlFaCirt+w58CB17qVZWkiOJ++N5arhzjZtI5YpQwL08ikXhTDzJMvDSyn
SbiXJWKHmyTaWdvDL41WF4e9OSNIX0g55dBr8xvHKw8wdJZTXH3q3FHeKc1cqaCySWoY5bPBUrRJ
/4Nn9XcPYHEvXLAwyD5nYvcP5EOUfNxrJCKV3lEAWc0SLu5iAxrch3hxXAzxRggE9bKcCKfgSSEv
IuT0m2z9pcsfe0cjtsP4Md2R5ZxGBscdmpzQ7HMd0+WxsKJRi1eCrweZnkDFvIw0BWEG+9obROQC
s5EuXeDEQRgBR9w5fcCrTjhQRYFRmaBJnWe3TovtEwKw3zJu0a+TuA5QJLAfo9I3VvEdFfx1HK1L
KrLJQoRithGw0KtJXcRXO+1dkAtLZYo0a80Qw7d1Hxru2bm1ortqyWmik8iTSQ8OFfoRES9RhPkb
Et06i4Vi9jrmDmbFLGqIlv1sSMik2HTUgSkMRmR1x67CKiz60jehTLTm7O7XyhVHKDZaTJZrTtlr
kDg4A5mLNQC0dTMTFCMM+waxPDRctPtzFPHcZOzL/HGjwxqCuLIOV3mPzKXlATAu3ILABZo+OoGP
Bzc84ywdnwFqZf19aUWhPqxHRcgvvKVRhj4XU4MgLHJMKeEowoK2LIbG7PaPAXGYe2YkCSLf5BDH
pjPjBIj6NYtQK60ZMiP7u/Dhzauln7s0j54tkYMFsNBdXJTWLJ1gWC6VM6S0TkzGgjqX5tnJGFgq
z30lwTid/4wAbeGltsYbaFOO+InrcrNJnHBvj7o4zmus8Fy0srkVxxRetE+gG/faENpzR2FOwnM7
rvfq+17N8b+iEYymbvzFb3C4VSSYEF3QCc1spuwDTyiUQnRzLvL/5siV+wA1dprmUD80fmcmeIQv
/9/d/8nAwxyOPj5QH1LJCYNVOnia709hKoAY28exhR6RU1mhNsKmXgy8fnwgsK00e7TYKKSdXamr
WxeIOBbp0q2p1mk1z6AhPwz9akzidf6C6d/9z9bzalVgQT1+gbFWQ8eVS8ZI5OWH9v9Ve5C3GJVp
bKmfvCUVX20KyewwsSXileeU0dTwU0SsHN6TGLHUbBRFIsyLDhAiG+U4M1NhF7mi8PycrKRJmStB
32+jWZw0HGJBoKPU3ip2V/QLTiki2TlhwsbS1qq0tKSq5WLU7uZ5EBpk/Pcj7Gs9Bz4OFn+545x6
yA0e3+73jZoURxq9cCG9JYfOJ5ubJOWU3xwcmw7cMeYWhcU7+KTJBScsbQlSnPZYkhpQFT+VtqMa
zhnxwKLaxXq9VAVSGeEpChuYBTa0xyIDTlDj4Vnsopz6lRwX2j8EkBpT/yOS1z4JpE3XyzJaVNF1
nZeH7+FVe77ECqSrOdFGLe3o5ZQv6hG0vFMEoE7dCX4WPQ7KTU4iLYyQBsH8JUYbKlvq/RI/dtih
nkF0VV0vgO4R0b1IDSDJaS8B82ZGGRxZ400PyX8kk+J+3LmoZBoxOQBiqqUY19JCt9vpORMH4UJK
QbeZnffIcTJjsIKhkFgbE/+z85Gv3chM0USKbq5N++eiv/jsCJihTcCBC2DyjLjklvrQBEoTvEY8
4REMwMtXSl7KEPo6Gx/7Sn0xBSnDbI0guy0UG1O1Xt7KxaHAv7kHu2frconBSCoKEXCJK8htFLG8
ZmAjZs/Y41JakOPHmxSbKPTfeKewVzS+GS0MJ8qZ3H2TG/1dxcdUpGd4/3BPAYyRKB46L+KhNN3X
5uYT6Rci7BxaR9+oc4+KaRwCGtPn5vJ5n9F+pebTrhGL0X3lfW2q+KgkNzAAYErymtTS4w6T0Ll+
hNOZS3wVDNFHfGbADGjw34TlTlq28uGpcRPf2Ox4BEiU3d2LpRqIdPNzw96rtLp1kA1v1l//iV4E
e+E1+wYMHF/iQRC158FcPnxJ1KLDknGtpe8wNqvcDgenucWLxgP0TgiLMD4Oba/Ylaxc6BhqSTsB
goXX40MNujYJ5oRnv0BKptk/ZwnLsJ1VAfK55zNZpPjMjYYhFjAzG8dLh3k/2tQfqG7RDw8Q8B7b
Yq1IXXvd63H6LzQtY/YtzSl8P54ITgGbE5n6oh2z3KnMNpiKXDCLwKx0fsJSevul0sZRip567fkG
KARJq0fxGTBcMRFVUHWLLRu/vi49+qnvzbZradVaebZXqqspnNER57Qud3UDHhwbJNQ+2qyVVekm
TgWMChAaatcX+h0qBLe/E5pKRVTJSEmiD+QKc5QT28NBvI4zAD08icEoZD4aUVTopqleexBygk4j
7VaLmejUDmmnl3o1xSY0Oh2TyyZKd2oEKFTEMfXo/YwuqpZ/YifiMnIZmx6N67ubonPjBDSKhvKB
G87OTew7aA5HTf15ZVvpJIMHfRg+lbpYCYmemfKXBLS8KnTRRclwaV0cAQ0xvBoSDE/gQjY+wv8/
o8oBmXTGtiqQ8SwjwYMNLf6kzVHkgc0DtNrVeIf6hGRvEs4jn2lJ1saqaYANmgKw4zY0Zr5o9sHQ
wVvlEvFxSMXPdCMlI3TFerbs9+Ud3aeR4rup6wvygK7OqZjLe8sp5p1f/criAc76vPgab9n0P+yx
jQEFZ8hhd1tjiT0wOzQ0b2oqbDEabAVDimot8Eg6Xb+preKSbD7bu7UA02cRTMD/f1P5aF0koUdj
XGX+wGorfXSQK6fjW5973qKWXT9Cs/gjt6pu92xFlvwNwYZki5CTqMU/SFJKZEvrJaRr2IAk60Br
N/Psv6GyY1c5sCS49bDZQNry6pdLAWY8UVB2c1Eh4DbYf8pTuTKvLwkRVmxTPtHCogV+NC3zc51S
ZnFWUvn8akJ9UoUTep3qHIfef9X4EkHTCpJTYDJMApP85B4Us3Mm9We4m2rv8Me6pvumAm0NSvYL
FbHLJTvZN9SbRE3u2PK4XyczNFec50xcLz2SL05rE9Fphp/EJkjiFTsXsJaXEbmOnE4Gb3U2WsBS
rQP5P3NxeyCdyNSSamjl+OlqVZeEp4SZfqomsjveBog80axUoXtco6qZa6Ni3lA/Bu7ZKEHiyjqV
KtV5Ts7QKmMTa53uRgAe3TEPWrDo/P5wdk8ZF50kITGSZvzB1S3978zmajAezQlXEBbyovvc8jm8
84UfFkEcdMrnLKtDPTujKLzV+eT2TaFVz+1DAqBqC25L6grfFG2f9REtQN8pbqX0bLqVhF5PHHmt
8zItRaER9Pw9SnSPEjEq4b4xWgYzGkQgfr6IqVD47uSARz/6Kycx7fL/5grQFmri0eO1HVRV4gUH
DbN6+tP1gfIEvj2wTNNfrc2QphQHjZIuIWCVSGSQ73HZvQdBTxppXEp5Rx8VGRg5PvlK8MR1Du9E
n3Rmyqg/xQihBNWrPMCvcmAwbKjfbX97Ih3tyO1n0+GbUiqrr6HGCtUQJ7cAoBxVPX10G9AQND62
pO+zTqgwOExjPqIz4Epek/CABCIpG3Y8QU2RaxRzIprsjI85yZqK97MoODjfM/l/6ng73ldlgZnl
04ZTLnkG+2jBvuZ9UHYEmKM33ddCznEsXQO/Nf9CLXNVkX3HmVbyu3gxHzy1glUrkRlYy4rZha++
zEHp1MEHEes7KeOga9zLooVbFfBEAkYLnH4Rw5ta0u8HQHoOx3QK4TotPbnN4odii8DCFvaOzgvl
nyge0qHnDUXUXvgTLEppuhqH3IDToCKefx/e2U3d0054LUin2J4tagBWdnJ1+VUhD7toPG4H+P7b
gIB7JClUd/CP4fxR4HOwT566TPS0nKEr0U9YAi49hG88TQbeOpe7VuLKMvjTJbGA/HFZJE+SVJ+N
7Oc7OhIdhZZJs+SFT2S/OhlTyxZm7Gmgl6xc7NDleogLbqyrWzF3SqpdwZ9Av6zftsSYBL6/LiTz
CWHnD07WLyOmxU+8Dm8jKgd58XIU2pX5oFXDKwTjWbMBqcZE3u5w5Qqv8Z5GG1Ykb3pMjZ7l2RxB
CfVIhHKqwsMXhegxB0ekeuZ9ViwDO3SULjG6qSua+Orr1fc5Lwl5rQXmvGvfnKECdW/IgZrmC+Zj
ComDogAeAC34oF78DljuNLM3R7bpTG3XHO0Q19d2MiSMMV/gPY4ofgKstgL77ZOa+ZIWKzAqs8du
gBlFYPuqk5dghV19snJSthd7QzNDscY06s6dYVBuiGnGN6JuLtOYFoCXJnBcMUcZm6cMwPujGtvg
u5UjCAQVdND5be9fqmauoPayXj97U6BVHT6BFxrBFolUYJhFGEB7f5la7QGs6XwzkUu8cfMpoG4q
mfl63enoY9fyQ/F8ADAyGImABGQNGu4qNiZHjg/4ukh4zXt9IdZ4Ogm7in463TIEKAZOvneKEClU
nl7MGmhSmGpJCZcLX7hSXeY57HIfTBdvfb1wQAlIykB5pCds1UrAfbXPiTKRgzWI3DBSWQpVcRRc
xa/iZbAi0tUxuBxqZm5fjCBbnC00di3BFPpM5He7C1/dgMw4O6Svkr96R9SidiLwu0YcdHJK+0VR
/cZLl5lGs0+yrlwuzHgobq22RPI1qn+FZ0WyawBkm/KSH7SnUEx/2JcTsl0SLyEVEzE8M217oKn+
BrxQLtZe5k6l5qsm7kmCv6/6qcqjuE/SRjuj96MgXtIxSikmaRVsyKFqn8ZoOUV1K+kFsfdXb8rb
Ji8BK9xwfqztrKvte84L6jrVPVEaZs//Fxvg9vf2PTzUb8gIbzMXRyGKxjoLVa3pgTmnHIvqKzxr
4eIlj+aHWZg0fHU5H73Xq2OT6B365luoZ6/+m6IdTA9vcIGEvzp9eg2+5IUOhScDByDGmj11vjfG
mX94XsgWauuii6VXDy3qJRJIg2Eup9x9nqBd0arl6t6m3V9s/8r4UyxI3TaQBOwL3KXDUbC5x44o
51MIR65q1JC77uFNopJN0mQxTtEhXGGHNm7JomovFnUbzNHb5fdNTQ1sC+v66O5pj0B0N/MJIFkz
svqA3GWjQY3PicfoyHfyq9dLkI4oBKft2rUn6cENqCeD4FtAMr11FogrEFKUnpA8Znjn5dgsKRAX
c1VjZPD54hO8prM9QRVFsDh8ULerPlkQnK3bx2XKFOyxAZOuYNYtenEqHYamOI2he7K9jY+wnyFw
pqfExVvWvdXvngVkYrKmTLBlmhWmA1s181ut/YnD2psfF0xYpQ0+cZVbUR3dVlc2QoymCVIE/Hnm
9eCjZz2Q8Ir3UZgRmOJoNw52cgFipKEExezPs+ePvRwuNKeqNcQtuxYutK0nZkP1HXYUmDvKtuOh
MjHDSylFhB24OmrF8tuZvng32plFn2H+ISNStWuSBLjim055Ocf6uv77Dp23ThKTFKQ16by5Godq
NeNs2yIHtMnbNKals9ZGiwktpUBEZxZHTFL4WWz9kV60fXHo3DjcJ2SFKfdvE5qF94+9KAR4LvM4
nmwaNtVTSTwuT6fT4FvHG+d/hRKhuGVWK08BFi7Ac5v9r8bP37/jRK1zsr2Xsy08OxkCfdWEMS1X
mF32UXbb1F0AFWOIaUiosNMOzE12473Z9LmsJH4JYTILHNNBIgmcSSppI8zLqNEHicoxOGAsdG2j
saCNfalPw6dvlwCBTT6mPjPxmPAgBtmaR+UcneIJ9l2IHc5oUqgZXllXmZKh3ID/NY9AZHsqNkAQ
ChBJibaroY6WBhcl9ji6A0ThJLmxhRHXuVfAE+BuNsAdAQd/PoFZYNx0zSO6VzdxHBp5oP62LhqV
b0LIb49PTzcb1oyd6fEGoJI5vvassxcgpXBqLlE62CsZ8M73RFZv7zR83VpzBRyYEQKx9yGPxema
yx9+LNYRfq6LuGJCOd4jtIp53LLenTirVEOz4aoy9Czz/ASZJgnW738Vo7ZhXvyNAEjsNrcuhaw+
Dqho1JdtoKCLM04rLwAylffbrMbycHq08/Rbv1+usFV5/c4tJLOgpSixIVPWNv9Gp35Vm8YEx8Hr
Qnj+rmOxpEf6vaGlMgeRMsKN4poQdgn6Tim2KChboiqfgwwQMJUlgr1BCwbCMbWKcXRwMXYHUNAx
4ktADg0LkDRY0HC+zCvtlpQdnzXtxnN0yUGYRuPbp0/GAOw8gr+K6PTZAmWYiCzfGX7GLIOQGSiV
H2Dvx2mgW+MTaO7bZqD1VHRA2Gi20anIOaZENOCvX5U6Jt0GYmts8bGgx8+XUb20R/5YrAQoXjek
8HQYzf+vdyFCk1EDV1v6IIR4kGIbbOEzAQKraER/z/fK2wU312hjEM0JVIhiVEJfgEJEzRy+aaWF
84iOuPBPwcMxbmtF7WYbzKkLQ/kWHM03048gjPV6OXFrxB9cVMY4nu+KepjJhLuZfzOBa3imImfe
ffy3pN4XyO2fmGj7OiIC5tB5HpogKJFPFKR12CeZ+MW/yk+xeyHo/pDAyS/Qk8xg4ynWYwxW3X3a
qC9at6yBUxMcNAiCW144jP/uRxR4Z1THR267fnykIVJ1YI/TIVN9o9ewcREjExMQhbJYMjWvV3TW
EqdprPnUY0qVjyvzZRfkBX5hB/NqBCHme24nPwCx17nARkT0YhKcvp8KJ8M/MhmJfGsquTGsXvlc
ekiXAPGWTdnww7u5asidIQT5IMVbV0/Fsj7brHAgAGQq10ynYQeBItvD7+xuo41rgkX76J2ST6l5
RynMh4tvUea3C81BUWyb5he96nH7TMxmgPuv2troRLE8d+tP9v2Hcd6S+vIXzxhzXNlv/5XPD71J
WKgFgKUbXSxgnSpaPwhbqByAleeZw6VMXIuIv7OOOZSzyr215FaPKct/Bu+dzN1w++hChgUMLiHV
FlV5Xos0IWfMX7QOWPUxaxKRJwOs22iGlXAdFCVgrjHDQIaLojuG7kyWLrJ8xRJHDRVrOoOEzWtZ
R8lzPzMSAcZwRRdyhPGmM5SEozMIHAqIiBeNxjortu4CcPavjGV3/Q9DfNqLer4ROeK7FGbNpXMc
t2dY3/GPrveFF0yaFYbQnQKuc/F5iahMGgDSsK2Pdd5lFsRuM0jFkePZgKn8mB13iv7iSbICLYDJ
g9gmXGWxFIraXlnLNSIwHNVkbC4dO+qpxkUP0cKS2xGHaqjOEwhv7fsX0A6nGv7fRVM1UTZYWmXM
feD0iim/vUmFJxbBrqMaHkokMVRYB9vBzRIMtn4ZkVvr5B6udmaCEYRVy+DexU3Z2qY2uAZcJRJC
VN5XSS9eU+XEbCaY434oyRY/ye9VyjqpfJrqBLydKUQ3WBVRxWGAEVfOnBWjkdo0vTx7JyWyJv+9
NqrWaLYTvhd2JN481lFNhD4mMnAVIJ+LdPXU8JFyWcnzSFxQ4v5B5HWZkWA65epYsNNA5kTtosZG
13qlW1Y3FIjvYfWvp9cidNGFJlC5208xEZ59IIGYOODX/plgIHPvGQJJdvm5946Tw+sQeM1syU70
a4t2Ehv0hQWyvKeXEJpoGNtv3k8kaJig3JQQJWCHAxD123c9G3ThIbJHwSw+06NvuBgcK9IqusDQ
dKQVjghe1/XSjKwhpRfqvZOg3ksIu43rT12tzbS7JwJOFjNMjMO6LK2aSE+ir2U6tBiUzBDXhANN
N/nJcpjEB2OUAGy4/e1jaagdLTNlJjjqc80luSLhEti8UuMpdNCXCDsdKu5wGkismvAChgu8MvZy
VVG0yiiOrk0t8SPSWRXSuNq9fugwk0bYgoB9pBTD+dQ/Eavo4E6TrzQYfDEjxavb36mLytY/3IZi
RqAQRxln1DKIv6CcX4G12T/O7hSFTx1dJsFz50CSlpxgWETn7dyPr60zYt4khSNq7spliMwFfWce
at1+argdyjkMdzTiDeedzwrpUECNrbPV6JVAxzmh8kIDVE7pfbk4JyBdaCTcTHArLsVhuh/6G79N
h9kgerMYkS5c9LsOscH0dwUVAJ01fmWTLKg/st7Byr/D34Ktx0wvBbc9xo1n/mc9i9fxHIgA8Qyq
Hr2AqzHJe16b2G3ofwDUAGZuzjMf5hRTCvQNUjt6/S8yXLKa5ueq5mLMwlxk0UxwRYnJJovL68P9
rbRZR7A3jMA+XdZ86HZLZ8jo8aK1QNMpB0imcIJnid0f8Ru6LSNTGkF4+dbYtXzaccf2P30J9PAM
dE3etnb3cieiFPQ9Gn1tevNHSHxTTbt46U0z4iQ9jwhOXmPBZOX+AxVFB+1HuoEo2X3qRIdx/9PE
9WFXHJRXy7zW+eY2ATd1JL3LpMEeQHyxETtqgTZiyUYxc8VtqwSzdh0CVeFQdBtmdmxVZfnTMD55
j7IPIkUNWuGDKqsIQkdFVn4EcZLpVlHfQ8jgdGhICbfhqF83q8Hsuy/jVqgqjwjpoz+547pk3ahG
6gydXgZHYyK78o7iMhhFvLO0cYM1N60p0oWgLKvz9yNWJEwX6hK01rOmXvx6CimmQFb2iQutTInV
fld7OutZjLxZx2Vk3ZHy1pkm2hhZc/k41h67n/cf+5E1zJNpPmW1Kr9ZTZjh5E8iZOH1/f8pp/GV
A6vJfajq0yogV5lhrDB/H0oeQMEMUeeI0T+4dcxY4adoDPP3Y7QgCpnODppkan+b3K1tQNvvp0kF
4K+XGxiYcVh/T1xF0WqrI2fByuP+8cWdnFgZvL9krf/R6PpGLrNTSuUciuTHaY7IzV7byR8oIdsy
y9g4QzlakxqPp6w1QSbazjcFv6u+QM/G9YkB85uazoS5jCGEquOznIO1XlDaPnfYEvFsCp2ahoFm
N1kALDr08hIRmofuK8nXWlPExti8bAqrWhPeKbzPE4cjf/WB8+WbavShZOqBotkudIeOEAG54ZD1
4VxcYKVCi+tvYxL7ft4iCZeP/whXhi8gPGCNRda0cjR2ZuVMRVastYylnNI5+bx3Xh3JlY5e1QUy
ANGQr1rqTQcp7wCflUR7Nyn+/WDN/Yt4s2qb521Tdg7/yy12IDx3ilNH9zSuLpqt3MUyfT+Gpkb5
hK5IwMqOXvHl7C0zkR7BWbR7LrSETSVTcDu3Bb2ws+K0O2nfqPAoBN2DYDwqoFtQ0Mafun+ABQLI
q8XqpVYZMuTzBr0DvEQXFsKOfCO3Lf+vWqUNbcznddOVAunAFqneabNrbDkO0r4Y8Qk+MPFoM/kE
AtRe9uYeOpdCjzXQRj+FEXTh2XwMAlhbwMDen/GQ6tqiQse0GXCCGPbYoJdwcwafghIaVdlM7YJd
DcPTNdUUzJDzmfOFJeY3cu3SnXVry8mxgj4bEJT7Ogi2gqBfiKOHrqDQzVOKHazkpGPJ8/4Qcq3v
jSlGqkSJFUwXTOBQx0rwj1Q9juwh/1W00KX85woFRGHks2Rbc6Eqx+hcHb1G2sQfnIWmvnVy7tSe
BX8T3a3nZ0P20bHWcs7h6bonyX/g/cQ02ui+Zym/mX4wzqrmTs7BY6O3PuAhsqnlb3/rgFnm4E/f
2E4Dpz1vWLMIKNcFVS/qvuL+zw+MaLnqJOgTZ6PJrWSv/bV3xAg7tJ/7XlVP/DVTYJkvpHKzioez
tuzPNqk6whHMTYEc9Pa/nsS7f1y+l+bY8pWufFoGNggz65TnEaHiZU8b22eHKmH/37D5CRFQlPUJ
DD035P23Fo+sTqF7N5DR7yzerF/G1Z0I99ACzTu0+GCEppHoYeweZR/HdNnmiYBC6XFh9pH2lM29
xVrWtGryUMvcNfd+6vry+2BJAQFdQo5Uo4lkx2bcTThEvV+V5AlDw4PxBs+AN3lMlenafGiwxS78
9M1NXI2ci5bWUafOFaPA1z0tp2bFypvbrnMYmVpHYIkvoHF9Hxede2LgZj9FLKrxrUla0ROFqTsX
7X+47dkl//nIXu+e3cdBbjo0n7wU7i4IX96jY/3xocBGYwOmN3GkXVVypQh4tFqHqC/c+9IQY9C9
sSRRwLs5CrS4vu4l6Sf2qW13R0vDv6WnaMew9GcN1JwCnLQVJMXQeR/jlTx9lH/Yn5L4DVTNh7/k
MBbiYyvFdjGPiUc09rll7VnS9gad1jtKrJljGt902zbPIsyoNA+CNgS9IY1Iw8jEDXu1Sek8R6fk
7eptrHfJ9tQXDSQYsU/alODpaI4K2x/3wWgkVLcKGhG7WWXVDSPmab81vChsFkqWVUPv3q0TAdlw
7cbx00dV1ZeBoPH9Jdk06BPz6SV3AoMmAlN2poimAJR97LCB5SwnXYRZA/LJO6rV9IiX6cDhilNy
BfcIzKaLw2VIDiH/3ndX1WNS8GXPZLVJGo3mMO3mvYBWdV6rOpjdp8fq4D3uN3d35h07gOooHy4u
MZDXfqRCMICFyxDRQTd/42a28y5//2yFLkBeZj7zcb7da71Gh59vLURabEFpSXzXivo+catjGTKi
vWDC8FLkY/r9ITHrHIgD5XAmH+G4/uEOzmOnQOaEhj83M03Ts1RT0tm6Wbkr2lBch4GS6lOcXguH
38xdNByV0U2hB+5jlc/AE0xX4ideaKRTwe1g/Acbz9/1GhWSkdz5VZUln8hT+CL68xan+nCh9Bvm
NQuoz/sc8qYoer7jbUTI1ByDajgHRIFEakV+3hrRZFYfOMRPEAg3jUCm/tppXCe2mn942l93wfTq
p8CPy+SgyjSf9NDT44Re2kamqxaArjS+Tp3msG05lC/Twyb5Gp77oHL6DAAnS1Y5StMFgkklE4v3
sjHVaVP+X9FJoE3RJ109Xt8BK8q1mC1uCzqPvqRCDpOrkeL5/byV2Yo4bt/aTn7dgAsQuvGBMx8x
4LUcr0+lLM7YVPlk6yoQxznP9N72Cj+rrDx8oRJ7wnbPRNN2mf4+JNJ1eUJl6h3814OJyAYpjGq/
pGCF29tznhxDFpwb2EI7LDlziwu8FhsuM2aOR0hVjnwlNDzInWmvi233rJP70A3j7K/lt9rfS/iw
S5vMikg7FLpKIq12gqlU6+d6FtHfHXiBZwdZqkhk0rA9bzrtX7dgepfNQxUdzG/Nwm8/KdQABZfd
exnpeMv8iI3+Rolem4rpV9rIz0bk3+9MrKG9RypbR9ChIhfj+yUJ1JAo9CbPxzz+XQev64gaLGLX
TWjgmALLN+g/ItsaOgLHqSacbjh3/rVgqWYQylCIAW6egxSoPtXG/SBypWV7C3bZv3W7ZD9X4d5z
0GwHMyoAxSUUMaYVmLSgrtIa8FFylJmkSTxsdDNYrThoJTFvu+RpxCUVHMEe2v5H3udHp3iBem9z
MlI/wzzPVhF976SBNi0f942puWMF4BC8hrRyyYcw6OEucHgGMwdfrCZ/FqBh3JBNbwgbxDEX9NX5
6UmLprKq+l/uQSGLDEIWsmUwv4jpNZdav+pnsDjFRuom4bwklAflAPhQzKNQ6Bm2VOkC8a0Jhdrs
wirwGDAAxDj1T1jzNF5yfH3EYZ7su1nYBgkhoC/Ej1NjLa3dv0ITWX3uosClbnZCJXmeSm5Ab3LP
CTHELg++TdX0QAXjyIgv8yz0ecoGmDuc8JfB1mlOG6txRWuyCUBeWZduz1OVpSaKLeFLT0vmy3jc
9/VXotvASmihi4Yid6061oEHIwyaJ1e6kJVKsWtV+jZ6//7Q93mrzszwvN3721jvf3PFW6UQMLp2
FRZY+kj49xHrmyTHLGN97e7GOtWQ8g0fXFCCxETXWSkyhl8ouLWGNtqB6S7GRu+mi1OIlXSTht69
JHhtSLbtFD15Hl0neJUOE1HOyjP5Yozuiy9YpQsTwDeQ3RQIuagMVwjWYgIpq51N9dPyHSiHTNXY
lMOd3eiZx3Qfe/3BnoNwU682Nl0fptnOjXNoHJR9XjhuYh4xOMDZIzG1MxDO4qbCJB1C51YuSZ/F
HBbTvk1Kd8pkRcoCLhTcvORE0nXNeyO5X8wcLt0gN82pHzjzLinpIb0GRXftO8KZPuT82UNMy1At
v11eSMyB6JMNcepZuT8lzeSSpoNvpRP5yCgVSAXXUA/5fRfisgq7c67dzKgxXVCj4YB9iLE7YaBl
oB/ELDezrerWb2vO6TRCWfRx+JGt3FzkuLbU5dI6XACdxPnq2QKlrFIKrbDyad4q+LkvGRNYHrno
Dw9EBbd0gClWVKznIMIZav3gWh6P2cUbFDVC/A+qwK2nzaCSs2oYqWvjPlJ9r6UNizdOcLOd4Kki
g3jySL8FoFbrbS3kD5gQL5Qk3NLF7TcSjNWiCfp6gIn5+bXO5F4/w0a8TEEibThAOzT0HrPjQagc
fRNcUFPDs2JemnmRZdyYsIgAlXVhYMgKyaieZVaKtUMB/DIEWn65dZZsW6a0P1a2kSe2HrNUInp7
hhSaeEDZ4gaJGnjoCIr7Gogro6IK3etkKuT/idZy6/c6QEtAVDGK4kqYdXAvFYQOi6JccypSU0Lp
q3Mqsd0FbKXkv5O82VYRXC+p/M08zjhRbcrrTcrzeVTvn6DC42Db8F4PjbF6n02KRLnd+tqcZIcK
AHFMfKf2OId+EZCEFDvGW+rDQ2EUiiEHlF6ZPPH06RtZNdfCRuef8diRei1fXL9diUDnXGqOmMMg
+2GDuciHV5BmAgXlc52vOTsxfofqh89BAovvNTeHhoYRMv8/ACsfAEVxeZrJ32/3gyhvgSWV2D7a
ck0sjBEnww8wqB/taX+xfdZDJVbhbFdlfImrsIjyizJdiLlwb78r4Pf4W0p8fPcwCKInQ95VNnLr
qbk0p6BUIpCZ95njPAE5jTTwGqNm8P9UAh0h2Q6SlZqMslQsGxsPCxuS1E0vCmgMkASsxEayrE3a
oLhZi1DsGLJGJ1hS7sUku/OTyaOtEI5nuxuyMiiMpiIc5bOQ7G4C/re2FJ6XhaL9Kzd3DCQX9Hu3
qfVMJpOwsljoVPQLDuemfspDKZY+/Qu1Gf8l1/rM1LsARzXCKLpdvxZ9O8lskXie0AlmN/XK/K7d
4bCJpK6o93kQpcoLO41R1gXIKa6AifUO23xN04LX7PCyOp4Dulhifg0qVwHYNXOU1PWl2DeRZ0dd
9bhrrbTG02m7yx+TQcfctb88KbvkmZ6pRj7dao/mCFq1R3TB127f5kia0fPmVn35sPtj3EICYSfA
GPaS01D3xiyvruHbWzJGPmj/nfrC5GvkzQpuYzN1r00XmnZfXBalw1q9wFJFB8A6frEtrze1Eiib
wrHworQU3fgw4Q9N44f3RVfYdOldVu6gDB+mbYP2QmG1zZIC+U+ZkhAWTdaRTkxMickF0DrJpuXp
K5y7kY5jeA/5csm6Dj7StyucUG4TPmxKqJEebc/OuyxAv9VFnYpETsQamDIynV4pPoOba3R7YwV8
hh2zaG9hGRv4+x9G+H4jGtwgqcZR1Q7N0shyNIECOF1aC9CbWxJTzqeSeOsBCRIw7B9IkPW0mDgP
Jcwkj6kQNODqt+YMub7VW00KxkksBISAHIBsJ4D1Ev4WeewY1hJVX5b+NfUvWT4VBKawTu4fhI0c
RzvEPZN087BkfPSskDcuYdcCvWCm+H4ti2T1B1g9cth1P9ABYfhJIJS/RtXtk/zBkV4a8z9+etTu
ulVQi0CSXMQtrbVH7AxFt0Ds2h0kqXXROXW/gEdQHdvDdyRf33jaGkly4HXuuv6juKaHPxQuT2+Z
qhWLdR20s9qyP2LlqQCcjfGf0wXamvEfnbBO+zckJOseYGZPu0wrJq50vmzUc1hVsjgGAFEnonJx
6dzkFFGhiYjSbcTIo4TmTMuZdMxS4554EheOVSmBXcwyL5eZp4O3ctPNXX7ZoIteZSKpKSPMXIis
Q7IIIAbW/1v7W6i17xfOt2b5BCwBNer0S1+JQujb9yeTNtLzzBmpYjpFbd9NK9Cr5Cnld3it7mh7
EMrBvS2ZPQcu/hY4k7+CXk/T2k3NsfnFAzsUWvKfxm27mKCw/5QaWHjT1QPE6rs95hErM7q72yVi
tgEgqOFa4ixGUMZv1rnRPzMSxLLCalA4lbswAww0aYu4qm3gA8mqplZHqHNaZhx+P2mWiy18n6V7
E2gQfpNfgScZDg5AZ0NJlmXILMcax8hREYxHfExjFdxxa4dKsd858IDrDamyaBuTLZCstkK5u9ba
CHjwyDnDJp+To/6hUXjoRqvi4wSlhRn6f+kd0pHEUWRHF0os0NNBSib3igPu73M9+QfjmTs8OHGx
Kbnyw2ufs1pkLIPML5br5AbAj1MK5awJDinW2gTJt27epDYh/OzzT3BA5nkCX/P6NuH4IMKLvXLm
ETmeeEnqO6pmVa9bb+jLcioYsGbYfl4ihvengiZvOWykx6e/gZj8wmYfkbcVMCkS6t/x0afzb79/
n8qkAQfougxymcxZp2y9RGFKxz7LL0Em1VMU9+x3lR0AQw+Ngufa3nR7mE003f11PaCltP7pv7Jm
D9r3ecl9fZaFyocE6TjaB/qBOCfGOm66bF1zpR0vkIgixj1GkYdlZGe8v5Rt5ZceI585X6uL11eV
+pw18JnKrOaRWHbIltXj+1PN7mm+cW5rF7OrIfhe2UuD7t7kQTuZpDpLCrXr/gtk/91jXFMboCNQ
Mkj+6O1P8EW61fdtWkBI8LP/GXH629GP7QbNE9u3dipkNxHL7EBAzvAJ3GypqZQmFEjtwD8aDr9d
bOBHgqosGHPlICTfIO+XIWAU5kq9/KCmJrDaYg5yEvEjpBjMbsYPWErrk5eD9hJosaAMX0+RlbWq
oWBJXGWui1V8p4w86zEJVYzyDmFEz9ZR5A0Ke3E0trfrQ7Kws0tHqOTbnHqDNhWGj/06sTn9Sgpb
xmZyxHH6BdWnAEKiUud5Sr8/861O4/7iKdRDMgU5BaMgeB6lfL6iG5xE9a+uKCP5U2Y8TLB1aNl3
06ffc+SdlF8QZCaJa0Vj5wMK+sCWi9O2wY24cac5VBIkPKKpR68Ri0YRJYnbkSwjvxMTWzmgTJZC
WDAT/Gn72oc324QojRImBzaAbchwuMApardwk65Ej0ZnzrJYQWXcbgb6C6kFnz7Gc/y4tRKFbHe2
JjA2mCSC35LqraF9OjWXaVRQUYr5JSRLCZIv9uVqz79OqPXd6Qkusma6Sut3+DNAAewUHoGu58yu
zlgRrz/0vFwSYFSWTrBkHOBYx6Z+s5C1KZI3yhCJoTXxr1onQLHBna8OSO6II8md2tGfitZD5swN
W5PtIeysOZFf75XcwGMDsPQwLyRjTKZSp3gysWi6p51lZQNvXtJ9H8calW2Avl/M7wEFw2SubzjP
sh0BQSIEKDDLxC8p03RnBRXJdBkggqWrHFVS6SsSYZuCNv+edjXysulvxy7QZ3t7Et/YzYDg9RJl
h5pzQCu3WyZE7vHpSlXsHcp5Si0TwHCY0/9QVLROHbnehkzdBsDhzdf0f1686YQB/KZRrrrBr4UO
0eqotit3r3+QQ54WkZeLuzbkIm0TUqx9QCmGV4wpQXCOSOZgFqoyauVocW72Rt2xEdnNQFgeSZTn
dNYB5+CTKGzAozQi7Vck1sqwwPQAcS9nL856omNRTKoyGsa9tCxEMWwII13HpKFcXzwmHIM4digw
EnamWal0ZU2el81rMp1p595OkxBvZ8rBiDjWxyVAm4yswUcYz4yh3BoFJQzEX3jYATC4hkAoLQGo
OMxrvHh5nUUmnNQvo8YkZg92x5eShS0DRkGflePaQbWMCF5kqKk/l/cJCJb8TGE8XJXLSfORA8vZ
qDiVWQAC/oBIvEBLprzo84orPnjcS+Ie7xqMSgQK4KUzV15e+GYiafIqg6xw1VROzWmsu3ouNckQ
Ei5jUi06/F4jA7HlGB6PvBQXVXnyCZQzWv3+p7I58p59odoXH5i3I0NCDE2TObjjTuBpG0EPdGdW
tAWvXZo/VGMK97U3mOc8ypM/s+ECr2fzgszWjkJ6WIVkd1GBpnFIJJRrmUCDmEx9koiuJMSCI2po
vjYhBnmgIENlwGXB0cnyK3ZZXaikCmXOzMNlqJfOsfxbHN8f9VncYQ3KADauZBSY00hTw4haQ1it
SUkG0YqDNcD4cgfftMhnXVcmJLEuQOuhiHpIL8QeaK9247daQd5mOOptfSi3+d36gBHUDjpjF8Y3
wBxa2D+2Yf6ZbBq8aUAky66J0nTC34W2TtR/BLSwe8qitRAotHDutSTJWacXFIp3EiXz1kURb1xF
NdsY3bRLchXMVlpVVrnJG7phNXMe5bvclJ7uztyPa2DzZLz79Nzhdo34NdDchvx2LiI10YTyKALr
k7PGq35QhrtA4t15nltwfk14pmPL0+c79cQu8AZ2eupooUPnbiXAz2IIrckHR1Z9MDqfesau3iG8
a6uIBtTQYcol8EbSMyCOenPSLk2wEmrpo6F5dsh4PaxEaVlf6yXKwA1fyslKfpH8U7XK/K7p6Bcv
LIFAvsj3L5+uk0Uk7sRAa/2ohF53CWPJAFRblN6ndYK8AQF1gY3eUMQMi/ESOEJO6IKaU7OzvOiZ
mGzV3OOOLFg5HB/pf3inMNCkPR7RMN61ZwzQGAg6kYpzJZLIbi0NrSIdKm3yRnRWfF6QPksR4Rks
BWbZjcdcmpTX7hSeDO3P6dFY+6wk5HJDYR5HyVQeuEgeBiKQcvLnCC6mUdWinrzmXWFQdJAN/5BD
uSuFC9yjPvXtOeQgiHiNdxLClLagXagohiB2JWNgQZs8x2vuhnCnb5CoEhrKx4brZvTrNhv/QUcX
JJXaMJXF3c+yznHMvFFnkjPlQOL9Dp6hoGSvy4gBruZnOr405WOqVXLYRIcd2kTA4IRGB9Mu8dT/
pwmRzrhkmK/qukU2ZUopCLHJbOZCRqeBrmjk5/CJQC16w3rHXDt/5kd5/ob0U9qMNXLMTMCNvf/n
0YgK0s55kvXJUCNFEsaE0fP05pgJk7nd3kbD6OnrWhzy8hYxFJeyh5jHk1Krtk6gJpOHFoM4ioyA
IDPWkTx7UBJpxvd4RN8s0W4LsxgepWXQ4q0G2Q5WYUswayD2+1uQnXucq7AsTR+0BETDvJKvr0O1
55VtpUx0jvlvi7/vpwvprAzHXBJYPvM7tVXsZt+s+blfsGHKNiE9aWD2q0ytbw2/itv5ty8Ayl2H
I+1uuR9EBe6BR8kkPfmczZONvaCNSv5yfNtYa2gmjdADgeuyROvyavz9AuetvJssWPuPsaeV77IM
l2dbxIRRpj6RfwjktSh4/UyzrREPhI2pn81E8Sk5qNFJioKOdjo9VQ3LtGMTFSJF0p9gBfdwTHHc
8scqxu9EXjhac0Dr0e5Nk83jtQ3DczhOiWlP1dVnEugm03VUKSh/xW+aUe/0Y574WiXSm8dXfsyB
0gBebJ5f9BXlOwg/djJi8ObAc02PXy23XXdx6VC2N1CY7l8jw9XSdGUFGjnjMp+Wj1xKlzQKrTCA
ungX04NxwNP13e41eolsEUoZJWC566V16h2OIxFMa7o+/GBEaX6RIyxldqBSL/kcUco00s031V1F
/BSc6gPRtSNcvX/pMBbRlDrneJiIujqc5uqPbd6n7PgXt9K88RQfKVaF7PS8dgTmo7c3rl7jzjZK
X599HyBsTupS1YusmvsDR0c7MLtt3phThJMajIbBfH9lcJbUGfm4or38bMyPwLIyjxLofu8StHLK
GnJKhZmogYsd5e+SR0qIEDRrGx2/2jZuTXroAgYPIX6aPy4hp4W62kiplSN0eQIZ3Evm7/hJTW4v
Z2uhMnLkhf40GpwgoYQR/WdvL/stGnt7hj/gLMiBTiMcMDgrzjJGHdnyqogfczZ7A918w65bVMVX
G+4gi36EM+haFmsxaWr5SpvHUrAHgj6I14hn400W5peNOWzxNJ9PUPy1npYKBKCObzf3cgeuW5iN
qesSQOIaL2f902SCsnRI/1dVhG+nTDcEHp78um0Qg3c+Nbk4xgMD1vnQExvaB0FpA/4RKYu5BiDQ
fcn0CYkY+3raT5u/fVW4oR2dYqzEuWTJ1He+o563JLzc+a5ii1YMohTzaC9NU7Y5YzvuYKU/eTEm
N1uAh6vfbDhmhkoLEHvA6UHbSNWTmsY/frrr2bjcEXAT8clqjbtfGuPSOz2Rf+oK0hPi7VRYIHJp
N63laOPKM3Jj3tASoTZgmqzj3rSx90+MONdc0ryJkAvpMblLXhT2y4mv0zVBIuWfKleFq+D6f3oP
DscvklcYV+kfauZTfzv8PuSDTj+rEcxezWtLFtfd8CZ0bs8eABG3nFthgDaopXpDLqwBKbn3IRPl
oibI+TW+++E3DFrPaqL630vAAAiDqYstFP0lU+izdZoiUHGX2WxHN3usJm3zp1hZ3wBOTP7ekMTs
gahv191qn3xvOvPFKZt9wZqh7wcs19LRaeR9Z7AQNyORKCn/nt/gN90Av7FA8LePaPl1ziODbhC8
t9iJWFKX08rVMnsmuBjT/psR2muIcp3CktbWjyr7Tbx8hPgNZYuKB4u4nMqdvDIjdaWtth9L0rNB
LC9p8nGbyptYgD6pLKaa+FvOySgFIByC6F77i7v5z8Vb1/dylHr8SYPU6AKCoXIaGWfToKmrkIqj
Z+Hw7b6VsfKuRVLwUEVQNErPapHDMX8nRRqF6MzVhpVoLyb7WqaeQUsmAZazZpOvpX2GCQQw7K7N
PhBKiJG5amggId1YS5zp3DSUWmeELvYPx/6+F89Acj6BiXEwuQIPbLsaTinks1jBKoboutTFl66K
DNmlweZjEC2B2CvPrONVwvMpzPbXWm+Ip2j/muR8gOpCIrLnrVLy7VqHQtcKGY7vauUO7sTM/XtH
JPXCyGxlO6MSjlcknm3IYM+GMXAAzzxFPmXUcIKWo+HL2GDXdCblDsQjRf4sW40yhf1/Ov1hcuk/
7iAfUzamMk2lg/YRqgQOYJZMihvtJY6nUBEcS2S8dkLHbavq49wKtO0Wu3PfwR+Of2mQvR5wXz0m
ToNJu667terHsJMsalakteHJ0cOA57ylGXXIKIeETPJUyoAHmvH0xrAW9va9cVxVkUbIQG+1hD+x
jDMIJmSLlw8Z6tMl0brcS6zVshK6d8iIFlmuCtdQkUp24QgduCGbbR927jBTqz87DcZ8sTG0aVvA
jGoFYylxhuYlT8JhkxunJuO9Cz1aTSdrjflomNsS/LY5t1xCbafQYqVMMB5/y/zB/PboLjOqHlHR
ciQvwfUFgxmLeHqVdLnx7y7jNpCwNJSJaWAy9h5WxqK9mE4RTf/ZPIXfVR+weNZ7CgsdvejDtG67
QafH0HrmoRhVJxxdKJuo0HHksYOdc1IS3/9lvibvXzpnOj5loS3c/LFSOowODDzTBlcspwr2phsU
eZwv9ujJN2t3Vvooqjdv/7cBLyzUt/tt50tsdRtnotjU+cPYDigQoj7+Y6IJQTBBOebe2LWOWkGv
fPqTWzIWQQDErVV08fSLjfSodSyPy+XN3QgWUZcOA12aCaPdNZaaV1jzYVWd4uKt38MKh/NcTt/l
woQmN1HyRgqZPqFptgTfSTRGSVtgFSxy2lSTZ6US0WQs7cGZpFJtonH9Z4hmdqZ+WpOOm08O3Jkz
1K4fPmSyZ6UVk0RD8smkAponFx+PJt4yrY4QXwRsHZq05vFhpKgy3smC2YZP53wC8ULNy4f8tYd+
QSTjOypaS+Xr5IHuWsOwh1ux051ychDob+SnvO2iaZrGtrxgIcFPyMQ3sueJdUkBOj2tyV99CQ2A
3V8ExOPxzBFQCZqXJvzoGnpf/LvIbo78raZ1+10IFOH/v4mCqjFYyNGYCGCFI2f0HBFfIAJY1/w2
99yJC+0QI1i18pxpZCf1ME+d3dMk4RFvOOzLx94430At/G6cm9B3R79B26bxf73wCEOofIzk0UB6
q7ZN7N06z5RgU1Z5iuUL19Ow+HsgnPXedvfqSpr7IanKMfOwgMgn7w9h1tQIy0WeUJZRw+2tLsov
vcfF6A1v0CmV4HYpCERxwO0zOyAomcrWSzZIaFsDdN1d/46/2FRhSk0URZmoAkpuFxZvMSMwMgIg
aIsrgjPyAszGMt552uOSlsTglmG/YJO3pgVwnJIC541hPPwgIKbLH9gU1oBw8qn5vtxhu97BgSFQ
nd41iYNsHUpB/sNDhvf6pf2W1/E5yISajjUxvBcPM2GJuo6WcWqZn60N+iUMukcxh3kfxDOKE+CD
HIrp/11CEq6JbQvRYI3NcIgLu+EI4fafLdLIrot1dyXu1Nocj1qFewN4eh5ng4hkLUj9dF+6oBFO
Z0/LKDZ6+qW7GeFrcXpeE4YffH9X99kAo2ojv9HeBqSRH8OtCZcNpUW4LkxPXg59Y5VuUFwwJqrs
Fp7lGGQf5R/G9J+lhzch62GULQQO/SVAN0VRkbSBkOU+vzB4zWdvecBOXjl3Hfr5wF183lQVuZG+
12rUuXG2iJiQWTJG2/1NaAIfr3pv+Xqbc7k7evZ1XkHynKnWRf+6eFZEJG8gLsE0GeaUeFRb+8vZ
EYmQIyhHs7NBuqrdPOqOYJtCfsmPMJKn97WcRU48t5IMK03rmiFQEYlK1AE3LqmMsB/e88eE3JFV
ibVyNCGnQCZqDecKqFJtl1isCltxygUAohAfb3D3VygZdrgRVzL0fcsZX5XBu5UYvnYyFCpKEDGt
Vya4EBTL4l15UYM++8DPoDc6z1gl1K9CVJCGmzvgqm5W2/O6YSN5ArDqHzkf7+PTRg1EVLMUxJ/a
iVjTUbfRXCEdRxnSgSJ/nLb/6HrEwthFBOA8MfPOVQGUK9FSdKi/gefrmO3GWgB9DOmWy6xC79Mf
s1P9RgFCV+qtNORYVEKGromyCzsRQrVkPDACt4leg2oUeOnG46i+jSbt27RZr5OLT6N68XLO3Su2
sBQDJH2oKHt7PbvQHfquBsJvlgGemk6r5UlN0uJunQuksO90N5gTynry1OO4Qyz7XfOzqixnb2gy
yPUwv+jTxkG3T8ZWnUXIoZGqGMs4ytFUysjom3EEEdMAcxsCtJ/gCDJTD/FkL6pIpvMzCoFY6XJt
6JA6XivLKtJBphaw+1mJ1e7AeP/bNQ8MDumjk3H7/ifjo+4AoSyx+jFJDBGIW6PenT+hlbNcCGo1
l/enYdjKCaaZ7QmspAQEGtOHZUYV5D973B2Xx9n2ZjyYIMO/64ZuyyYfJ4QndYbVBCWxxhMo3MP5
fvgRRMZt0t+320gxLQQYEuSekVU0t/uNNRE4n/ZffOwgR/w5jCKBr9YkI19s0RFMgHi2wKjLvt7n
Gt/R+R8F+9DRB8tgV6Ejw7VRY/kVIg0nxmkm3dSuD4a5dJnILDqB309HNpQw5m0DqYiZ7ZNrPUgW
uCrZFm2p1kM4HTIxAPhU1bP+s0W7JqDos1dpWpsQSqpemrhhGidJ++2I2DbobvNCd8fbJGMijZjU
DmCSz/6Pm/Yw/tCt2Wjs8rOAvlJxE2Gnv4si/EWevMKr+AkP61IdLO58Ajk5WyTf6OUdeqwE2G3y
1sNOgmkcYcux8gILZGZ/qA1T1GnlbVDdsWkg3XywEpbtaGCHh7hhsoDZtec18lk68dHv2jsKkuCJ
V+VD3Hgo4c8CVQiK66TQiWoac2SApojAcj7j3R1sK4/e18OPsUX/mulPricYisrddsF7HC9E/Ptq
afYYO/1vJS4KGQmlQ3i/r9nSSVhXxFczVpDrza6VLtu2DGEsQQtucpqHMj8JX+yAAYbFCKJ6P6kx
TgJh8qigm1l8tuAIT5Vf51G2+kBHN/g/46oQyxGkaSjXX+tJ/a2UTJLNamUs3WPmUGPVejFNA3DR
RY9JHWWPVdEQQ3F2cU2slrKZSErx2AQM24YaneJwfUIg6z4Ohur4vfWiZy6NRdxMbj5SuGNO++L6
YXI6qzSrluKFIdNdHMj1et/v+Rqxe+x8Np5/NedA6m49LTXB1WzvhhzpnL7Zz9G0kdCx8rlUIUmA
vrOkGJpw/44ilkexz32Inaq0qvws/6Rk7vTlKko6/42mTZD3xwhjm0nN63NBFe+V0LLX4tsJEL47
yomQiJIGmQPMVgtiWCaIJJuUF8/StVWiP3Hdmz5NknsB/97zfdRbybD6+gSzXVYQzXV9e7Wvwmlp
US0Ab0QQfOKrxE14ZgGyAW4Z5aLFu+G+cEQinn/n1TKql14ZeixKsSXNNZAw272JFCfhc6XwoUif
ZuPcOdlVyXOT0d+n5SdeVvRBKuAMypdXCVRJJ3/b5D+OEcZewuFBitjvVor4d/RI7vfe2Ef08AFB
4piAEIyoIzeS3hpLga0LFGO+fwoHDP9YZpM8ZoeofiZLNdYWG45EOTZloqtVgP/oLn1mQ5aVCTLy
vuzbZel+nLQv1yUwAQFGAfkrcmO4WCaz50Ece7oJSmuiYgmubvpmhyvynGxCo0Jt1rSc+XC/3CLF
LxcZwshZ1C1ap4aKT/QNUt8me5fOleezBdODWeysLM3AnOGXH+OvkXByF0nhtvlvX0iJZk/ate6o
VcTwxQsiqTIFpRmFhPHMo5QJzQUDfyfCCkhOOypFp3K/mGf6Egvem5gbsCaUmQaYFm/cjBPH54kd
5xddS3l3bktafrHvOdzK4X/wH8qyNZ4Y3F1/KIs8e/TgYUix5Ohyc9t69W/lI1fptGFASUOOM80c
giHzZbxCQ6A7spvSChNspcNSj9N9GEK1BUxI40zj2Q/9ewyVNvsFGklrn/3mHgMjq+jfIxmFPVsd
ehK8Az9ePnJQwIeUhCT3LZKdTU0jAFFBTKqcKIAlZJjePuPIezwyIe4+6xaL/ir8/Matbzt+S780
spHV5bNcKSKJWffp2xR/fA8Y6U3c1WeOS/5hXwKBGVnMfF0kpkCLdm1ETAjHqvzacqphwvar43Lk
KQNTvGrvdrR4GzHcD4GEIHJG/UE7mWL7Ea/MgBQko3sxYDfXWpdQSmjtY15DKEAvIOVDXzVTeur3
lCImAO748PbSA1OzOXRq4vzsXiOqM4xZQ2xBkiiPI12ffz1Rux05YLNAd7Y7UcYpvvfc3h+Qwyjd
yTaRSgbh9+ojQZEINkpaABQnRBczzkS7IppQOsvdIuoO6TqikWrT5pyhQr1uSmHvv0gO4B8CnqE0
fFyC7YUx+w7sbDm1Pq6GBD7+1cwQYMy2PpP3cpYKUO2MJmvuCmo6WbIRCioAliXpvBpAzg3J7j5J
7DnsxQ8a+vOT6frKr/A4XZ2EWGIv1GqIQ89mX91WeqDa2BoFnhHGSedMNt2x2GP2tfd4+6AddErW
TWVeTG6gOBzOZxSZeO/ChtqDxQSmHoRCRmxq6kyNxdnJG1lad4Xasy5wxMryDVsTaTm9MQM3Xfvo
7pXnQUC1J0etCvT5HhlmsYl+mRPjQjh+z4EdI5BOEaBghHuucNNMu6xYnI8a1g3Fpb9Yos1iwfmr
ruHwLLNFD/JN+xx5oUcOq3zzWHKDwkXaG+EDFLPH4qjrv3o+wsDFYRNOPeglty4FLO7INIYg4fWC
6yGSFRHH7qDpn2lVacpioAoTB9ydBUsAR2ClcodLvqEAzKmp1CyU0ojjDfXaSdm0rWQt+x4/j+ec
NNFTa3nNKyN8dsazPTS0XhngrTNCdS/iw9Wx9jj9s0SHpxmRmRgoSemACIRa9COGXiiPu0Efj4xb
m/bbuwyRZkfMvNNqKWQ6dRL6gInKyUUm+Q6Owk83qWB5Fq6OBJbC1l4fMIc/XRfWN7GAFo9w0MUd
gnWbZrHFqKEuVl679F/rLinzoOwlrWoRC/zmR/OjqrQGyy3C+p6CWBxqEJmksaRmypukXFv/osgu
6jjUzeZv5XPUE7zO2Cwj9vThBIMJyUBgaiWEahXWvNR8It1KV9UZxb23m1XD+KJd5A9mR8S54Drk
UYUguYACrs/+kAx1jnrDvm1azFHHWt5MtpcfcUz1NYCc/aiwdNRcpM3NCZgA/AOongIx0FecIVjQ
N9rJOKY4X20uaye0Fi6Xk5uBiuAwyEs27X6rNwl4xC4uV357RVdDXBU7XPehOaSLdZKYyPamfPSv
Z16OZSnJuxg4nxkgvqan6KKaf9OUk/dKyR127PECINzT+xBttAdDxPt00Yh+sm4jdVAgBLU3PME1
l/ZWyQC6O3ph9ozZplqfaM5dvNjT4Zu5vEFjVdvAJhePtV96RMDrLrY+5OofoC455i+CsRQG2By7
5Y5Q3cPIgtbJ4xWDdbpiN7bEnp9WcYvNvReef3KyXRZF2ebjX3JJ0t5kvy3+u+2liRk61BdGZJwh
wjJO6h5wyeFQA8uNdw0xg0DeItR1WcTBRPoaJXKPLWO41QmzUj6qkMUMcMk0uoXMU2fHU/KkhPmN
0G0bMJrGMJKRFkVOMBVkSYSv+dn9y+7PLVqTcApQzRDedlaT+jZv1Od5TzgJKv9c62IwCCCj4IS5
LPM4MRM7ivscC01hko3Fd+aAo73nIc6qOhowwstzLWFZbO281QfWESugsebo7WynCAfCm8npGGFC
01fY0CzBAmK5/23pjL3fKlzPBLAQyLPbp9OfldTtfFSgESIt0p7R3I+AbtHMlmZZWWxEqLpX9uUQ
hoX1UnBfsTky3AEjR38QM/29VUANSOTr0kVKUySPDfYzAKOJJVKGbrCgkAEkO3i/mFicwkBdfUFj
5nVaKJ1yHXAJIWj5KirhI9veHYNzsKah6bNfqldNimRxEZyGQ0wH/6IfktVaGMBZKTWOSBQF0BYv
KUDVIIaoFmGLNJQ6g8PM0av4xPZhr6uwTm0HkBoNDKNVRdtRB9SFqqITPsy/gcG2DwYtqKmg5l/R
p7dVQlzl/EwWyGXthr9xTJ2/7F6ahQG6yq95EdoJzk3PhpuWMcxCE0GIEv/3NyKkZL9UNWatfcAo
rOcxXzlUkv1OAJR7ApFlnOVcKSqrwLslYjMRUPQYrU3L36jUtPf6yVZlW2G6ipSX0W/NkieKCBKU
ijHpRwxl1X3/ZoUEzeVZTmPqFWMi5dd6xHqdDrN12nRmOOnf7yVhuQc1veuTfPNhnXcYuJTT0YqH
UslWpaCORv8Wc/VD+gpVlVPblQhk5UUpRRRWLHs41cFdoTV5bgGErDuM0HSjKcDEkBz0Ecd3BODT
ZHqKhT+Eq0/AGclJQA5S4xkFLeg7AwNgnVYGWD2d9DisYZUqEI9AP8Mtv7btPmP/mW2jeQ+q93EN
feGMDXasueLK/L5ffkDbh+IHP7JWgePxOmYUSsKonXO5O5eRvNSpr16O0a6zlrCrAMYSAkzpKnAE
AQjEo9L8JYhlAVzqBmh2UwA2fjp6pFAWX4s7znyV8tkYQ/X/YFpilZ0LUA/k7xq/o/bj+g+lFyb8
bsIeFR+9ToikVe5SoDJ7Zq7dlahSRJ4WWff0BhmFC1BanM95Ue5t/2dXAE9n2hJE2iryv8Ms/u67
OfGKjuwvokExOfvK5nUkGuhl3E4LgQQ34gqB7rZYyj2FN1fLMoVj1B+RLiSfxkS+nNAuh+m1/3K8
pS0nDyhuHYBV5eaMxnB/wIKAiYq/liMt8wQ9h5KRe+Nj8UV8DS7SU+gR/t6P0NjfKnz6tMphOtNV
0qCi+qiYAdAGm2mEFwqqsnvvO94VhptldO9SMQ8d1+Ir9fao5ym685/8sme/JhnqlpujvFsbK5hO
7ySXHGQKA1itiBNyhT+8jcBUtz48W2ln5rfTqOnp0Jzq7OlpvnBodZoNTbNzajlcC1uJ0KtacE9x
aMRCk0m6OfslA725KchBUBiPvC7ODtFuH/eShjXJ7LTu2onkEc4icNqUJwlpt/beaCYFbHkqzxHY
csDehRTQ6dV/mS8436fD1o66jTOxBvkUF6TE8ycGoJS5oo5z4yACK8s4HEhQ2Hzl0zvnvc2LJS66
fUzyu5kFrjNcS6gTpD3Pty8uCH7HARbTt64zxlVXz6/88AjO1sb5rVj0wpQPMagaeVXsAvKyrUX5
xifAT4WPknyCvMJdlVxxcH2BrD5Tck+NW2TCCzSxqO6OCh9U6qTUee/Rf8p84AFO6s36/HOupHAN
TtjQ0Ggc5fyReJDK4eZmVE4wt6iw5LGMy9RuKDKzCyAfgSStv2sVHZ6hcPUFaRyPqgXUUpclLFoA
FJl4J9s1x3AnxY60+KgDCQcdsyDh3KtBhX02Z4DXBC2mbu6Sw8CfWK47sIRN3na9aWKAZDnUW8T3
4vZmMGZ0YXrSmxDt9X3T9pchTCJL1dZYcgt5+vQYqPhmZsamKYRL5+sDcXr2idHodDHv/x2/FzA9
DPDTYUTHYGKNwbt6Q7MSKlBnQYdkgg8JC09lDuACTGDs7t+SkWCEuZ3E7/LspB+WApPuQiHhV/42
rbciuoKB3xPWqxNPKYQE8U8DxkMqo1lif3l9A06/jKxtF5Zv5QNZv7zi/XHQ5MvcB9QvOFw/9j+0
nOPOqgmh7km+wcN4Lrpu/jnIeCaVGoG5zEFmsFMNhMNv5aOPNHRXHalJKZSVsal26TfTY6cWlJXY
SZSfRMkiSKu2efkSyRwkgZCrjB2DVjSk5IvapiCsIZwl8zcTvZTxq3DGVwt315G3yaaHUE2+xif7
gH9zZ+y5IonqvbuzpgnqZgI5KU7nMKuuyZdDTORC2zQJgEd06pk0OW2wIMe8IUAilYIkISCD/Zbz
71MgFPGA207h3SagKgOnoJ3WJxq29Qj8mepR8aAgL5hzRKu0sBcox7ZYGumGNER6ls4rgiy9DnzQ
2COxwITC4tnGrjEGu0htA7r1Y/mcs5mBy5lInobAByicOC9AYChjwrEoaqNMyH28mEnXdWCv9euZ
oe9QDAwwjPNgoa4xHFsd76NNGbiLETIwVlexty0CkMASdgH+oEeSfcHrTVSanUPzlYgZ5reJuGH1
HDGOJ/8Gbv5DJxgPy/P8yj7BRx/Q0oMWu0Et1v5BxBOV/C2EaLBUVoWBg9pDRNZr04CwCwAWO9aA
gUWhh0XaJouoQajFGKTFGeYsicq2752p3xsZsLJ2y7NF9YLlQkdMskH9Soy7mGeTkpmqW6Krwvj6
0CaBtMWVsrlhvzFRFNxZkqFH+gAoJEFTEPB6Wr0ZQgc2p2k0lYcgCCz1pbLS0T9xyjpBSJpWm0z8
Oq4PuoobxaI5hWuPjsmjmeGRMg05HdW+rhBIMFxK0eoJSpIKVZ6aKLOFV6zRay8LsMrMBbQ0VRVx
xmQeqEo9QA9QNnjPlnfpHea3tYpBCJwR3kPVECyS8gZGQOfa66438j5f29dQAeV1/HEtcwG1xaJa
0z33Hu0OiS7Ka0ptpCbWFY+jvUudLuOpGhxGrvZS+lWzZ+lRP3UXWomLpOiuQ4sQbDmKXOUVkRwx
9nsRgVAgRVYCWRJCTAhhhDuLbi53MUJ1JXAR1//46TGrhwbGJnUB0MdJugIc9XZt0JkOiahWmuLE
MNknYwug5Gi0eOmeJWUCSLraJfh9hRBVtFAwlnIYxGs3GNnHKm5qwKChmzO48GQHtdHwyFoGz+v6
fMbqRA9uWr3Dl/dSqihMmBd4/G5jM/yH9O09oWsf0Z7TkNUV5etMDBmiiPzpU9fl9UY+9Prp6iSP
A6WJei2glXBPhTC9VNks86/YBTxsWu1wqYQfgkqH9In2lBoKshJ8r9Ky3bfTZieKDcspyzqvXq1m
PoFh9P3NBNvI2KoT2dnC+zP7vJVk1Rmufz3Ykb11vfQCegxwFF3mswADRw13fWFOrRWAgoRAECh4
asifyDBF24YM+oba//dAf3hT/cZGzTaeVUKm/Agq22Xt38Lbs95AghKT+s1/OPzw8CQvjae84FpF
6QB7dvIEDwZW5KV4fULGCsh/U5SBEpIYE4R1PUKANc8anaz/weQ6iw7wq61pXS89E4gQ4aSLXYDT
MBXgmGuzaMRWXKzBRn77AsdIvVnsmN8F/awmmW4u/S+jmz1a2S/aaQpGO1Id5vJ+mM0tzDUibs0A
Mlk7OxB4YUtBp5YqIUCFFMXf6sz4U+MxwWMdLh+LnAImnr5QMINK0qNkh0knDtTUF3gw/9/FrUdR
fNgdlseBmLIIOSM2RW0D30HsY70qxMFn5uiY84WhdnrCxA6c3NVmubuzeIHXoWrClsjDMvd1Ck5t
z8rqWuBt61W1A2B08D8z7+foIpz3FWes+RRz330c/5bKa59VTAxx0HoHOT66bGvyFIp61uYh0vNc
JFGf6BRBl/AL5nWSsa7K+d7Mn65zv6wWC4MA7a+hE5SfhhvHZ7Ued33qpAMDyGOienXByllulE2d
OrOvM/qEtDO0IihWg54v23Tr5iuUOkEEWfpqGFDRzorBy2UaBNYDcQNjveSQVhEXHT9evnFTUi3k
TqUVyaydUjvSl6fJb4M+S/UWIVGrOAMPPMUANYUGAasg8jwBhMk6mx2PLd+dHmwEME01xq7ueoBm
Kj5Ii8dEg/5rbJbZ6mA695VNN21/snJ9R67AKWTOwjrdSRwjCkggOl50iwMFEIvGWBi1OpUqIUZH
YkBkB3PnC0bH14Fe/0OB/2JVI4u9PFmRr9Qd3SMmv4d3Gkir9RXpgxBGt+yGsTkX2TOVA51FyDR9
/rW0Q8pC8PyzOSy/Pz6gUFzxq0CL/5eajg1hf8Jb6dxnEMERS+zvnmh/0YGbljrs7NP/OZWuHlkJ
dq5lWuA4qqIziDPSlQKu+3lXgd69G2rl0xwvUlvYUwwFApSkPt8VQlq7YqafBvTw+HZUYFiYdZ6O
0vOqjfGN+D5MshnOzJHWawrSsk+v6g8VQ17uG3yLHssMz5ZmHfaTGPijE3mU7sPkUn2koIkTThg9
0uDtPAseg2oYpCIJUVWQPr/elO81jKfUDB5+1zLV+KJXtSAaafTxBy+fj83+z0sfLGQKBQxjJQLF
S0zKKVQgOttoR6sH1NK/TsnwA1+jml+NAI/6/sweKVcQjXAi8SVmg+GGvlBAnAKFEDNai1BDGt7u
gdH14uV/HddAZvcZhuUhjr4TAEcQbmJg6M0MkFRtYSs1+vLFpJ4iJ4F47pTYtfC+DvbzTxURiJh6
ItJ+tuhKpxoIcYV0F100FaTam5muONMenO+5gUxH1c0BbM5Jv+MnPOstPTeOEB42qHWRXuj8JOU1
U+LwvRIzFPeoTTRvCIhIDzOWHDpbKzxh1SmISaDEDCCeoVIYNAryml9bsbuBjTmkRQHd1cV0nBG1
u/wbXcOsDY1Dw4Sqx6cJIQURtWPMNA4tjgW7bSkjrwp0ERImCRQK8Lyx+mtHRPIeXCT7MOlDF0+8
EXNyXhll7vxOnVLjvbyJWsr5uZ5PuqbdnCLsfHYtmY0zh+nNnfSel4B+ErCET/6u9EYU+mTnb3HX
bLe/qQc21i5XIHivF9kvMxxFQSJsApuYuQe0KbNxxHo/6AxTXxqdcJa4f4qz8zwRDa3CcvTEI5I0
wC9Od1Z4pKL2Inetb/kvVjUSIqC3tkGY0v24gxW4MMNTKdj+izvX118VfdnlJYiMvXZgAfWf5TrS
hRJ5SSCYo5nB7Rs92ki4n4Y6UQcj8DAbZCjlWt6YKxEPYGEl2NgyL0vi7Ku/EOKqrYcyVR6QzDUG
Wf9fQDgHqra7d0u4PxfThteDhEFrW49K8qVxVQugZgkODzn8+UjliYUkLGfuFoDMRh4s6UwNdiwu
9KGBnZpG5HB3VqUMbw3CMSkSw0Mixfi9MgxWMhs63i6XtdlgP4Wl/1UMuyaovBPtrjNdgaqWie8+
nSxzueZpjjDfvxAKQpkVDQgvii47DPF0ngwqeKoX/+QazUmWJLnEN2VsJbYjU0EDWDvidHko+092
kWsjr4enJPip1NsKyPU/oWZ/YBdICryt5P4seDWajN3bMOn8KkatoJixyO5LRpFKhhET6fkdgdvI
hgDD8EAskrM+tod8qK47lYe5m/3XBIOaqtfzl0ojvQA0GOXfh7tKc8Xj2nJ2nQrncyLEDbjLf6HG
TNqtDHSb66mHeFiFKz3AVD7iUH6gZ0gIqfvX1PnfZPe9MrMdiMUd7rk+NxDoNE67eYlyufuYErfy
Q5Zt9ZQN66UoXaa3pWSreBAF/t1g+2mwXPoXH/Q7dNS6dsmQZMVgjojeDmVz7mZzfwZ8ruSgMu4i
kZzZRNQeTkUXQJJvv7a2lRFktC/SGD+Wcnz6MS/nXbTItk0nODjhr23h2NRAygN3ZdEbl6Bbw73/
n/Beq/IW3XV6eOu+yp/yHusHbReFMUJnUWzyL7VBnDxbVYsxBdpObBgDRhER+r4i0WFE1bXD5WdV
h1X/ZCDIxpk3VdJZdjU9wRgkEFCUElLHEicJjlwlNYH9qFFs+mYShBzZYXBfOGQ0kmSndOEU8dWZ
UG58HtQC4RzTcCNve9jP/1oGtI7vlJAY2XEkgJSceFmuZT0TB0lWucFtwaeyElQGmPZPrjC0g0P+
hgx/CcYGGNY3RBGsXB6HjblKaLd7uof0pYHDztd3ryZi16RjXwJHcalyB2W34rMRsaqrLTfGb0yw
9Otqy5I3KlIn/xXXTAoMVaPceeLxjc+zq1iU2VAzySI8RV4ppzAsExgT1YJJ2d1Oqbc4TQGRUJNS
DbWFb5xYT0ZA7nn1DT4RMKkyp0LStFlSfiuaxrvl8A5p47WybvHxNIZaLFX6AThPsYUoi5fAQWZe
bJEAnIsYBQs8OKfjeNxkCPW9qwM7B2rIuwmWgEzpFc2d3LVtSzeJDpMkmix24EXHCOZu+TF2mqlF
843m/j9Wno0rYML2DpkJV7lLbSLvtXm9R76wdjEGUb9h6EeW3jMWuZk4cUMb+i7yGdSNhd8X1x7n
jtW1ThDxHCXyd7lpUygOzyNJhPRk/MWuhK0d6fU5wwvfU85Wyko9kw3nyiIxn1RVI9/KCV6dmlgl
P7Ah+leUOcaHJyl0CDJ/szGU4l2oPwi00zlbd/xXBGyX2ly3pE/S2RueFu9fOD65HgyBYFFqeg4/
Vr7fViyYmFAJzTv2m65pnNFoVwIrfX4okgSyrbvsM4pORLxkdaikOgHfZX2+QsmMwjSa39H9FrCr
TIH7/3PVzifG8dmPgjlmCkBMHEYAyLoX9wrmZ5s5VpSXgapbtenPaonCTBXL1Lvabr9p+1Z6BB3G
rizXUACGCPeSbeWW02xWwEMtROvGUTNjjvbiRKgoy0/r56WuPiVM4eFPocVulpTAJ5CjWfyswq5w
4fheFKG7uFGQzbMrlY4nfaIyD/NTD4YgIeeWMnpVKXeZGDvhu3LVTS5yaaYj2TMBKkMLcuI3YatP
yefAo9tyXcSAXjul1+ybkVPWtZ+OXOE4eOq+POYkMiKUiqYA6qnj0biOY5NF9aRdrE+Rk4mv/9B9
H9AsZCaMqgBeh8ErecqxSaC9QAb5XBqVgq85lcWku0cf/8I1aNBrN9nAWQPQVun3YftFqrF8nYPo
hvj3DsmCvDH6E/bSSba+EsBPbl2jBNP9AgUqZJlNujdlnGndKfzpHqQjCDzNnnBbtReqRmaUvfkk
571sM1Y2PwVVRuA/a6ofn8kTD3QjLH4ZfixnvGSHjwm7GvYX/glbVwgUk8LLzBrZMM/skk546V2j
4iVFL5HD5+dHVsAmNK8PhtZT32usb7fzGJUUeKt+5t/otl0ECTWDWTMFtBYBVYtZoxR9nF8qISvB
3v67RlPNGoMeCdlLQoC93rk9/sKLB/rdl0Mo0Y3NEWQEVrUf+rKCDmiD1SUrbrm4UyO6yTiS7Zu7
Y2Dn9kK5rVkzGL03DycsHeXezEs/g7bTtoLWx8jmFJpns974V1HRYqUtdjZfSu/f+xmRTVnjQIEs
L0xlll59YSwCxdsb5gQqto70VMk1VexYBVl1r34RNXpVKA1ZyKlJxUDKoov1/I7FV27BolCVYhDm
/gZisE7U23oJFut+yHVNZo2DRINtxLF3mZvlGAjcc+TU0eCkAwHRiXSWZsivWFdO0Ina3WLnt+8b
jEqCP4u6lv88FQmqkg4dmOUxIe+b1dlcRbPDMZ12FMNHSZeid562mw1CzMJIQxxMN2PioDvh0KRO
VPzyPW0AtvtPNmLPGW0XTudtcMG+6NYVOqSxFtpjLeOkTL5huM1hABOgW2WMjeou2b+qyiMDf4Bo
Lik6OjDnPt5Hiuowj28jkak24+6WuFUzXyM1n1esZDCdP8ZQNcGDMoXqOtGhOh/+LVcLKHnmCwY+
73ac2tu4D82RqpWZRnu7JUO6NagKebbhsSSanlxw1r0iBf3POK8+7Ga6FjBMXyblpeai20Lr6nQi
1/2Se578K8CIPz0s3UyXw3iprMru4RaWcJWEx/U0eYG2Zmvxxm/6JI2MuZXQxrerlMIeKKz7tnOb
JJviYgbqyl9Jd6GEe2hbIhmipk2+hdqXjSrgs7PPslqPaQNA0x95hMO0PUOdWjV7wuqb45sKzy63
828AIM6fvZFSph09qqc0q3bidpJPjkm4gwyTGiDpyiNRUMXkLKd4z3Q+8RqyiPrNeY37O0B91mh7
hvkW74BT9BmbsVPxMgpQfqVc9YT3jp59W6cA78Vh02y5jRn7/1CqwBBfmdS9z0uYudhdlDl5nCui
yWNLqNMrCFto4KdtkagCh3ezJ0fHU7mDfj17BlNcakYP+j/+B85/sTgcQ4Jig5l75GFAtGkfMo+u
bgeC5uBIMcwN7PEr2feRK3O9LOzzm2bMMxRtHj8pHUbKJXajDfQqGuR2UVqdWrumsHDZ8R1j2PRR
niKaWcTosf9FfrToh+TgiAOq8LK8UYXt9K5Jzg+S170c6ASobcJIXSiGXNVuzsDQDTHGm0lrKurF
Xk/6zMAMMQ1caaAJ8oEbeb6Jd7/7cbO4kpfp8S3Go6MRfks4A0BPQ3IhUBM7Y9QfGSSQ5nUEjDy5
55J5GeDAb4CtCEvLyJujperx/V32FYQSzYueikTpBOYiwGS5YT/BkhT0NWHg7bsT8gSSe8mPJavk
X6IJ9aanUB8oMQ3OF3FypqolkpEhcejWHFjf27yi2Y0VA6HSgAnD7NleNYmBBfQi8U4hDjGKJSnI
8P3H4p8JKhf4T35cht4tM4fqD1c7fx+NV9Q2f0dkhp5f0j5aDCdHL+WRS97SX/Yuwph8R6lnaxxJ
2fQWIeb4bbXY0SaBYsjIoMacRSJkW4MxcIBbYjl8oP8FCsZ5GQJbMF3nXbzAcj+xkDsqcTj1kOP8
+Ac9WyONBTzmRo0X/2rTxgUp4tKAFlZw309a9j30xnbelje4vQw83FQPLij4WEDxGvVKEyPDZm26
8mR84uP4pPHvf+JSZPAVcaHlo64QxB4TthyLmApEm3v4Sqgfg2WiSKy2YuP9D1rGtss62T1qAB+c
JatkJV5VlUyFaZW00JjGBKD2Mflk2ASC8B3bI+XN8RYVt4f3BHmQcX47kg4mv3XhlVbo8QWj9fTd
O05GTbyH6nBY/meU+ftqVVq3djnhQKVWowSFHc7lSaja0ONiPPmWI49h+2dTbw2xKT57onvlsF1b
o62eaCgg3C3zzYkTzKYOksoeWtaW7S9jjgbGxy3ppezgwtUsJF9FVhduHuMEFtuTpB/uIxktuMx3
zV5lC8QBFAae9GNj6ugbLJEPYlyz8yMz9usWcp1cucJkys6ixvWYDl5Yy4WILgZi/mY7Mex32Wyo
9BxdJggN224K8b5Z9wzcXBMntQuCN58sedWfRybOw1maXA8GHmNzP9R1og1U1Ro2ivXvSNfov5nm
WlHd3lqdTEeJ3X5lEahtbmteVOox6Nq0waCBOXLKs4Z8/qm3sdTRzxDWNBjPRuox/sE8VYCD9O8n
4v6egO0Nd2uWu9XiZmX0Pd6iRcgm34tqotIcICSpisnZDzYqYmZOY2Q7eYwEDpTsivEe5R0VZR5p
oJpfOo5kqQq76z049NqWgbOh6hH5XAiE/cFrAVPPXVfNQ4kZMsIHK6a45s2zjlpE3uN7sc22mbyl
5j1fRNT0m4LHLktK1kkG3jYq02C5rcP0SBndXywgPn8LgT5yuax5J69ar0ZwJVTIhdu7zzZNNZzR
0gipYraFJiCYE7qTIynE2XrqP55wrTlFItqEXuJhMehCjZyALQeQyZKIl3bvlxZVOrg9EU1qGwQ/
vm5/o2mVPQJrSgLJ4HooRX+aw6Besf/qQ27/Q52aU1qvLWpOnaM5lzpSUDDn4cat3swvFxIRfonA
QFyE3APykzftIxOFvQzHYjoLYJBkTFs8OaFQf7CIsZnNt//GIQTrGZYphRJKMB3imGt1L/5ScsAv
+QER6qewPRp2SWtdc8sv+58A+MATJqCUqBylXKiVyVIVKZLPPoUOYh068vQnDqZSXRdLvJfJphAh
nL/gR04fEJyYisRXRtfM6u4qoEi8JMqf40pu+7k29tYjqHhjMhh1qmszG6fwsSi6kwAXXB9hL3L2
LBxnsyNHrBoJRhnneRJKUlPGjZZBjwUDTIlwiCRiTTU5/PKDmTJNUpY6lkfAjDXeXoXRV7jcul/5
vDyj7g0eeEKcSqUakD3bnxrlfDezrHvzmJhfoVuJSPdOKIhcstLzFiQ0UxNb7kvPZesYzD/A/0s0
zbbdgCcK+TBHHPvBthd2QbGWRvag3/SAIk6Friip6R0iiBCbLbCRVLrrbZRTuLC6zZxnq8c/2E5J
bUr5upw1XLX8YaL25dnxMd5x3bnWgTvkmJifG+cLjbQkyxh4m7mY1SoUwfuhKzMUIv6ZUjrVhVjP
Kw0w1oeo5L55ihXahRzC+YWgXgC5SKJOM0DL/8YUBnwHr+SsrMomk7NH3gLyICdPqIXcVVo/0CA9
6Qs36TUsqrz6zbWJroYH7gg5sEGHyKiSgFspoc+Q9IV9I4tndMT1Rkru46ltIWMaPFaEy/TaqAo7
RNtF8tv4uijPUCPntVBwaRkZsuMJ5uQLSpCCEHDUcM2DPKORWeHRcg1F5McsC8aZ1vWZUrKK0K8m
oc0vR2A92rPVvcWuYoYhiB+1PSmidonqvae26SSyfZL2i6hKR/5GtruIcS+Xc3U2Br7mQHOHZJqN
sU9uW/0CXndzHhfmKQnOhtB31YIsfnSWsgsmYqN8uKL39dCnMy7FN8IakTh9MFr50NAFRtvUKgNh
c9Vk5K41sx64ttiHvG53OtAD+RKwqtYGda2o+ETBcjN3G8eMUmXv3lfBFXxVshGYy3aoT5gq9fF1
VtTFvQ1r7SFK6qFKAbNob0PR5Srd6PXe4M4sXm7+Uw5F9a/5PBH2DtSExW4fFey4tL+Gg1VthQvt
JJXT6Ie/fdaSVAgxAnaxldTImJbk6RzwucvWjeI9mi0D83vFfCKQDFxkvAGq9ddGm+tTkd2jSWir
zD/K00OYKpcrHpir0Y/vh7s+lmIjAzSKLoxOAIk8dn8cZAk5wnOYvf6ure5Ylxop9ry+7t8d9plF
BCGsGaHlDhwP1xDefMiIARlgb+6/XcrdRYgZ5FR16pE4H7/UbhOPOJXSIP/SG7xVgW/BPPb5zXae
24gOgZoRkXlAsbp5xmoNf4Rpr16jwaeI8zWvy86OfMaWKE/WHXGVMaP6D4KHZvZaMyRELTMRAXiu
U87cprUhwOWpCPtHsclFmdG6mxgYrh+yauNGdvHx2pJcJ7q2XRzBGVR1gP5GPHf7ZPffnSlK+EGP
eNZpDSXUODQpx7BmYyLPlVoGo3ISKVjFoZ1gPtucUTnKGDYAmiXkeg+ek2QKY++u1XOyOapqttLh
2+mvUK+FmU54r4YUuIjqVTjQyQSvpiMeRuiYIDGFuiZVsM2FatTsJYnVRenklsVpG/R+7WUNEbTN
i1UT8vKy5KdTAk/5sOx3xGsaBmAVDDAvawuu0bI35fkc2sKRoZd+2V9TEvfKHBDsP+rCizzMR70i
s9apfmvdApw+9M/E5CJiCuk0MeLkizqvlE5aWLZEwRFYHan13954VOfZG3Rly1Hd0qEC2RdkLCpy
rrLXRqMpTvFg9ulNgTn/91ShJ8jPR0hmFk8znmIpYto1wTyHaML/oVCPq31ZGdgS9ZxeCMGWZy7H
GTVLoVyVwafOThtIZfoEa7ScoDnQjQ6rusUIsaXkfeizcWV1SRK8CQnnLDa50JpdN+u9MYLVjsRX
BMg1fuUnXgZCgXXI2vubOnSKQ5Me18XCZaJIUcWOBnSc/aeqqdoGgRtt2/a02Cs2r0nt1ko9HFqV
n2c8hr//DSHr84JdeaPpGZK64O5961YczgBK6x3aQac+0JK+f/dm82QxU+QorFsrovBWPEvOwvFx
in48iM44ZizFknrpNvvO6PJp1iU2IUvKqd0gL/kxuo6EXdBIQ7Wld0qO0dKktYwZugsxtz5liWlj
76prdawffn4vTx2vKMsvcb/3IRYqkD/Isxp0/9Yg36tfzdxQ8urQCM/W12WXGqWHgZN/HQZSo9Jq
5QDkrIMNsUS8w/uu1jv2eUsxnqa2r2sDOuZ7+FO3XfjBUpfa58fst3qSRvEstLIXNzfldbqPALGj
QYOciDmvKBV5xtW5DAd4JLmaobe+6pzn96/yxzU/fTwzI5LGJ+FQ7QRxWQsOoMQvU9d2enLoqwsH
7c6xyHBsAtN3O98yJG9qF2kD0nyezSwvYJf5/3+JLVoONzAx/bIrfNpPldYmpE6yv0DMx8u8EGj6
brspJbBbeMyguaZeUsX2pTndzLCShhcBYEu7cCKsuyJSYX+QvFDDRpFLVCMdQsZe3wnLFCMRQ1w9
4vd78YKX/M2uoC1DKYAsFRmxfS36DdZfV0DRbzsltbwWRosyl3WyiufL26CpqTPeIPLv75rYhMXS
MEtnuwamHSeofvXgPOxZu0pwudyj9m1JGOa9GOr2c3g5Y39JsqNdQT1lGnDAucuS7qnlk7x2jSM9
N9aXSctElu0alOVXoXueTSSvm/I/LnwMoqEjvXUs7IXOW72K3n/zkV+RTCcdJfiKYU128IZMmC/m
P5ohPm5UreN0MflTqKTmABXx/TQSw4YiBiIBIx8ktLOytK1a7J+b9IDRnJEz+uynbgOa+/LvjoKg
L0x3Ex1KPawL0FpIs9MkeQVjLXCt1M1M08jHkDHEFaXl6+qSMXp/dRSd38DgytSiFscBDdHsQ0L/
nRzrgMWl5EiVVslomr4Uq3m5KJkKjkEFkrKDF37BiWGJz7Wgac/VIruM+ocV0RVBK42JN+ebKdpI
VARczz5rIfb9a6QfSbhTbBX2EQCNrUwX2bsBw8Yg01+WHNiOIMDGio1sX2yKmybvF7JCvu0vpye5
CdBFLLDj+ZszM/H/yf39l1UMUkAq2+1pwMRjiduFlHKi5bBnJeBla27TZTEija8bSuRO8cyXiSjP
I2sqkiTqe7Zz3VGAFvLq7J5voKAUcU/3Uz/PbqZ2N478Vz5IGDtTv5Flb7Irz6zE4m1hnR49568l
G3g3r1jLDsQwJ3eYJ7ug2Clk/5x4DuVD8Xd3B7AbWN/K7yqdx13ToSzk44qN+Vl2kWkMjbOBOveu
fzJNeb6ZyBKx142PYfrHliWNmAO+Ayq45G/hksvHeEXWzZAFjb+YjgX7QaskGFBGmmZ/Uw1uCysz
r0fRlz/6195lDxoxEMWnz98YVmSaoY6DOUB1wyzL7KaxIVMIsm8gGPy2NzAvbBT0Y40WWOOfHpsN
nPR589sVwvnYZtafagEoBOzeWcp0YnsExuR+S+QMJR724gboO+VvDyl+WwXwYi7PfAh6fyenP01d
sbNMpBS3OtHF9MU4WiBVyBb+b8pqNlp8utdQIGLxXuhU9Ko7r8iApUtTl9eTv1iAqG1LYjPaJyzl
P88kiRSvf3YS1CvUDZP8/YkWuh09dqPX/dEq6/2FISEIiGWPetdLzK1djRz+KA3D2wO73OmbC/Dy
LGa0ctHJ3+jeUT/CKX85b1PmrfqzWVwvGC2FExUT3FKy/79VPxYsUKBu7dJlyyxoHTPWp58SoHHM
L2dTRja6BOeM471mSDNlgl0XeUZrvFW5j9PeaHDyFfbEfkpqaBuqyrn6mgIimBCYaYQSw0A8HLNY
rgd21wHy2TmPq31Wip2vlRK2Abyuuueurj76olG4o701LrcnlPI2MJ23BAK+sRupAn7OB4bQeahD
vazrTanGVKHm3Z2yhiwYTPwDxat6d/E+JHj4H2Ov2/TTtnduUyXXc8ojyvPVrZsaQ6IWE46r60ps
YTKha5FxL59KsY8gEPzJOFJlO69IjRzfOEX6NwwyBdgPjcMT/UNN05Qp0bEqlRncG86r+xh568ZU
7ZxlnRXMSaN95U5Qw1kUkfO//drp/sZP5YMpXP+6fVcrl2+g/k4OMXbtgmM8UiFpRpfwa4uhnvHv
eqdGmdYnfeMyHiFl/VcbkIym/P9DkRLXT+Wf6PNzvtNd/OhOgK0/9wbnaeLh7BxpdIXUnJIT4vT/
fqQwd6yejbit3CBBQmJbSkI/QWy/GdPZhyyzjCCur42JkMuioCYnNjKdswlLRNItgURAjxcuGLpK
uCh29c4I1SWPvVz90/ti2pEQuskWjFG/KTQ5j0Rjeg4cCxtA52ffC4+FphAmqb34jaEfYxb3nf6S
L7UYHsLNWC+AihVuASpSUur3M/+jPioJRffZ4ZOR0lKkFEJXb9oVEs17Xx2yeLlvDzzVq12Sw+/1
aI1oDO/sUIZo4A3B1ddCwAjoQxrrKm3etJN3McGc+Y8wn5Z2B3rVDZ72FhDZLgF2SV5UBo0iWKdY
FOo1Q8gfpmZ/1fJpv7KFaaW81FKbQhhXBbIorl0H+wLKKvu7UrsLQohvDBtCv97xh7KmzU4kVHX4
fwkU4Yb8FyEV7s/8FVOp8c/oNMLXj6tmppoZSdnkx3Ec3pITRclpl5K9XKl3Idw/YUwVELMti3Y+
AUyD0OK8pCrij/5hYJG1+KrUjw9zJKbWt045VK+hjfx8mFFeqmfPh27MpZdx2eKTff0BClCHqYhW
7q64hfKYqqM9NYUcUJNqI8K5uH0+uZqmvWE2fJ+XtyjJ9HQEysrVw0qehdy4Bb34L8pQD9aVsX72
1Ei9yk/DdfjG6PXeeJ8SGZQFFq1JD5rWJUwm/E+T68bDMTxXmzAckD4yBP5rpfgrngAvTg9SonPB
7qFKb4J/YUiFEQ5U8taawUoiOqZ7Br1w6iiMGC1qebStURIH9j2ZNU5XzvIbmGkUExfNtluoOBIW
Qew/hHqTe7hBilOVTn4Vfo2GbKje4Hx2LfVmnYNIIsg2ymHIOOsk5jXXs6IfGrtNhaGB4hZ37jxj
E48u24rWP4l5zBLKa01dGcKVyzLLqQpvwGfESrEU/x4+R7i4sgfCQzQvAfITTYU9RR/UcJNyuV8O
JHYFAvdfV9Jtd7SFbMt8aDObknvreUd/jGanqeXtvlJ8snbHjij/vynQLnLhpO1xWDiYA0lHzXhp
8QXO9xgFkJRDY67mtTsGaMyOP9bV7VulEIsSOhKssadDIUFcmadEKwT/i3kI7NJa7RCDrd49/hWn
ziCNo//nCh/FMWx0JURb2FYjK2hy211anoSeZ7ZdRDksNjw5aM6vDW+WLIJwVTNCgWlL/PTOgnbl
jMqElDBFsGd4FSLI/2/wFuEkz368yzxkTWNRo1pTzt3tO+JOQX67aXVYk7OtwrlKffV8fN85KtSt
gSmN5B+HqU5t8n05O5wp5382iWN31dhm9052bgQtzALiZmA7HxFBMzVhA5fRG/1GbdoSXkXTrB/C
/QcfQuhy8og0Hp9qvjE4Xm8E/It8sGT7VZuVdXbPetoQMf8y3IgZhIaEKPpEMLbGMUn72C14YKtm
p+oesApnlnVw61Wo2nIIKShcLlc3eF9R/C9mqzb6VkTBTMuBhd/Lx7zVAiXMxKc4MktpnJaey2Cr
T0g1pJ4YaIS6+bLzRy/aFGrqOKR3bpF975WFDuEF09f/nrbiJAXcUy5W3qtTDhvuyE3ITkJq6AJY
QukuyR2GkxV6wTzxEdYeWj2RTxJm6D0whMHBzAS7QSdak24NyeLi82M96nQROZJCCt/qGqr1gTnX
nIHCGbkrhm+8oUGLPTTC2LoL3oDxbKG6p23K3dqeXOONVhCt/FT9CcV6X7AQ6sSZnQp6DdEeyA/g
qmSJ7elcbOrftuHLMNRVIFc/V7r87c4FQNC9cFI9KM456dZnV1z3IazpbslrV4MmOrseg30v8+Yg
+z3C00cVPd/i0LeGyiEefePPx4XTKmpE/7E54zlZsj8VQjZlb/S58+ZM3gpUg8Y1+tVKREMPH10+
xzJC0IUaY+UmmeU/8eQt7056zbCEttcvyh3VmG2r7rOesGbsatxK0yEA+Fpcq3OPBObInRNU8WRF
owaK8dNSqYHM4AjUK0bMXNyLvqpxqk0ehNAMUKKhmTDlNKHMs7w2H619u5oaKrUQEp5yfvvJ2b2M
7tlpfb2AFVOpSX9HlUcHaW2E0x1q509wBzRoRlnus9oWNiT07me97hcSxjpB2MQJygqNHpbJ8Sxu
0jaqGhsLyik+2rHVUxQo6ntJlgm4XO5B0sTFVV0SMnT2uxg91k2Xvi5yA31ZMMARhfZ6f/aa9b+Q
P/eBfdzSK3tQypj79C9npPpoaVypgNATjl+ROBEXPOvZ4ankqF0VVReJPMK7cuXp+x36mbTjSdHs
eh831XEfvDhnHGGXmazYXIn1J+k569HunAVroQQBAcWEgLyhoRgKSr/ErOqtHDlbU/ZnRZ1svf73
Kg1uqxwNODkYrlEXdI2OvhLCQDpyJYIg8ok2/EUAKpPKQmV02bOVpMTL2dq+ESRVXuzKvREBvfZm
VWCFOd/6tX82UGus0ZSzxUw8koQBUWJZvddcqQRwZ13Dc/Eorrab8JXa/gsWng4ocdpwUBJOq3HF
/3RwZ9Gv35+PQSW3FHkLx0BP5xrfZe9KKLsEk+LlHQJXYSj1s/uQd5ieA3QfxL5j7ljrepU6brVY
FKDN7QyHEx2SQW8cOxACADQ3E95KzCYEWm6Pe4EqhFm2vO689nzUaFQ+RbDi9idz8cE1w0uR1bG3
mCNmVirK1HnEubIL57AwsZrk+oMOiHs7ebE7FUozNsxef0iP/TYI3EYrebHnJIDZGNeQ/ICJGNnY
X1JNbDA2NhhJmkH00sQ2soffA64mJBKGByS33gQQ8kd5sjD1MkXaSK85aXSRsMeUd66W3OLRZnCu
jS6h4fqYyC8f24anutbSkJK69bN1xz0p2c2CeQ1e2JNpqy+GynLSWnNWajchEp9jrKTAjGljjOIJ
WMheeRpWXVAV3sC96K5juvsZAhMR1eYoUAMSfjesEt24JTyzkkA4TT0g9rUh3M3d3v/KSWObJ1wo
JRIKReGqJxErBgiL8HtILyXWoX449RM6PI29Kt5QbR1kHoROrF4qtREkFvZ9Wrux8dFL0XmkaZkP
ZYyYFee2SuqPoExNL6u6K2eMPUHXR4n7uYB9wV+d/iMGLRt7+W8cBj2ZPNhTRL/At/qcEnc5H7oN
01mxv7y7nEKyKi5ewdkx/d3g7T2EZjB6HNEeAfZZBD7r0HJ3ifp2/9FMEOYM0Yg+Z0mMgtfoKdo8
9Qz2WHE7irTUm1wBtPPYbQ9KD2J1zqbjR7z32Kk5W42xS3ukODWu7m42aiLVTNe7A4pLXOKXVKIn
4VkPym6xlEna2Kh4fk5SRugxscxN/l11XDu/zVT2hN62pI9kQ8+mLxkPwBSwOvk0YRK9pLdCAbU2
AwlevapeuZm3QyCcZC6shbCe7G9QE+vAbJoTtyMJWKza3E6u6ToZUjwE2E0Le6b3lNKnfjqAfM9d
MpR9o0WIBx/PhsUygJf+aKQXQcXe2x/uZBr+LNrxfdta930UBMTIIDHbGHOX7qSCvyjtmGpUffAc
jmw5AS+rSXMEgv6SBQXA4ho0KuAKlU6lB3atRo3oHreWSKBbaS2bp+vcPoe10yW06jfA7jHTecxC
C13BPyJagAwvh/g8J+4C05nD28CqJv/szL6is5HFcYLlN8wJop++6FCBe198y7bRGs8W2vEVdeQu
njf0falNfJkprJNv8fyj6fzVD0gVSpnDcsEoPad0LUWVkrw2lY8fbGikojYg93kgw4lr6eGwAJma
Qomd5y/Nq2ZJUTq8MUrDU4CoHW56MHyBfmcjRsi/61so6+vQvOK0v31Jv5aVAZAQVb7vMF1jXaik
UpI5PCKjWpLLnAJsTFmn+OZCI4R2Rtr0fuaonz/VCXXaAQyJ62Q9bl0qC6+H5IKeRPmcBBcwkFr8
DF1a0qyzWYvzDzhlFRFcbVohihjjJ8wj1RAbvE96Wz3nBYScGW+cKSTE1fLrT6Ho0r0g9SdAhaoy
ROMC4hxKR6j4OFZ1+UCUtR9P4mm2DzyUBpI2G8RK39kxh/XMRFWPyL/T0VgKSWV14N8KNU3pyYtW
stXv5vQy7aNG9U67rXqLyEdsFp8l9FN5TBxuTLg/iFSek9xuHD/R0nx6fKt2eFMDy1KN4wYlC+wL
hTLSmII0Umubtp5aylg2EmgElwW36JWrb/cwaLAjNHg/zU6XY6Ujg5N3e8gi6gUO8cSh8bW62DEJ
pKlO4Mq1Cxd89s+aqVTYhS7sg1pmuchdzAcrpbi7CIVr/7luZAf/Xkh9IGgbv+axbRq0I3ecG9pB
brsPHOj0ZB+FIxsohH6fuYFm41J44qIRFnHZWrYCwZUSWGRQsarZyr0msMnoMnxWnAD6C476k+nY
Onc8rFEbpLP9iXpNeS+MtyJtTeup5F85SqiSnqCHE+Jboq0jFNtGsVepB7BtkcxS+vMqQxA5Vr3N
vKdqn4fEUVmCJszPrRAmqrYTbZKkQGZZqu+Uw0sQDDXVoDRt5NxAUDVm/RuHn+Jqx3WrME/zfp4d
a96tudBWx9F24yOuY42KUwC3XSekEehdi4jfxtqTVqah/NEQkvXBKqxQf2CI97s0efNTPj8AYa1/
ioTMFtfGw6o+WyLEg+4SO8INQMieIkwyYflg1UOyP0olGMlP+R7N+vZ6KLGTNYejkw9L0oNJ4S52
u7rEijNg4vusRhjJLkNAXsQj5Y0D3ErUh4b6w7Q8xkKP/iiDpr3eNOxfWE5L+XUduSBAUrDo5LTM
e2rw0/IHM491Nwm0Ghdbi9FG5e0VeWXUhmvTOubmoRufmY3ky5kfUKVisPfPyMgNe4EIMMekev8V
gNwcZpQAjFPsHObUW4t4Wdv/oZFPDOlKOxeNLVnHKoV3VcHEwImkIP+AYsb8XebVV2GFBEWEA3iC
teFSXmxf7vL73dd+PBGJW72sX+5cjTJOkCBWXIEzzqmmSgQ/OyVK02hPxkGK9pgXE4NaZ7ibapqi
xCdUy6TJDyOOwXk6mkuwuQNpWdmYHLCc4eHFtjD++fuCIzYGi89x4BA4Cmw+VKLnJr5kOlyzus6H
yR8lr2uj/nuXIWwDsC3m9+sIVzNAKPGZgG47wGbIuj27pQIpUdnQCDdaYuWzLerQnEAHvTkWfnRF
imf43Lqp/7I0gWIkJ7wOpzyW9H6HEPVpi38UQVpXsnk/6JU3uBhUsoUmLR1wAOhb9lvSeYm/EQyW
ranNt44nOtxUDi4wZG9k86kAU4j6Rc+ujXMZmOyKPmzIbmuD3O7wVXmOYJyRW8XMoFOzoxY0g3wo
CNnM98cJYteF+s29h8ANeOZyq9AQm05N4FlHyCGcKNX/GUy+++QU4AgE+b7mDYOq0xRLiCug2V+O
tkZB0GabK4NkpchcEBZ5HRxjVCidseoqvSPqfCBIuGmeUsnPe/I/Bkibdmhp/TehkHhHyXYpEebU
jqKMev8PDlYMCiJwd9T8gX8N3mbBUklyCUKq/zMh+tpOkjKixTsoguIyfm7UEVikiF/H68VHNy4q
a/KaF54QgzzrxA3qj6DX3FTaPAN8hh4Yn7CTiNAv9t9V8jw424XnLHw7KAEvOy7TkcQuSuNFBy8Y
bQ59S1UNOnJz/TUN/4TVM4YLT8ohWjIKFO4Mp1iTJQVHP3VsJQMuq+hOCPc+X2d7KkszfUkjxOye
x808CWgh5tdn3xHU8BURdyYk8wO+JmjOH6TBuCDicrrfcaWN2XKR5RPqpQ1+5QjO47+4KdkUOdTu
VDW3IPZ6MGw55jZfYXb64NcSFvBhhHzv2p1+zKnDRvxIZHjwEmDtMHqOHjzDqM4uve1h3y0NixDC
Ze9y03rmVwBq30A/8qdmSSSSQd//2uuTaQ4twxg1rqPXZF+8b3m+jfv+008yAbhNg9+JoVLhwwy+
BDxSfutUxEpgwuERO0micrbz0+1/UKmwVDQopoOgLaguRqpq7cTj+YKI2mQYBDT3kQYL+OpJV7yd
UnkEUBAgQjOJjY4ekBbgYub5uHhWkBGtP739v2mEcmCR2yuAWI9d7T+XwnfIJBUVK5nWva0k+xC6
8NgfNN2rbK03zxXd/UU7u4XwMGrCZ/7KNOdnKvH3Co9NE9AKFwqL+qdgQQxUfy4GNljDC6IZOn2B
1oCnq16RN3++ZukzRE0mIJeFuYFkx3tYwr5trXLS6NefNC5lQ57OvIaGb2U1d8xUXFVb2xDQHngL
w3GdrIqHnfMUDG0uaMSr1KrkbpV+zKBt+0CkEwXYzQHlC86DuWYsjOgiBzJOVFtZmEmNTqHgPHur
bYJEB7tumPDuvjhcyupDBDGb5Y79Dis74lGC2mYo7iiYKn1Bv/0rxIAgLuQ3F7KmorhmuXMcRDh+
H2SBNd7duH1bZlZgvLxGganBUdfGJg6i3ZpSL4MWUvcN/2ROgQ5tG2DCMUIQqfi8TnN13YgYv5pl
HBuOrhCC1xke+mYpjFLA8PreFg0U0h8JUbYcAHvccDHjMpc6+FapudzzG3wSJVSeR2suuK4Cw7DD
WTeS1LHEKxcLgfXczlIhuGGM8VVmddAZCgRxi1pSzIww920Mrdcr+vpsL+kZGY0YeisXFTYZcEPs
EtgqzIUKLqi2mVKHFDHNGFk2aZXA5uXX4et/YdXAOLJr0TuwA5bIyrjHg3Zp5qI+7p5luQLOFPxU
Hjk0NpkJ4icWMoOk491L7QBJCFKSPVF2Z4K19jMa3YSjY20kDS/jL+vVZqqRPacmvgCWrv8bquBM
ruAsl7JhsPOuSDECxschztSQXTxti6mdED3aDEJtsQqFDAxz/Ue53UCoDKo6ymZfzX7wrcOWqiPY
usOebppxaSWYU53P6VXO3hq1CsAUPfX+05kcrzLBxuyCkRWa8tguqsZ4SMOjK9Bv3hzoOJdafWor
EoIVBmFvOlvmVJqNRzwwMIrPT+Ac11wYJ0048IKD+ggNwl+s9rq1OUhp0TlkRggLqtpDvWjrvSUk
XLrPhaZITKzqAlkBUI8p5XjjFny9DNkzxRaKs3z6G25qDcoyn+n26zhOVDVLWj4hrDeNjIyR/+Zn
5Bl0N7Kd0qw2JmsE1xs6Rn87NKQg0BWIPoI424IhO2/pPsSBtZeZvhkTHG1Gm8UGlP2bn9FggYpe
TjdK3ZVuiNNIfblgSrRcqKliX7lY7QjDCXudhyoiqfUSyMwX9VweUMmDC7mKkyr+w3Xl83y+pF3E
+Cie8p3OJsVLVEzTy5iZ4EfPE4zArDVio+qiTWwTuoei5I2Rvl1YHhuiymfiuNAkYgeXhzgioz5m
nSHbX2Ls/9uIM/sX15Au+H19rv3BpFo/t4nJybGDPXb5jxUsw8nfzcjPqGMPkKE3eZYz6fOxlILX
+FDw5YJwahDtgcjJ7aLjsilff0z3WcXx+vY68Z76b9Py+NUrdno5y0HbLP8SYfMfzC2yhqJhmqfD
CPAmlXC3DRac0QLsq+kbOTRCN4qJultJ5T+rYNyp1Vo3u85o34azlFZlH5JnUdplBA10zd2veC0r
2jmXVfTpjldT5r9yCPcQ3nGl21gQlkYGyxDn5FnSilVtuHaIrUte6P5UpSCL1RT0zL2U6+EuBNKE
rFeGWKuZbyACd49UMMcQaQWDrvk3csUqha2b4ec4tKjuJksBdq7nBJv3UGBCdsbpP0Eh8icwzUq+
7irxoWxM/1aDB9Suh7xZfRcmWAPuuINAanqSQ4mQSZ/rlX3EyKx8GWNLzQqsySVGQpUao6KVhYBK
AXOu6x3kMGrrJqtuH+rhDLwlvsuGB4m/oXzrGK741cK0wliGtxxchrSEgkGxccU9o5oarSUZnJ9R
qUl6aneeSnlxZv5GQH6/A3nIBNvqs6RvWHyaTqTaePaide28KdMFbFN4TFLk+MdkpHt6HukALJlW
twzwRAoInm0S2ero+Y7mAKtgjTMO3+01rPZoRp6oY+cw2cR7C4UaI2NGqqsG6V4tYoi21O+i5TZd
87lWucbz8DFzO46ONmBb0Gdcww1uxau+alhT/rxbNTqlRjaB4iqUwVmOR/tDxGJU1YsW8faU4vKY
azQRJqCGQ10xBW67heFR1rHx4tewvKAD2Hv8MIZSYIZLwiiruV6E8qcxSTkcnxeK+XqSxX5TOJCG
+Gpl28zTbINORakRG5J/kzEFD7Hztw2Hm12el43VbF44Ce9EYtx/yKQjh6qNJ5q65tvum9bi/zow
Vf9YvsG20h+tLCfu3Dva7AbNuP0JRXn088dybQixsFp6H19GM6jANG9f/2qqH35GrLLfK8sF55AR
JObIwrrozibgSiHpLkCX7O0l8R7mbXhAhkBakzdUSrnAjJYFG0tVRxfrJBBu51qAk0n33cdlKxbd
bsR3s+1sTcDD8DuP6PxGVo+XeEYzBHmN9zXwY1gsdfcKiBW+9albKuHuocTx+iXFtSK1IPFdrXbw
WVmApX/KhR4LkaYiRYRSUE9I44TL4zD6r4f/vhGPhJmxo4ysiSM+wvpm69HVSmfNXBPT1O6RvNqv
7WlYKyWpg7wvRq6b8kBcRF2QR6F3XpLgRsc85amsjMQnZ24/uxRPaS0rhkQzCmwu/qkiyqx+nTZ4
zQNzTUwjlVgbQJB4i2NTxDa4ehmvyGh66O2MlG1NVTvkIz1puHh3XHvcqcISzPesHu0JYwi8lhie
pFaCSnKagJ0TEHgqgTKY6OAm7uVNGVhMZnyIs/rpR8sjwLkd5TU6Me5ApAMUbi3Ezjc2m54hEMlb
3qGdvWM2YcrMqgBItjx/9XcKef68yZyOl+liZS0in33MYMklqe/xHtyi+6oQ/5YCoyJkNyPf/jqf
2lZ0Dg1quWOiro2VcSQKuO1Hjxe0qCI6cLRe/x065JSXrUDqxkN9AcCEol6zPSazKTikusjbSqqb
25nN5TVXE1k2gTrg4Nq5NpUdHL1qFRxPZskWVkxN37CkWf2R2bhXQmZaPoUW3Mm5AJA8rej22fXQ
nwc7r3wEYY1o4KKmaFixLDQX4bxKEUkssWRIiM+llOHbRZMpXHQdt5xVeEwmSySNZdc5XOwOHivQ
fJ36Y2q5hgdSstaaPtAqvvj3jq3B+ma6vo9m2TGNpBC8bGA973IEhkAVqKCssVy+N0jXKdjnfwEF
8dXTZFt3ad03qWkIU4585k3CWiVE76km5/rso8E8OWYx9/vglj5t6QdDgG8JgIsyPmWRDTphgEVi
P0r+ZC5KavJ7bzf9rAiXvdllm0SeU7Ni5A9qVX8rvVgbMcYCSZiTiRGdhQBWcoSmkonQMPeVH0VW
UTvPxUPbE206gHj+tMT5f+fSVWdoExxDF8hmS0CE3fZPMmGXYifGjh6NNfhFsnMB4jlytdA404A3
KZZG9tsExoRXPxfoAdioaUzm5pnFWe3iZRPc3Z6UNO8GMF0pJXH6D2J3PSnaDzAu6ko2GGSz5OJV
/hbKNw4IfbcR05QrHkrF3M7cp+HBX7DBaNWeixTXYGd+FpP1SdU8W+kE7IlX+OBCe0VzOmKtTbo6
bDNLb5pV4oi1bCf7oF6QLtCkNYYhWYhElax6C/2qiaM34tQcCoUS7fq3uoULXpVLF63Nl/0jDA7u
tiOedc5aqEluHepgefTL1+oNiY8yq5kpYSBUVM++/inlBqGZuvfbCdfU1Hvz6h2FCU4E5/tMcdW7
/nW2/fOpJlZ4P7E6Woi8bEm11OzkXgvua5Rcff5OK1U5R6+Tpha6qUQYaKTBqCeRtM64S0vFGeud
eivpsq5+xucXO4Ppp9dD/MiciG0dKGgmizzFI7cULo2tg5ZOkNH9tzHJz0N6q/RwyWzmfzAVnwzM
g2ad7DuDnoCx+ikxbk625JuzZZ2Ptc683iZzLpPc0ROUI0PuHh8tpUYvheE36sQ5j5FPZ2R2bcjo
mDQyiMX5NSbNCgSRacLaoqta6/gJWhiUC21XGUH4RUrO5VzDYC7XTwBE8WARxuZSB4hSEA+/DQDl
pGZXbUSOOKZ2BXYcsOnEG+ua0OM9MTfxiSRMbaS1rXjgGUplWZsspMwtLAC6/2LHfU/Av0KYuAKl
Az/mnPSy0rV3q6FIHQXqBWk1SNDKDw8F+adeFYO/V2cHFOlH2j5sjTRMfp425Jg5faa6qxXQtXhv
O33hPMcjX6Ihsit/nmD5Q3GjKDjGIE4L4JEmFf4C2MX4ZQk6ELLkMN1aWNYVoO1AQlUPcXAqqu3d
Pcud0zgAoMhmo4tAmbqVnNGK6fxX9DF3eGuNXVOL+vStpfsgbWkIBKUr/zZUzVQsT76Nl11BAQpR
aSkFF6U0iH/weYiWZF4MENsqRZq5jnJIvfSYd89MyywfabMyHM8hBzkOkqMSp9XQjeP4DT0SOgyL
eFuVati+BqEqwOPAjbe0YSKWSeY2lgrm/ZoQzlJfjt1nUnORF865wGVBdO12maWWRpzGtmLwXm9w
I7hie8rn1EBie2d8lYOdEDGfxwTrz8pmQAl6ckuLDFW1ERKfqEuE3ApABZDsMJbSzvbxkpDC/M2X
nxI3yG0sH+i/hu1XhUwCXDXkozINKN2V4nU43L0vz2uaI6MeJQZQsEU1FzG3emH3HSgaRmC6C8kI
KjpWeuNgVa0o2FXQr4qpmHUmfSvkoTfegBJ3oKkRj4oQgqbLFPLzZgidSCzgJkgwBZaVN34+yBmW
rTikuySbOWYuK59DiNCCIKnrif6Veh1iPpFOtYEh5HEEhP4bvvCY/CaHxSw8qVnTihc0cwEhY/Fd
zQkVrDu2IIjTNIEKPuHQURiqZsE1qH/VCa4D0wQWu+ehuh45+kKCiPSeMxgGK0JeVCuBgVTYiao+
TtOQXtN7H0NaB+nA4D2wKdaPHYuV5DEE4FmRXdP23nGXO/dS+ad21Y1chHUnsH3HT5omZA/8I1Ba
jPQsTn6KZe3SM7IqTiHfb50xDhFzXD7wKxMgy5rUw0FPdnfalN+Ghai+kEqSJdJa7biys9ss26bR
2I8r6Sj5RPup8MkaLay5xU5aZWYm7ttcioVcY2E7x+sLZu4CHwU6cCfUbczF6jmoJSkB3680YXIR
8J7qOmfLA3aX/o/nJZwdMlGaC57/tojjEkzQB4g+w+WhkGiwjLYCrPq/1fmLAVWS8Pf6I+dCBvOl
zH1qhDG8OrHKjXzUvjl4z78iJmOLjREM9tZ8r8aksaHW/8xlDDbrRTI8H+0w+d+aretNMib2pxPT
r8k22a543YK+IUxZxL7gUAUAYsiR9r+PLK+qoTwLQzZD+4jOvST418JKeEyI3FCjmGvbVFBE2waN
eug0vzpae49OFiCSubNLtwW579i1BvmzJUGliv3/ZEuLBmT9CEhURZ3Yxxex0EGB/dxjTll0O61D
+4FwGFF3Ea6eX5gwXprm/2PvkAYcxh401mWPHrQJmiWScZjwMX9o9tAO1meRTwow70CObqwY4Qsn
kifzQJSgxmNoIi/w7sxQyfvZ8vuurLdJbeZScCSX6Lg0Ea/cWRZtYzhBa5PCFKrlayejrXNrZECs
lL2WlYhc2If8D1NZn0mlLiTsfGXvv7Tk2TT8poIbZyTYt+zEOBI7uCPRJugTeiwubTIlIYqDVClj
wp3i6kBUTGBkEHj1wW6DNL1+SJD68nkRtvAOUnTt+XJBI9g8XdthkneOble93h+x3lHz5poj9GBZ
wbmVkHZl4PwjWXiBZIhQ8MOdQ4/FwqypERnzb1f9xI39Wj+L/0u7EsAzK2XoEIfFKJATCFv4folK
xqiukLMjJmZV2TvDXPGteID4etMxxF3F2lZX2gt1puOzSuF1b/UcLFrgS4kCYbpEMaH0gdWvGqSi
SQpWOPxclxtkPaF6JJFGkQtB/WMQ8pmtRMzzO/0WK1PIXlUvt+5vda1pNp3zgLQuGZgS+CGfVs0X
t2/g9wMkj6VvUDX1q8TLQGwmusBYxqvF9wWg/z5/DwYsrn31lAaWNxKcqE3zsqFp8ID3lD2sL+Sy
65XET54ZDXy43U43SWR2JfMrCOB5X22QQryW6XTwEonlzUgHgJfZkHF5AGLz1vPVrhnXssZSL+IX
HH2pLJUNaijaNFxmldslWcLKGGxKGpoGIkqrLo4Vw+vZFy3SbiNMaVSL+SCWjSicoPYAZhR/cOdk
KDXTMGTKvYeMaHf9gMORCAq+1/+BOiQCmCwboGo0rnBt+43CCx09mQLa4kcc+3l27dx+ZdsuA62F
yTzZL/+1PRIcdkE9K9/2BbGH29/hqqIryEXZbOyIuA4BlT2xh+RPcYhX6YJ4bEz5eMKUcwS/OKnE
4VvW53YLEjYyVT+1nbVaH4zaVg63nWX/J6YmASB6cDRZaVBQh/MqlGdvLUhHlD+/nHW+bXYvR05R
UpN/ObU+hbuS02xJOYVDZZbugo73LYd9vRnLF+qAAOsF84ugJa1HFztAx//KA5zH0V7dDl1MMQz+
bQ4opnMEQpPXMVlQdN3hcsCKLnbDtkcYB4tldrCryNgPezRV7u/xrp/oG92pmHFwX9eOC3N7A/Zd
YuRKZ2sJ7zWXgWaHQqE9gr9t0ImQDCsXDJZzjLR95MMi/Dwry88lvp8gRW6DH1S98ATszHIitGjf
EjkFI9wILD9CXnh2aWiVvr7shCDx1dMeeDZEHTL9CuLxAnmHjayjWLbvxPKMpviAOocLGp0EfzsL
eVyVV3mC2LBz59pyU/46y4qeTmCSWcrmPTZ/HWNdISibW2EI2gZ7w2cXRaAu8JcgQbn0c9mwDhQK
UF/zF/mhlmwIKifaidFJ2BjirwFKy6XVqIKyIaugmDBzTKCavBh4XVvwsvLoRIkdEnwNzOH/X7KK
qltLXE8Mk3Y/ukEMAmyMv76M4M4GTRNeCkTR1ahJVcNC1Fq5VfKhpOgSUrkVUKvVA/2Q8KNHiR4N
vwnomKzTRTj3dYxz58DHRGXXQ6HTPzBo4KrmTlo4NU/vkl9yEO9NeuopJ0Iii2rBZtJQ1x0WiTFi
sNvxjUVHi6HRBv80QYLad6jkb3zcAr+9dRRUVwtlNCWTF7I5TLxTUmfayJQM5usX2McgfPObWkF7
I6qw3Ngt+IHb6K/5peTH8QiBP76KpAZW2lW2GvslE1m0Az0G3kEys9DULn3cy1vwDi1S2BHZEZUA
5/+au3N1rvhW7fiWgwz404AFCp82C2kA56KGusj7a2cSsOirhHiNYL+U/UhbZ8srwMOOMqc3IoFU
3G6oHjtVcv2VmmJ6n6oQUMokVtRBb8Tw/RTrbJFM6hqTzrkHKHahFchRX7Pk7niZQumZZtkGQCNb
4JLsqh6pNMHkc2HsOd6N7yEPq7yHPpgEyS2o9H3o1oqMgT68Ao5I+DujfKDAndgjPTLXS7tnH7kf
6W14EfR3c9tPHJYktWbZziSNcMfy1d0LLEYe6YjPsTFlFPEeP6S/72BQ3vUwAylEjtlAky2lygrD
/bp6GzHZdjcRGkGBuje4uqwzRWgusNL7WIsT1jONukx7I8LjDf7om2RCI1OqoF3Jnd3L8cg69uNB
Im5/fXqNwBu3Q8loRKfD3bqEtYYURfHBXF6QThpxg02DUSJAPIy4I3M5wmLGazZ/2kXRyFkT/dLY
sM+wSjLCzt0LpU3sFY/VuoggQ7NuM5anyyav0UCuzjo7iZp3q/RQs4SQQ9gCt4xubhhFhqvWBu9F
msaSLRZhk7p7/ys8aVa3p6h5RDUGLIZ1JfXaaXtDoh0ZqBqrfpvwNNccqG1msucyOKYpzdxmOVAL
shkxYex7gOUyKpClvtEvxLwI6kfZUknJN3qlBDj/pl1PTXwfJRQBJmTE82F+fK/we7MypwyuK+wk
ys2UiszlN+tAPFpzw+cXI5SoLeEyCt4Vr9OhAd+uPNI79F5NQcXj7xRZ841eWsO5OEqQ0fvqN7+P
xr1/jkmpcnKGBIAKy1nH/OwehHZctshAOZgAzBId76pZUhBGtlbUzqqLHsRfTS+60Wh3sWecGnzl
9K0I/Oh3KufWA3a0UDDfnbxf4gzgJ55wYJOYPGJh4pfqGinxNegreFvPbNO69Vbj6wJkxVibOp+2
Kp/JCMc7+IE2GbxdEEIKImDMEQ8dxoYf6dyPzI+bb0qQ1pttgCTyHYG+fvt4dL0ylAMlSwdIz+af
wLKdetYFCt6bZmlV83UWTQG4WmllYY+OjJdItyPRDmSxte/VICrS1d0rsUDFUspI7mQibJiwtLAV
P+2lYqu04s33Q+ee/bT2NrpyTOvHXj1a5P5Kd1/VDdf3++auJWVGZM+o+GKp7MyegLL1Mb4UhaFR
K6V+062s2Kn4U9lU4jouawduw29JTs0hVpgogf53rLpABXYqiYbcA01mh/RExB9IWgzT8dx58LqP
rO5iY4XnIT3JppTxKldiKATlS8ec/0eya0o01SuubiRuYVB0ZkifDwYDi3OQcB1SbU1HzcbZ+lCQ
FoSaaM4LbIosvzgIuoc9AT22YzIltzahxRJG7Twr5opLhFqQJLtI/sCEAfoBvUUCdRx0/XHlRL/W
1U8RORLAbcx/m2NOJ+DNUbhAvVgZNhbikxwGg/fLpemknU5cG9++FtgTEaqxS6TL9EQzHdx4tUVE
lGaBCsOhWbryeUCLIa/BUwql1pnO+JSo3ydPwc53a/iYe5E/EN+3UKtuf03nZpk/lnKBiz1iVb71
u2OKPyQ+0R1IDdtNSlH6c8b+9c+xRFaEkLeX67OcgZyER+MUCPjgeh/36OP9JLusrTQB/gsB/MCD
jw/NKplJo8JzK5cpl2cUB/7pNIVjiYOoVY9uk1WVdpmuKyiJsKNJC6h+gMOhmyFaqMCp/Vz1ccak
y+1HaAsiYOp8TsNBBBHAkQeh4kuWga42+lbnEBoS5bnlAgfmEALsfAlhJpWdPJalrt9fYyDOijWY
RwrqZdOywTKewjAVNL8Cq7XgLvJ9hLdt4b1bxEVyupw43grb2nkfAr++Qg0aKwLHF+1XcOpFZTmR
09FeLReVvi2QA/b+/pPKDXiiKwLYn/67U7WsJ25gAiqAkJLqnko6eORAMGhvnN3nlOF9is26SBCj
49TIz9VmRSW3JThRXIp2v6jV7T+OPWsdZm4HdWWAgLK3EzcXAIIPLvQ0nF9DmQ7cjptk4HdiDooT
8bV+JIOMdvW6PZxJCUUtMi4GfkHg0DaF+x3OLyV+fIqfVmt3+po2e1cPf0r5fQewzlKzk818G6JQ
CVOfm7md1zaB73+VhdSIdD935sigSd2m75eDVIuIs5ThmRpIHbLi/3SV4BXlY3texjTuHs6yWriX
RLHZHXKCRdoniXTRRjh47CRAwNCjLVJK+6qfllYryTGgBHFaTRIuMP25L1Njw+F1/45eWT4V7Oyi
/I4jh5+6E9QoE7FhtLtJJbJnKZIuuNPyWEUkGOid1bA/P3/2G3QhXBDhAIbASjINC8kBlNfzawWR
/oyL6SCeCaI6t2OssIiCXnvoDycax1eRutTOcPbF+4yOn59umcyLwHqonaANAKbSv7YF0qYQnH57
1yN04RRjR5N5HnWmKG4uKICoPGStGvXu4t+SIclhrReksw2vu6KlMRnQkMR3DWCSyTaCALvSGv0p
JFUYvvRlkLa5hzxSENx77OJWmtCr1X9D7Qhhkk2Q/4eoQb49PRCEAWxRPdDIkcM+8ZUjP37xoXrB
h78F7eqdVnxbQp2/w5kk3IV40ATTjkT1c9lTmwdQnzi5BKz6xar7sEsWyOo8TCMwS67QPEonowSL
/SU3fYIl7ijHVVcLDmZEA7PfiuYftHKLa00ZiNxUOASJU4y98w0ftmnSWoiQKeoOrmN41ySUTW6u
7SOKxhyyH/n+sAnWkmuCcPJyKAGvP+u2SHlR/TAZJy4/y29Aa73xrsaStEiTcUERvgWV6Q9gJDQc
4Aiq2VxpqVcHf/n/Q/cJLe/1CwylBoHwxiUZdfYSjDew22gNJMurTP0vtpC7eotlzYUMc6nMCPeE
XHPEBZflA6ZQaPBndmZN/nY/RdCHf6cVFPPpLrapYX0nEZPRIRwK7WYXR+15E9CySlMu7xn8LXky
HnqvjJrsl9arPQYXijIhHQG6kr32vJNq/LIpwHxwpZseHtC0/dXOCNevVm2CCmbqzRG1WWiFUap+
b+ncVrag2KBjt+wJyXfar7duaYYydADC6OasSUEw0F7YJGUxHBpOOU92HQhIkfsTQIKMjGgXgehK
JIiu9Uh8RdNOb0UVQNO/uD+5+zKXcmAfg7bgv3lHgo5HeZ/pzhNR21Vbaupgcocb+B5OoVAaCSld
OJ5Vh52XvGqpIWWlrX8heUgERxm4Dkl8UJKdAQtWBbeBjDGMvui1rBKFqBLlPUgXv85oUW6beUnE
MfFeJl4ZBppJL4iE7Z+ysXnrTUBY40FHJNJE3qdU0SChYWJ+oZ1JQy1mGdPMeNq+0u9fSVW4rsfC
ZAoSnAKNITIrWzneMGVF0dnJW+S7pnTXQnNoZtilJemh66Zq0xK4zy0vKVYwyj/jGiHnHLx+XkLt
5bsMPK5Z2+rOXKzEesK4puDGUZzvXUtHQW5fu4Cu/T/jmuEEStqOeRqsxeF7DC7p/eBLNB5QiXHo
fUDiRBoqw0eq05C694cCw8YcVzeGa0gI9i9a3E8b+N3iVP7Er0oT5XNv5YkXoVHKfoJDq4jzBMc5
dfs3DHcD+XO04ltlH/QxbR4k9pePl62v3Jzv2CP1DA/sLtza6ZfIMSP2OBpz8HrZk41qJ4NYNnP5
4MzTVHP/U2OTeiTRME8KKqLt7CMPqzMVpf9FC9NzCwaaydbnReptTryi+djWRCuWIaT8s2MfnYLs
sO8L+eUN27Xl5Kf9oR9hO3i0yvkQT5iv+DO+WNN4IUNLdnJ1DtFZl1vqkby5bfG+nxHBXMkNFftG
qosVPkxTg2AyDvCqJ6yNuTmTWectkK7u8FnwKjHzCTZ4DIH6/aU3h/4q4frGopcJyVqwzO8dKtzk
9lBdMThk8D2sfSr65gius52tiUcmnBrxixloDnv6++m9NjieV+BGx1q/1nHe+EUR3vvMClurqJdh
40jHikYozpWiBRvMtbeJhRTyY+tbrjH2WTBAkeZ/Qwh14RSFkk9tnwL9u7nl9479jRzCxYmlPyja
Iyna/A8QG53yyixyXMYtTyz7Igh8vu7cQ4DPKFwl0B3X63XIvvvIW6in6h/ntF0KxU9/f30M2+Uw
Seowf5qYqXOdeqW4G+3Eqe0M3+1Yaqvl/LAKay4yTFnJ+Sqp+z2u2dRNRT1YIn6obZggAvrxKn5N
7JySB1zSKx1VxoVyreDzjuJOOcFh95MXUHUDS8Rw/ACvH2ZPfU17aN1BoTBnj4UGbsUYpwT9KDSu
WEw9yrpGVrBSZi2FYEzM39p0to+T2grZHbEoc4bnjcJF4uuzRd3jA8qnyKKF43nfhXewKwZNqwe/
fnW/urafXYLrqvUbUHRsa7QjTc8O9tlPtjOjUTbHcmyHWcpvxtQF4xvsM60TbnhP99rLb80ZoXQL
Sgity+UBnYwwQpHY7QBWwcJImX8RVl0GHdgwuu2RE8nxBjAnM/4HfpkD3egCHELj1hQM2oA6qxvx
Ma7NUaopVWcHyBv3X4CGLZ3yZgCcNrpLZgitMXYqZAOnbC2l2Dw+b0aX/NAbLCq++rrfb57qaO2P
sXIeMHoVxU1wcCaPVDGG8NaNukTm4udmyreLDErgYII4/yvrYwNMj3Ulht9QcmTIUQqqf7RYKG3T
GjpV5HUcxHr32MiceppBeNfT7U0IJW3sUJnWs3HTk5SUpKz4n1gHVrC4nYbjxLlljcKgiE16cn5W
fGnjSSg/A/zdeeBLt+SZisYVKxWi0Srza1D3UNVNMoqN8CnBztQUr1jymDlcZf76nRqQ9mRSKLmF
75NLcFEgjvV1tpUcf3KtgwNDEraXBwNkSqtyk8cSGacmxvmIk/+uS7K3MIWmlIwKqqYDo37zoqTM
A3p7FCM5toezZKHbUqIv8Dg45rJXq+BR3QSDGd4nOzk7WQ2HBvw554CXWiNn0VTnBz9YqIDbdwAG
8hSOm7ys5gZzpYpPLghgfUvNfZoxeMvO121p6rZsDOYXN7HrhiXQfgeh5GfPuZsEU2HgsNbv1nlf
Y4yk0I5rwzskCztwcUlp7UWT5xEe4Fwsz2negrfa1X4bB8pEE9xvPiKfNr2g9QdnqhMIUAsVWqXX
+cJiQhZhchl8rbjjH0e3w+Z6gjr8tPM2+v0POLeSaix+02IpP05gNRXmsOAmEUbFMiI1lev8bRh/
oUIZCw1yMoglQBvxnoeWIJqAD1QD2I3ZPtV9Yj6HMNSafj4tIx4VZ5TI63W7/CTMgatGo0vhddLN
fbkdzRYJ+q0C2mD3NDY7Cmv0lvWv/1Dd3JMK5G8YEEtX/8Raim1knp4ExVrf0ExFS+4mKArGiRW8
0g6Z5TMzKLmTuBozsBVIe5w/oyrEBYrk5k6ewXNwxjg9QYax6s4A5e0UF3lHOk/l6+1g9D5R7KJJ
qk1RikGZ70FphYqpbCMJXHH0zwFUFiZGXonJHNcUF4EcTIHYbJ1hOVPKZwqu8xwYSP9E8s6eDDBp
ChtXdonyFCjuaqV+FlqxL3jGGQyWXOJaRChlJIeD9vUORDYurLlSqInvCo/kQI51V588+BivK7Z0
9ja3LW6EUZ5HnpuRWNdJiLxnTkdim9cm7QM29BQ0XLNP5r4SBFM5xI/x0NwGcE6LOkxB2L83k2aL
uOozZBcc96QX+rXk362M9zmf3mc8idxETZ5ONX16ThWRZPgM16lxxAjGAPK94GtTIErMbXP1fy/D
WgEhMr4g2M66qpsHOHLpAsRCP63uDGrg7k7rzQpfATVX8UHRtMEyxS/7/t5HHtKk6ki+a3/toTFf
C5gbMLAfUesZaETnov3fio+mhnKvQC87hqk4YHHLbrXICEhypW389ej6MAgtbUSxcu0r6u4cOVlx
1y0cPdzculB+4pkHao7gs8p3X96mllc0QbPYVNbrU8Qq3LyNTw+WJHVysQyFFGzHqZb6zerTp6W2
Kecl17H5G1G7nS/qCyMeZnnu1KJCeYN7aZCkIs7TXsPA6IiSVXiaSmYAQZoORwKhJrZxwyHvZvp/
dW8VlSIwjtfOCZ9xdZvv8icqoKDFVUUZCJmeXaGLHG0OUsAW8hcRQO5870Dr0Tmejsw1AA1GutZC
AkIIothGxVomMAfIoKj2yb0GlQwwRLoUoT0p2O4GRUT6hejw+mnnEaJfEHHL+P9o7tztfsAOQm+x
ZQfhmrxkcrqGmqSdKCjObsCehEYdIDWjmsq7mXBj/54QpBL9Z+hFTx3W2qZeFmbr0K4ZBuUruTfh
AOfYEULjKg6MZVAO67dl45LgVr5z4feThCtKSPFFjP4c1BW7jIt43nRjGMFE2S/VMjo0eErw+9EU
sWVpZwT92keld6HHl94xXtbrHDUi4anNwdt+LKI8TBa2gbUG1OtkGhgZ0L0GKESeAH7YAkDvY4f6
EywHFtzlRK0X9F+n2INnJDTBpYj00ZXfU4asfoWFlmkJxXaTdo8ESSKRJgAxStKZGBhPy6zbJaH2
rhKvHrSKZNaDTTf1rdSnspnyyokxAKq4WxVLqdWZzt+MJFONvS1My0i798rbo+NIbeCQda1cGWdw
MZkX+9tuNPgeFUhGKO02esr6HrLHWV74uQv5zggjDSEYeZv4+MMIa4q1y41bPn0wFCsCLlhTgEbg
iBm3wFgytunR1f7ZeGOWN8P2C/pdVsIZNtPLKfujenZlpmkGmd8Tf40BzdQK3HT+v7ijUBUYfqnO
lUBgVmADLYnQXPIOjx5XU8CiA+/O/QdNHP4Yqs1NjzCCrPt6HWhaGid/qPTZqbaR9URXjf2hW43U
/hRoUK23RHI953Fc88jiUJxFxa0Vp2+9qdCyG7YcaRzsodd3IqE8c1XkzfgjeUxVC/VX5Ef0/poF
Oq744xldgcbrNq5kapD4oSSKKKyYlz71+B33ClfkNfretVaqigos2JEc2T4KkxySfW7ME49okSVn
jmKboV6YbRIz26ua+UB07cmDJ1FTr0LUNM5To+WQGAy6rVOdupkaL7pi0dctIl/6Nl10eQevQdI2
JI6K2YVHRt2Bk68RDoZo8HYepkiX1JzrBqbOAtMlz3cgunEuhGylTMJF934d3cMBk4wUgaZXYT5M
dVVUHHSMxIeId5rDHZHBcxN2GXA2TZpz650gJ292xshM6Ebmgj6hPwS4aBBF2S7bNakmrceJpRy2
dMHVr8J3fzehBUzys7BhTlThKtDvz+vvdDsQtRMe+wTlwBypWa5MoedLL5+obnn+7qasRNr21DwW
tVARCLdu1/xiPdU/ldT9MyyahqygfC4iQLVUe2+B+p6djVALwTQhcAAz2zdZG9E2fuwwwDmj3dPV
PB6WPcjm9PFBUKUmlMDHiYvkhpOJSuvBh1nEkEZFNOUCnRJhdI32ZiOADtaOUfPpj2IyVaTaUOPr
5iXq+mxrVYwYSLsmuBua2VrabAswCmSklL2QD7fsXPF+MSN6rY7HkdE7C0jN7NEUuSXCBnfrQL1/
DBOhWsPYfWMKqhhx0hwhjOpPg30uizJQtvjFGurMoTcR1HCEjkNM0Ov6v191u+Tmavms5HdI2783
01R6DTZnITeoyj9+WFiaY9nAXje4KRDfStLmVaG/NEGJ5PdHoBCWRigl8N2cx73bc/RsFwBmFJtw
H36h0uJT9sXgfsOo/zJCv3MV/w0lyjDQzBTEZCJ85OB0ze1s5HO9MDNvhzyIfSqcAI1hY31rWipv
1KakKMOKRvGsIs6d2asMLt8jQIOO4KPTKqw3opHKZh5POOK7h1JFgSYPDZb7283RkhSAmbjr49cm
WhhprRrHfiK7BZVJSVs9RHvFbcItxRS3wcNskF1HByWGlTQXYtBRNaCWm4subhVtHryTqUulUt7+
rFWGwlaOsIlssaXsa3yfiDXmbnKIN0deCC1WzibxBSkGXP+IeOFjXq30eDYoscHVYkoY03qRzsCu
O9Vdrn5ltHd2pRR13qQTYpJWZVYHiAg2VHRtxTJunPRyyYumKhzgkAdXWt4LiAlU9EX6Z012UExb
i9s8aIUfYMAG4wltWmji2nfzbo+m08WXZ88j1TnIsdvQEteCjeBif0m1b8ZnZrJZh65F5lNxE3TZ
noQFP/3YD8iJFavRU2ZR5y2OfAvnIMQT13raaj0FARWab/uVGR3k5y2HLcQkv3ppG4UweWR3FGqB
zOwS1cXNJzrG5UkzoSIw5knjqUsmcIC3C2XuWlQd/FiVGGqEWp9xRUqXlQmrTL8zeREnHFkubA1C
NfqGouVir1izhw9Df1N+jJ0JOAmqGmYzYCuZQAuTVdEGVsd1d4MhqdqQNr/aIZlslECzF4xKfDC7
Jp6FtE4/lb5lkAcD/KN9NQjN/3q7NFPg4m0mHOTPmG0jtoEmDkMC3NYCMNBDmQsldEmrInKX/cow
YCnyW3neENAqlFt8qEmCheREPzPei0GwBF5xoTFe4x593BD+3yeifca71+QuQn3ie1U7U2sut8BP
lRivBJoji8ti758bA+uLcuxctfqOC5zu5fAjGHfL7MeTbFAujVekxIADSOMT5ph0hwZZwH+gCHoZ
/XZxSIsh5x/c0ZCFfMHCR2/2d7rgt8SII+pMrEbAX3R1Slr/+LVJlmD+yuQOYIkeWJKGkg6zNHPE
rEodm1M5xoZoVFDPLrksTNy2Fk8VUzrFAW4WEV6OziSaT1f3M2KVK6cuka/AryvJHp73+i/Jrss6
EyLrx2QMgJxUV0q1F9W/OYOlq+jMFNct+YP9h49R/08oOhLD8fm5yoOV173hM5fAvoomOoaGwaJe
KysqsTtCcTOeBbM3xYIPaHmIfdPySHis7Be+iuu07loGTxCmvBoB6H9EaOH33T7WiQWDMiDORzDA
WTyw9do3v/oFYioxWyoYhy9y3ehnwntmAJBoZ9htJxcPpIa8t7HUDhDMD+CLROo0PwtZHIQxE51D
+7b3qxpB5D+ni/Jc6qefRoqLXdYjV5dYB28N/zlcT0pFUO5DCig3dwDqW9ljZt6PKfPMPs4lpms0
P3whTvS8WKG8Ip0Gf/XrlYDb+3H2703M4mdlAY6+sWLK0pXem4bfUdK6BamzpUAVlO7p7U5pQIs4
Mz4mDE7COePd3rQdeK+hKxNiKL9i9YgevkY+arFp/1K4VVihWtoBzz4nWRbFTdCXW4K0hagNTMuH
NxIGc8aJNSOZpmm3lqXXqW2ATKd/PUrLP5eufYq79aUqsxVyXL2pAdxc2hF62Ftdc7OIo6YNigso
yeoyBxEmDC3Sy5G3kaPpt2TkadrxwSMvj+GlSJ2wjpC25Bo5prOg+ZLIcW8pbqjAY0QK8nd+dFgy
VcjiybHDRUbLtTJm8mhkAiwgXVM62K27pPOdl/QIU7ZVgz2KAZvG3OufIrcZr5Drj6c8O37iQEEw
lo1p3yZOMKx+w+0pYBw6eLCQtzOfQrf4uq7py9ZI3IQ0XMm+k2AJ3A+grMLcwN5KYFQEf2WJFa+8
gKwBQVv/xm9W/Fo9bHT/3goU16Uz77yzq/6H7Lj7wJNXbBBPiBDAmysr2DO/BQNrlX2K6cwjaE6d
+LYEpAjqpldWEiVKaXBYrelGAc4tdu3zxAmHsSESzOaCncc10UH6l21Kl8PkEUNmwsM+K4wec1bj
oxCBZHFYSLaYekBhatL8e4AJ5yOqGHzLAdHdoKHVLjOcx4B0xFPOjk8sobM7pX5X16DedseFaHnV
jh8iQdGCPPPls1Tm5gCva83ayi1nDefuZ5CQBHdM73f61u+fPu/EzfFo/UzNcGeHZ1enSkiGATvb
Y/7zFLEn6tJRtv+2Bkmfw5uEAUfbEqh9fY4vDHdoxVMxE5AV9i0ahBv0H9x8duTbxG2c/2dANEyb
LkOSge+UCM2kzG/DTp+WDq7ocQbANje4vLqAnQKe71POrRK3PRSc6kILGG949YF6S0Y38jAUiZeQ
zrRsQQst1NYCDDg+FsjXokj/WtZmG0MEhIHaKayp9gfVM9Lud9eVovQ26Cp7NJyZsHfGJ5lvF9wI
DkgBd/yOAKfQybfnUnHBk9/+QrMunuSFaxlZWHg4phakMOzWOLpxOV+UsJg68tCOGQlNXT9MBTRT
YfxvYX33eTbFFKxjNDEyz8g78cKohKk6QhUXVKr+FsHf2CCqsHAfM6QoZTV+jCfWv5DAKfNPGt0u
CrnOEEIceNabl6tUl004hbhlunbJWo7SuXyZs50KYia7ofjyUeiOlbbFmVQ1rW0B13pIb+I2TpyC
UAiNJ6fzxUBpS3MYoK0gcgCtgF4Fk/ga1yBYIKRVZElHbuHgJ++nmeZIyYrwL4zs/KiA2btEvylu
/dKch6jp4MB/xFdKVl99leUJPT1MZryKoL7bhA7szu+Ql6z0S06wIVa3IcpOJqvbTF1g6Obcb+E0
om4WKqR5bOP43QXO/jp/igF6aBH39oViGG0Uya4Ze8obPitNlFSjNVKr8fuuulb1Lc/Hf01KoFTX
xzJg4x0CkgykaUPn2GjYnUDkTr5OmacXbhgnOkBVu5oITjA+cP3NuuBClOAacOd+3GsJFeg5vR6m
GELmsac501QGSuoTnVPWOs8J4boG5qJXzjnJF2/uVpg7PdsrEgy4t4g6fRzAAFFUOyzvfhQOBz9o
orsGh1n9XCK8K9nu+JXjm6mNIBQyYxuf55r0wi7EbW9axYIEt7NeKSZZW5vkmvmVB8DCjFI0HVp4
pGYrRileyL263uZQY+5bayiDxQ9uK3Nj3ITbWLHBzEwry/bZpkbUZWHZNTxEIMXXeqCC+ia64scc
5iwbx4QDef/7oyO41QLKYfP0fpCTNZC7zeKkzk7Lsg/3KAWHVHt41r1DntxgDDRCdWCfkOdlKyRA
Vfi2lJmGBFcUAy+SHpztHnkLbZIqQ+3cYRnzT77fHjyzRfyCWXLMYVtFSBVfBepj32uVKQijByZR
QNg/sh5UqSoqNyUORE8qrguRbwT8IyXpagFrSfK55mfJymnHeKV69DkMmoFtUJFrh/RhtWXp+10O
/0WuCqj/Jj73vWMoFiDFHGsR+kVvPDUcHSH7lJFx4Dwt+QbuR7Lvw6FPsv6u13UVJeC9lMf2AFVT
n1e/7Am9/Fnx1WqklCkIN2CfAzxkPFL5sZtQgl9ZS4VWvyUuu7wN9bueF3O5ojyy1CA/UuR/u6hr
4Nb+ym6tD/8fnWIMGWFvCguW3Opi0ijw6Di8y7X2NZFEEsDgkCIqv7TTqXIfQoo51cHSnxLLsGgq
z2mNUAMkP3eAX0SLAnmwUWEDxqTHnF46ZdZrQCE2KuGq+hJBLa3jZjyI9LhKu13UAMLNGntsYnM9
O8n9g/n1Eo71wYvqs0AtC9TfKnVlxmHTDYXmdYRtT/dj8UzB2YkIh5j+sTdYC3p1FwC011f5/aTE
d76DK+yIH1A29PdP3Zb4RyT2SU0KtxJcNrRkYKkxErzuM1/SMT7Shxw4sdMFLbDoCNyZhQ4Og0wZ
wzPw5ErJlyTvC19yAUO7N6tshLrqQkO5ODkjNRvjOwFbvvgmYJsU8tLCz1Z9/5SxLwTwfYkJO9iC
uYLGjswtLuFWyDog1GhtA4BGhP9Y9VLe/x3PCQfNKQymauRQ0u2GooGoqSyIx3tPApr1HSv+uRR5
OpH9arSOtMN64576m9+nwMCQkGRQOr6V/nMXPK1LR7g4Tm4HEgacDOwh3B7U22gl3v9Bwqsq3MEj
z3snViqcelQgz2eccznXTUSkTB2QTdMqZ0jN2H/oQSUQlQAynWpyBRuzn+SiGZz3f8Pfa01IhRFZ
NuUCUkpqdXwz+Bcp9M2IRBkjbyrElmJEynPX6ixZJjbq2rjpyvPnMAC0Vkj35pjIUYINwbg/dxDF
Knlj0YOZB1lbqxHT6+IHuCCqjQyQD5WENpETc3anMliFD3Lg4rS3g5CJTq/SyG/ZZ1RAX662bkYM
1wkqhJ8kPDcx55XtDedR9rzjCTrC/BOvYm7bsdrp2i38K3o0GOt2B3fSsT5y+U5uRmIcP04r8MIg
YJ/atuyZE0t+VDjRdCZDdZ+/r7DziHAy5TRjjL6ubCTJB2ykMEbct/lFtlk2zDD3VJwYDP6I2kr7
x/0Hk9F/t8BO2PszeGPwCP6ckhwtjudu9NQsZVuzsp8YPgVyZUmGcc5wy4LQ27SgSaEgr23MQPWB
H2vhJF8cwyUt6GU97+fKOrAE3oPLZUFhqHm1jCHIM0uztH73Mh81T6eGFCSzQ8QFPKUiQaz3gKE9
xEJQWbLOjcmrIaSaYYMJwMveGxeVrZgQ+7V6TPA/S6ESUKj5iR7pLsE06csHjn+eYAUZazh1d7+7
1GYcbYFORUJk0IU29HAN6U0v99OhuyhCQL6GVBwKW5GxEf117Q8AtQLJGO4C7JoUSEBee53twBFW
vc5CqZUFa1kj3tsKn3/IYqW5LDSo9o5dfakTrMJftMhvlF9X9HrC0BYmgqEY3l4dSSPWiwtSESyd
oUQd7XsxSipMBPrhrkFOLcCN2vGisSGuDSqBsOCayuGWAVnLkuRvzP0JT4n/bVMnDTC3gTYbp2+G
7qm3hYWg1NKXnwJ0S3EUZlf0ghmsmF2/TW7aeAaSdup8e6EJTTQNxdybiC6HmxPrbnZbgemCp8sK
9R+6gpB9IfJBvrciFSjBJL0flNSFGq4K/XMTmPuv3IV67BW/5s3PsIdAIBfclPjQgkCXev+NuIdI
d+DR48Nx5/DqKXRLxrW7xncrFgcpVt9zl0YdjzNqojWB6sWYF/MVUDoxK4GXalWF8zhVl4u1pUSv
nGD5jNNPpGHtriyD1YbRwRb0rII/GCOpOKiWtOnFr9rl9iHGpKGS39PzFUk+v5lhT90wCTp6VAvi
zx4oRm0zQnD/xvUq7l0Pd6FCSQQHdMP4UAnHnEzrP5caQx0cRptdGaHXRMRaBZuXG27JB60IaeL3
UDl5wXccXIVSud1Zauwh6OE/Pzr03ouW2/XvqQsiQ4SAwFrhlCYRxNLqG1X018mI2/J6BInbubjA
abMuoR4msliucDe4mCOGI9SYYgdCMclOUUTirsno1AjOLrSquRo38hg15Y0YTZXcKRtunhOaW41P
xi1UYkA+aIJYeX74i1Ve8cZAqywWoSwF5LLivHmEm/IRx7umacv/TSV0ohCGyb02RYNRAwU0gq5f
MY6F1/1QjNC9TubMx3ZQBaUO7gjkxgfo6jNZ/TiP7atr1mqs6jorHdbZMB1/ldrOcB74+BWg86tO
wzmmqgNrvrViN9zYRXD16T4dF+DgXVnkMRsOI8YUh4Gn1QueuQGRzdeWbZciumLEYJ7owjMDoC5c
UzNPlyO2ekVXWi8Vw+JYYLlUBPWZFCiV45VyhAXM6lYOUIgKQhYzpsDNZ/AeN6dMjfG+Uf4adaXn
IrmE+yXslswKL4eausuBuqBv4yNMpwyfFqVau8e+V7T3dULyCIa6cbpu3pDjmUfXOJMqB9e2cpv3
vVveoiTkCuZ/wLNiR0KTn/Eg2RCwI7IOIonD/ir9jyy0M9+7Y5ClzY8jgyz41XTR9GIytDZr58NU
m/UCUIO+0vvDdGr13cWL6uhf7lT0zMiRtDWeVwWpezExO23fy4f61Eu3rGdpsU/yZA8tJ5i+AcAl
tJSlVg/UszzpkI7mnQ91blpV0CTWAbkAd3u57xiBRPUwUGIbZJOBROxUZWYtsGnICpXEQ+QIqrKs
aLDyuC+H74Ufq9b3Dai+1sBEYAP63HTmluLiG/dnhM8c5wtXWWzdzQV1djMsDEMMKBUGU926J2GD
s5lPRNblUc7CyKKWbJMow0vZ8Xfv6iHutqoiEftITLYbeFUFsUdTAy0ezeo0v+yrfZQf2THJSO4w
IYXd60XlMq0g1ZOF+W6ksLUo2afezcWJz86RLOviL6SzR6lBCTXv3axzG+XAJbhzsBIWqRWAosVL
RoA16yxDze75IGwvT7v6dKBQhgKs44CQH03mWFvaZY/YtU6nUvgJv73XfbRwEeo36eDJH1GQA4Hb
Z9YpTaEhX3bkLnYCd6FhPU7MvT9qp7QQImccKlY3COw2GVwK6IMgLc6xo6/Nk/ufYll4E94PldEm
JKlfkLffRxQkdbERANPeEAjtHeZtYR1PV6xuvkJ/z2MLu7QdxHbnOg0QnW4iLU/WXBhwbB0wKq2p
pNY2ESOlwGnjEXey+2aXS/TpLoKZh620wJvQIzSlZDGqg57btRFRZ/pJsz6qBi6ihnaz4/sC5i1p
DR3lic62FOEUekAuQbfc1ZwSQ0WOXDkO7jYz0kJSJc9JJ7KIm2JCZRbwvKAUOvnVdSS+KHg6OIXb
Kwl6kfBO+HDAdtpTHB2yDuiK049svaDrqrhHyp1APqJUyrCvdGvgle2fRQOvVTVR6ZBZFOMTha9d
i1RCyH6nFWRUUNYrz+t/exKbLUPs++e0ts+iunqTq7j5dqMHFtjLvVcgne93o+b5mB0zhAMhHfNj
o1cHuRNZg4R0BAwdwaFCKsqKyy1FFWkFCeaUoZz/SnN2d7O8GIxQRevhcZXwi7lbAZ5wubg9m2/T
NWtd1fi1+ytjbfO66tyQ6tpGxyoDzGzHf8tiTNXfSVgubZ8Y1625msIsxkoXTXHkHTOiOyfebmi1
j7dMuhJyIi9fwYtJ38vzfYoTJM5DQTX1rvYyzcUGCARegM8uk/z6IraWbs40jC6MOmdNWjRzW45w
Tc8QwQz6lg7He4Vd++7Tizcd2w9TTLteYc8oDBlSu6wYAoHrJ+sxg9X9VTrusESMLYieUGSk+YKX
D+fb5PIgID9hJrP8sgAlIw399Pbuq+x8q8k/uwIkjLHQDrmX8LgLrwvTaDt87Tn7IWA4IF0amH2Z
OaSKnVATlo5OKAf2SfEiXiM4tY6hTe3tUWT4+nY+EUpmwNpDB3cjd1ERCnoaHJB5ZFKkD3m2Sawy
Q3+fsEjuMYfkgEgDEmen45W+E8IPliD/Wuvm96/5qxeChf/PhQIqbRET093aM+cEI2xoUyQDKkaU
zDjPAe3h0+wkYIoU+d0d2Kmzq9tnttc7zvFOoJC8WlaQt0tul78ulnpD1L2q8s6dwivCaPJGLVL8
lBJH4TOol6XjgKHxoonxWeTucIuy46pshU0iy4sNuM289XPwT9Lp1J2p1+Gn1Cm0IXA4loJusReR
OHgBTMNWhFT3/PBKVeFgbCtA+lJm0uyW92TxvPH1KhLkoO9LfrtBHWtaGa08HK67edBLoyCqpJmZ
veY1VdhJNNhKHYH2++bIBGk0jKNxlXdZooUOOSpljSkndp6me+l8QFfagpDI3UbeWygpkZIwRg6Z
bbEg4wfGBiajFysD2F/y0WYDi25/kJCUhgyS5vZwuF1pKOkhnUChn8clG2tyyqvSjnPv8dB3JEcf
wGm137o6TJFxDU86cAEkDHtJRZmFGQ33PLosNkpFRJr3X8FK6tpreG0NyJI3mgJWMPaWMrwBXBWU
gfP4uAE5TDQDVoSswnoICngBAsqxwBvEbuHXrq5oiXh0qpAzbEfwv2qCie08KNuKspoGHkoEg5x+
qDkms7vxUW2rJRHR3rh43Fr8TwyXFWu+4CB7eO00hJ+Xzl1nld0g+lj/jK31F90+oR+iI8W/Fd6o
nboTnI1Ur9vjBN5ZA1WhaRjz7wGrQ1L1PEWoysvrn277E9lygjeKva+nf6HcliaBLtQBzijiAhiC
JdoHoT1YzIJKQKR+gkXEXFW13eNqd5RSlJzwLHzsYP7PTsymUIigjoG3wsxYSCsf209VXjKZ31z5
Qk1t02Yy5gplOSqnWpR1cH5LeeWoIyBCEOeYD6IRIgYsGKcH4+zKWrGh5lzQxfOEk4AKnqiL+Wty
6rz1yNq5a1+5KgZIG/v3qR+e2buXEqJr1WYQFFIMCiqvjdcIU7c0lZZTtgEU9R0CsQey/VrFePIL
jDS99wLScnIQAjxIeq1A/zzT1QdG/iKt9KXOmyShFNFyk77ZsxroKzsyHeGbu0qMGnB5cyJeoLrj
2q17Glg/4+IpzkKnXYo+YRUnfuo/6QzCthXRC7Rjdrbcry4WowQap3zDt6DFD0vu/h4BwhyDZLFN
idjixkHFjjob/roAMi+nwqgxqqlpnVEQGrKqDRVwkL0/duHj5j1zh1un7xzWXYGugRyub86408vv
DEbssrXQiQeIdHtkHKXWBtJWPHO3ZsSoqnjMFhk7mbBJI3IWZRufc0jhdrY7iTSVLzRz5ki1abOi
On3z8EefOf90MOE/3fjtwMJPTQFqCkU+xKn7CQDlyiEvIFYgPTTz1fXSSLcD09JNuJIJfb/fA8wg
2eTjXhCBaOguElg515M0aJ3Olhcm1C4bxn6fo1JA5lXLb8bx0E6QysVzo7XgGcICWT2jR3xiPmrm
QGmr4AKqwHQVVbHeQSDeYxIEUKY/csEVVhrmxtJrJsdIhPnUvmAlxGsNvYq+5OmHfsP6uulv9UnO
Y0HI8MT3547nNG96IAmDcYq6jeGthf3RGT87Mbo+KiLB1DoiY2vSaK279QE9lijOuZC0lW6yHlZD
XsOWmbpvf3dwHVP6+WJ2FuzIx9drYGkfpmJOzoYRXYK2r5lVYhrJJWqaQCyNDsuBd5cKEMJW5cnS
LCU7Zx3h6mkpmP6UKS1kcKvz2b7UwRPlh7Rh28NL4F7gGvtbsOasyeC2/vOmQUCarsHif84IDgEb
VN6ahs4J8OhQrpnLTNxLzCK+P5Ax7ebCpfWR28tMuF5Ceik/4kREb7twp2+Olvalnz8IWlH9RK65
QgDeL7kffhbZVG/AyRbJQYB1tP8pYDWZj+/fmq+8KrpgKAGyAa5+H9bAnCnYNm8b1sQS7zYWBAxs
ezpCzo4cfkx+ts1/7Dq0RSDDdK8UgieYU+UtNAgKJpqNRDOl9OwU3f5WCPW+XDMZ31TzOKBhfs54
HMmdl7jbPhugv0qJUsIL8XEUfzO6Nckbn6FuY9L6eZvp4LEtLtwzvsNDZ0y2DHwav1s7DU3/CBk9
azUWNlq4y3fElpqlEgOid2fDvo/57dEz/HAbRBO9nuv8nUfokjrqFNEZJYzeKVT379x7G7e8M0NR
9Abqw/wqh6Mvibg/BsdZA+o1JPQuXKZFGJB45Nw2d41P/EsPQM2981c2mOIbL0VJ+o48rcsNadap
BqrrK9hPBsTuPpnOnKxpyTq/ISaj49tJWE3x4HEE3d/O+wOGs+XeJ/IY9tLCicoZIL7pAa+CHdiL
bRkJFCiKv7a3NTdF39kqHwrdvM3azxf/FgIqFfT5B2uD8m9VVuZVDvZBxQPaGU8xo5iC7dQfKpAT
B8FLZFo3nvAbFwrgEi4nvTiiWEjH7enC0qYyZNUGlnYyav6pzQWjf87D0btId6CcE3edwv1vqMPH
XKQgjIEeG/aeerLbUMgF9lCIsRtXI5M46FfLFvmZuPbJGHr4bZKCz9/h2CXzgHSUlY2UTUH5p7GU
it6MUDgIgCVlkwEj5JgKsP+d+yWvKESlam1ulXWP39rDE2oO9eQr6g7UnFaPMG6dpt2mghsoRIFE
qqzU9L71FX8YBT4vWlNIBHnciWLCEdypczGZmobzxce0Hqi+W2a/pt/j3AqJEr1SpnkotIH/Umhg
Ip0zXzkPGZsihPkj0pialRbaLZPKJpLVMjdp+rInctxHYih0FMtFYPfYMIv4hbqJSzblOGqkwJVk
saBP5uTWQMRl83BbAkKLs1krMpWuz+E7Fb82HQSGRxl1GaYHJMWI5mHF0KTnMoGb1D3hpQUiNJzw
Sw44pXr+/QDeiryg3N2LD7QBOTrpA4TEe++DeCNn3RR7bKBOzO7FFQseH/mTSX7OyNPI/uo71W7K
eM6TL9rWWmJ1kgVLrTkUkM9RN7QjmAJlcPCxs5rLRn/zo3kKdu64JfUrYhsjWI00VYWZnU+046Lg
C4fUaiXB9+VmbSo8L0TOajglzTMlQuHl0z/8cFimhfXGQdYSEfYPtysQspyiSjWKuDwm1QOOkLEw
+v1Xssho4md1UUYsfljGZbARLqEzc6RJir7nFPLqnmTba5T4w488HZDQBqNr99ZwuUVmxVptscRr
D09tjFKrQCGrKxPz0Oc9aFIV1OowP4GHTiGaRrOm4/l4pjT5894vHjjI4DM/PLtUvnz5WVZAXzvx
pyBAbRnWgBsXnslJot5L884tqAoVOMfr2MS9R3H14XaIXhJMnKpTu/73YxMPMER1osISuv/OUO20
c6DfyfVNgX6DC3XsQ+KWBJa8jdEOxa7ng3YCnPj4qeXX0eNPxoBXLexp6CxW7A8JQyI3RjPP1HmC
F2CQf9mwmIID8hUUMwjyYDuAoXrESvhoyYWVk9Ot1B/qm9HsovMKkHiOl24vCXNRfFHHLpPkwS6M
DzwLXQDC6LYK125+8msAdrfFBESKsnMOyXSxV8mt9dx6sKmM+cQwlmMo8UNidOyAHrmI65U5OJwz
j6m0pEVqzDMhwiO3WEWdZoeaHukSbmu4Dv871zZj+YLBauQ+hMAxSwc2m5WcGU0LTDI5Wxi3INMw
33IPvAltv+CiqZM1Sx0fkwHjafWPjPi7ciQ2FgZaPoEYdbNj6dClTTIWqrF/vTtXd84g3wF5K/uO
cN1AXUBJw7O4mh9+CXCRJ1LtGcsih/M6pRokhJGuIUA85GQPifHFC3A2T3S7kLOAdWSKxfOZsvFW
ravCuOBCEJM+CYJmB6ztgrVx4Z9LfkybOuUEbxcsO9puYeXhLQE6hjDELr0siTlyJZuiJdAE9M1l
GmkxTHf3OoHqsWMSOVMuRky4epGDxOaSu91w8jfX7AX0syP9u/tnL2vjcMdoh89Ik5+HS5T5PrXA
P2XEvDll/A5rfNBXLkFcp5EbkqHYRlfgIsnos04MZU7vaxZMAv/Lp0rmCsUaynogB5pYRGprRvLL
bSf5H/FFMzz2peYkrBY6QmDNfBsC5yRx/XVaFv9KEtqupHRKRX6X7tIfpZp2Wq7cKiw+QUk7ogW5
1JdPWGZaT+YxsjkIyJml7HLKTJsYHqy9fXpTeJ9BX8Smhxl+lB/fOxtPjHSNR9KKA6L9Ykk8yggp
mhcOGlRDp9H1R+LoUzDM/qeiHDY1/XA7D3VV9/BK7JSVZXswv9KspEU+TxrePK5ma5HifcI+QoK+
OOXRer4h8gAH5AUk15VD7UemgqG7gQiHbljfGTcNT5GMm/IlOEjTLaBNWu8J5uGmeaPrJcZXi8bf
1wXadoeK4h/oF4imv5pc9548ZxWXkjoKhvJdpVn7ITDwYRijbubNec9Up3wEtdmN32J5UFQyhEpr
M7DgGpWWDqyKbTnVMAjoKGkCl8+fuq3TzR0uKs4un3ABPiIwUrn+z4I+wrnNMa/BmNoAfpth0qP1
ipXFrdz+Z0H5QgAFRcT2ZQhXPA1euyb6oTgONGHHpO4Ee2Idcp3VJwjUBTUnQZbZwcXlR52UXyYg
q81g81ozZNbvbSFygyDEA4VO52QMY48KXw5tZJE3go/iBjwHFoD4VxtOw9a+4mSFWU5eIZxTmjHf
ASSxvr8pMNjb/RyZcpbVAcyCmnnix0DWvq6bLyKDlWU48bR4s1/OkaywTwz7yf1DbeXswSaB44gs
N1pDu92hG5uvcUIavRIyO3zsxEeifFFTXubJCaRa6FtYuwgBlaFanyWnxyE5hUGmdW7tfvOk07Ds
gY6wvq2/yeMI9VFhHt9DoVo4S0otwRZxOPRB++5pwDTZmiMJk1Mn8p134pzdJdI0f3omEUtbSShV
4IOA2hsDbEh+13J+fXS84XsSNrKnYRugV5yh0rXg+1qz2f6v85S2Qo47q00+TVfHLokpdbBhA5lE
RiI2BlZMRRcwXcxpAmJ4o4vZtUzxUymdFXxjn2ukVKMge8zmSKaNQLJhHFqYirYE78ldokFF/psZ
+8Xj1YQB6vsvSUdMN+zhkSlToF1uY9bKWPunPSbmaZOC94eRx2wyLoXUWmPC6UxWI5yYRduds/ZL
/lgzlnNVBSlbSZjkDQZJvZSrE0CYBrQfPp2gfIxHnhxuIIc0kHcBZHFcXChn0TJgFE5IVkodqQcl
QMpXSP402AI+uLePszLZuMm9ydJIExbZ5yz/EUF7wAO2boL1XrntuweAr7v/FWrbRRmmDqCpI2rf
ZixE9E9Pyh6G85QV0s7FJull4FzPgtcjJ1lhN1LsG/1q5cMAkbP5np+mGnd01LGxXT6tfL8nwJNK
59UMCo6ymROeErF5jbKlZHZ+x5xKtuvdtZx/Dtj7k7m40qkBUW3gP8aSpevGDfxRRGvn4TNMmO6Y
X5MkYFwiWD2sjXzLMFSz2uoV4qZA6r4gGHGucYbh9LabJRtQ3MzDJ7yidyKUK75YHpSf2ReAudHd
LQcwp6OBKA02X4WxCsjfboSw68kZW46jFoBxyoP/fslKMvqVWLWhXw8F0fN48WuHN6d1BYc6wu6+
M1I8n29vazw+2PDAObJsmnywl+HYz8rZUKqmVGz6utFZ0W1LbEWj2a3KLRYKfGVCMgxgfRpXh2Hf
UHNeV7WzKDkDjuxhPjXgBwejdwCjjygaPBDQiS41juowoMaUqtyt3aEeOQ2ekPKcpgFcZKPJl6Sb
zPBdkz+sh1gaA6mrH2DVrZ7kzsrJNh/cSOiRFR2fnF0sLvQOsM+h3a+NrKpPqCBZhlXYSnFuOYyP
JmjvnV/iFnYcDfjlnfgHCFsVh278UcVpkbTPVxhaUU9EqMUDkUTYfyxgbfTEPrwEX9T9qM0l0lJb
Xn8KvPbF2tHEPNttv6nghf/sFckPFhH74YfiWH9fezId/HqS0iEvQfk06tKwIH1e/gWIZqVkAevM
0Mn58+gliqEH/KlMAwwT5l9OZBOD7WsXPiPLm/KHmjWBIY9CalKyJ+qfnAc02QO6c+PHGeIAAYcP
JW8K4dUDAcAIYcIVRgmE2vc3AHHeeUdEh0me+0gz4dY2yCmELE08woWhnBbRVfQkjS2uIZZG/k3r
B4vj4kG3V5uWd1J43tRMT9sPBXDiPIfaU7Di4+O7H2UOUHlmvQDpjLVQbKXnqL8YM8fvKL4H9h/u
iFSBMOySz7GwJrVDo9ie/myYy53y7dXI74UCQh4yAPXQ63vExAepAurXyALhVWCHnTSPhvsfQSzl
Ssf8nB0roTye+Dz5zZIzvIvDTiQQ15SfGg01plGSgByOMMRfgIp+v41wxd0s/wEaZaCRRKEbaUVG
UMJp3UnPWZT2BQ3Hm+InF3XVR0bEp+oGG4uQA/S1mLik5T+Ae9jy0PJnw4GDJ7PqbIH8cAuhduh3
ypp6Hh/WThAZU7VgyhIPzTMwTfz1ybVmyUhf57qgihLI2HbUN1yY7BOmYHVxBharLBT77ZaPWvZa
dAiMrTueZWp7L9OxggQsVkj/+TB9xeqOhFRutIamrdhNE+C878wENwscWm2qzYbtlBlO225E4co5
MpueOqXRp0ewYUC4Fy7Qu+N8NG0XEnP79VD23wy5UQkY1mwjxxIzqOEr8FAfe37lhD8ZJQump6yY
8vD67x9ePauq/qYj3iRI6ckh9CJhU/NIWzywL3y+BwOs//uyFmAf/HIjVeKRZ9mqxNqhAAQYq9EY
jP4RSF1xB3B0evmGe9eVrlkURWMG0j1oD3gjpBsIRxR+7EUDgeSd7KEhE9mge1SZH9q0UMzJI1/F
BfCY04867a8VH8znF9ZH2eOdKR0OlHHNoJ/FrOz7f2bXNZYRieWlu3ObfOqQ+c80v3Mx6RJOt/X2
8+3jtc33inB3sKjZJU564NIUdvUosNrr7pbdwRnQv3UlPgGtYaYYKiAZN/swa/QTGuAV2D+Js0qq
Y6b/rEi3T8Smc/k5QWWUxLAk6RYoMhLkuyseM6+WTblbdfknefOX1GqSHYkkSIkPO7xfU5ZK5sQs
HMMB21IXNhff/Jovou0qM7oW2lWMhIKq7tpukLIZfsmm1FLerG7aX+H88+I9ORv3APwfkprZEFi4
6DZvmwiPM/5BLq9JYgCzGHubwLFpQ5Q/d8NJwFOjsPSc8Xd63WC+vYj/mqeBNxGlI168ZRGKIVIa
7i/mVZHW+j8tuEBcApaStTdT5KpV+AWfft31f78Ibue0/IKHXkSwymtd9qgM95/aFf8w17tLAQmZ
hzL5haZ4pVU43g5EgwDmMxKTVGCELgeEm6PrpuEx44vqkLjAAdztOHn4RWQP4A0zU2NCXwvR2YE8
t43ULRzS5AdGLm8DVs1YSCilbEZRL4gbdO9a981InOCuGrnZ7iXA1sSutd7TzjETzOgp/bqWeN63
im1jo0nD+kaSDqLbriz9L2PxEvDYFnKTuvAW6nqLOypSc3Koe+aJ6toq/SfKdHdfzKQ7c4U7XvKv
8sPfWicVSBqhmbCU3zUNgl7GNWn7W3LJHpAvxt2Nd79fkqO8JVTVBYzZycgW13lVxVsCycz3X4Gp
sOFvV+hzsQUxKwsvOHg4djbWbe1x6Xs/ndq51DtUvDvQYg7zEYhnVbBhf8JLxUcuwfuRxMNRJJS+
W95AbldcZQuYs54pNyHsUc11hfAixUJZB3+p42wO9Qdo4l6LEzki7tAEDeW5QwM7NDzDHh9fxNOo
gQp2UeVUS7f1sA1aY4Ma7v7tIqnXzxuHIV/5Mtt0/UOEP5anUgX5auh9+NVLx/8o5Qymv3dCUW5/
tgJdvb+ZKdimHjvTrIuClAcBV92FcPHbiFOittcyd6bc2Lj/b2kIsUBPe6NS0YSAanIfvX/KZAp2
oCK/c9CDApFhOKb2qsaGVOGh5wYMoTf52lrK3VZSCIKtoVoL1oZNQ3rxTzIc9iqHn9brX1QDF+XX
zi6h4pL4BtmxNoeAJ0J0JRK4+dC43OAdunB0AQY9ES3ddJSjSwoEVahjYUmU3UKhperhQUommMlY
f1COOLgx9hxGQIyeP1/sGmW6zRUyNYPGHQT8GB7NUYfLsqi6LTgB3R6/OkkOzxdhUa6el6LNgpq3
EcCy3d28I3pEbgZtl16KqWti3MiPdX+E1UGJEYX0aevIJe1UWBK+cOvmgq1OPNODsVf37gJlKBD+
SZhsPXCXTuF2Y40hts2drt23H5cZvf5TxYjZtZvY5e1OHQJ7K7EH+QJl3Zsx+hS3ADndWQC/imsr
864b9D/jK0EHOANfERunAozZ364W3bAYsNsP5v0lKyP52xGe2AAO8/teiFFBpR6c0OQg/zwM3suN
5LQ6ELgoM/GBuxrLL9l9aXIQX4S5VV8kHesKxlzd0K9wQV22+eM0lG6mo5gm6b5hngEPkzvjuYym
nsunJwGZnEToIelwLJ+5pAgG8+MtGsqJqCgFV11Sd635J6urzdd/yEwcFRmiM4Yp1SiZkFzw5+4E
qGq6FjfdtmX0ak6EL3JHne8aooWKTP8AdLMOns7z0DMnYU70eSWAw3kWLGFhP3WVtZ+1hxXmsSuu
cjeFMd3Aq8gsMfQN2netBA5I1KouWQ/r3jLe1/FaIaQcxAi2BWBC1bzyK2dLF4rzvEVRKONJkcEW
TjyTmGab6UxY7r0EnI6GKTyLKPD4eDS/FtxIALP53IZUvkhJFH0/uqEACZI7katofTOTsVgJiDoN
pHx9FikT5OvyScyiGXIxPpzDo9l2RheS8Ejr2m7qS3hIQtd7C2tVyDr95D5ZDFN4y+F/ksf0SFRZ
zyuveLO/V6pifGycIMYB49p71PlSibwuoN9PIsXjBkixXcFyx+liXqceq8WduSL+N9CJJwKFkFal
jtOTi7AG+HUc41uV8kSShXaKLseSuIhnz68YMH2QhueVg05K7h/hbZXnwSPo42loKp7JZhXNf8Va
E+9b1wD2FK+/Un7X6QF6aYhIwCuldYt6uSnq0bak32FoLKoO20ylIFxNaE956BioFNRKLaNzSOg0
+6/b9Dp7NBjgYPVElb7af0qym2DwhJhbVHSaqeUW2/+steWOPOU6kZ63lvE/J3/xpgvzVfTkDEZT
qxFsvBH4JJiCj768VErOjmh5KNqgA6lhM3toghWsMwThr1I4h0TWSqV8rLyGlDLyCvhVSyGONiz9
8ZTtmR1QpPrjk1hw6OArBBae2rWqRYTcuWqqUBphkNPkCo5IWAU8kQINhfVLQIL+knQdElrh1usJ
vqnjg5KnmNMyu6RbWMEaY1PoJ+lS7+ueQU07pxC2RkBsyMrEzD6BL83vvsQdwalJIkq1P9ezCSfo
ST4OdpTdoh/tPA9nwyyngHFGh2FFEFwrNKmAi1ZUZ2NsQKNem/CzP6yNUyATNohzTAbTqfYLA+o3
mj/LFzgj3NRE6EAkWnDxuP8b079YvL4GhCFSHdEOEzC9+FI+3y11Dx68Py5qRsIeLccq1nYUK4r9
f0Dxe4t2WKwToN04Ffn+sDWyK69xmaYpWIz9i0f767D+9EP8wVgfLY4tbzjjTKOS26UyMP8aGTbZ
MJ3blxfeo2qNM5wXm03H+BDpzkps03GPvykNgB6k7mzFpjXyl3wTMQTnK2c7I7cHj+C2bemjU1Lb
8yaSV/nSQa9ldPf/l4Go4o69t48jwydkMgb2S9e5w7OAl+ENDFbEUvlfWL5T4uKM7AnBejgT035k
Ao6lC+gjCW9a9Kq2i/90KoOtYfz95xIVukgUUH+kDhZf1tB+To/VSJyv82yDSqWPnnr4EOqOSilq
CaXUg4JvhzsGuyV+9HQ2UYUQby0w67bB1FhmkzmU14caJBDFXv0xkRyrBR5k8G3NtL15zloTguMA
cBDy+IOmVVMb1UhTyCxrJ5CMsAwx6KLlPhF5L/MY0blWI55idcHrdL4cADFogaM/NWtV1Q7bXKGi
8qcLmh1QrPp6W0oV47EllZq6LCs8JnMn4SmzZ9SX7srnR0djernGPCqL8/uwNxexjO2pJcdtLHHq
PYtZ7U6stqXl8+s14kFjerpJiLfDfyWyNcAeQPtbS6FHhsO1txdPH1YFt6mKkfSaP1V0EmN21Q3J
GmZlDsnXwLbm5cqKJp6eB+k/F2p+3L+g+8778EAxCsdA9jBHtlX3mcwLQ279o5GbcqgkR91OPhvU
i9tW4n2TFkzflWhXfigInqSdTENupVVbOpWAxSCccBU8I6OpfYKDEmLNGBsAVcd/K93b1cPpNQi+
DBQ4sv0c2Fx/N4tpd80TCVx7IZmpn/N3K6iAD2HkeMMCxH+T2dWdFo6kbcKWfXFKzeap+miMFuU+
ee+dqpbk+kDlS99wib7g0nDNIfwMoMk1Q8eXr4fbByWmc/PdotXO11g/evFM5Vi8Nfxr397iXyC3
Cmzyn18kOxTSvhEPMsskxRwUVhcCIzVLdyJERNzljvJS2VoMjg0RxeKiU7Z+jmjntOW55vog272y
4qkN5zKsqcSzqpzpwcEGe1MVKfL5RIeUwOZ/QOBpEREcK2Vh4yT+F/CUCfVT/aetQUFpcI+WkOO8
huCgueiqKCPUvl0cwzZYI9yIUt2u1MTYCXa+UA8LCKDjDVtkG9XXI89TXrg0xDRWSllELrXxk7h+
ccv9ezvV6GBTbSa/UKF2TIsfJLScanhQWC246Cj7pioY2lsmS+HvT2yGBfkj4a8svXSPBynF23yO
h4etXB0RqmU8BbIWTe/kd+rXmLt0y1t52m0xebgKXSHFqX+sEKm018V2C74+HegDGZZIr+VIDvlo
DxGpg6w8swNlAX5azbbGx6pVv1uFtUkLDPpN28TIee7m3dJyhzf1sqBg+PmGEaw3mdht0/zYPsY7
3aSFoxtgqoNyMpjQw05V8/xCWyQI7gzElwB/t2rvQbDHNVAzgSFBqGaknuYYmAshnFWfy0UjggkY
Xqa1ca9W+NJui49rYggy9QPaTe8umj6Kg5IwXQs0yTyOMmDFdAl0QzXmGtqckcl8Ygg9LRPx2hiI
mcny957q5/vEmPquwXXemdrM9TdDPEddb73gE0YX2R+WrTfuFINI4kSCPKsn6C0rZA+xYdwnQqNP
7iKLwudNLHqXFmZSXVcFrRDBlBE/cQSL/D4OqBvfmxYWAXo/7kq26gZK1s0V5VDViEablmukkufw
fA63fPA7gC8zQTtKq20wWp0wjeKs4U3hKENnPAN1sEfspyWgy4M6G4lWrwfol7o/Y95MmxNxpbL0
Dxq+EXWTy6bct6c2vt/hdgWRc3M1lss//AgpjYBu82tv7ZrHSLRSiuoLnQivDZFyvyPi2YD/cJRh
ROVzZZkb2Dfjj/sfZnsJdV/445t5SuniXCGb2IL8VDPms92ECJAFUmGz0Qt9PklOxq5cAwtVS2Jx
M5xzoon0cD0TVpD5w2d6QD0+X4Gnk5N399Jv7+tHPqbtXHhxgxLAZgWQKF2bbkR62R/fyOB1wPDS
5x/IGdnQ0e2u80IhCelXVqzAz4bf9BHr9B5FH9nqBJJfFIkVLITsDyiUvGHbicad509VM6qtHBvT
W5hPYt7JWRpQYdkyMKkrQ4Be0xgnZjgEsgvgOyYGOxcyx8XUyolqBZQyhLBn5vTeV276mAthgaKL
S2S0j7R9+TLKw8hCvmNEUAxxQvqKHDdWQW1PQIns2w3+ObszB6yurtMODVGBzFrH1BleTdM+GBt0
7uji9nyK7ydvHpFytfgxc2yjjz0zXyJHfCMl5FiyfbMT4qM9KZOdx57a8JJy2HbcjDfQbHmodEEX
r6OvLMmHwpjqxvWrYxsfkockGXAR0rwEw96A1aLFGJHyXpOMlP0KOkCiHONpHHaYs9JZzkm5Wz6C
jbhb+CL0uqjqT++Cv53EbNktRh9y/yerzRIBkrBVHmu46PViuHRa8Hx69NMBhwPUjBgSLRcpuoUg
Md6911em378MLZnWrSmor+wlrS9OawoAcakXFJw77u8SfuJWFUUimz581BZy/G01dr9iat0HTEH8
MZZ1LMQxL9eO8lK3iENnOhD2uwL9ImbRTvUXb6AHDx0gS0gvhRQGx2D5Mh6B2Kth8n8epFbsimKV
NOjPvT/WdOE224woeycouC+zjp36/jX7jUQh0xLap/SGSyhKu1xsjtKEftQggIqWi7FHNJFWhy9p
wOaid+47EoPuR9fftXpZkJd7aY8u1+nmAYhdGfhTtcF6XNRnNSZHHGABrq0wyeXL6bJpqF8dSGa9
loJmRaBFrfuHUt4w+sNuVkNXATQ32YonCn8cjp3iR9PN/ke8vglMhLSVBthR6pePI3cKWaiQneHn
FCUcoApfih28CzVzVihjXkKV4M1mFyo9hCVrzgQGODwle30YAZbnQcg7kIfxOBgUjrnv0Z/OSZgR
LQU+dVATyU1yEA92rKUGr/hiMFdA1GuyaUX/fOEqZFGTMs7WPPMDlw+y8ZZDinH0WrF6IfMYNql+
ZgFbycDezKSFqt7ijpTJGY4x7cB5rT+a9x9KiPpBwnQ5I2Ty71uStRGX1yKwrWdFaOglZ24XNT2b
pMPHE3gmRGlLjuACrJvfQXKsIhuQzYnkUscZNHzVags27wQ11pgeFJrlpiLe31GG66tcjwpxTuye
3RTe5otiC6LpTJvw43Yy2Fqg79O2PqeKRKsmLLEs7KigSuicGYYbJPvf2b2dtraIgn1/1eKp24XX
dniWV0MeKLogVS+BZd6lUEBRTjhpuLUKpMlpWmeJWsakSb9FOgY+PN6h+5tG82maPtR7jV88CeXP
Bfkv6rapIRMBubwWzXIh+qqVdWKFVxfdsEVkqfclYiJ4C9oi7yhVLvphR82YV1GivFeAfzec4Byx
VIPXi8utdCK4rkXee6zU9VPuNPTRVe0Jrin7nvRajbNNylPnlYZg4QLym7aF5N/RyAN9bHHQOz3+
ok4iJX/gDUugMOt92e6Ll9SYes2KNB2nHyYBh0R6pPQxYrBpUO7AZ96cVosc57cs5WYVk3zjSrhZ
xp4TsacrB+0ZY5gnpgYGeCqZ+L0Bj/7tpnUoyyihio10nE1Q+xzsbpb1slrttInAhSvlR/fDO4v2
gskt9Cg7+hwfdGevRdq87cglv5bIvOO1EGNV/cujfAnSlFUgs+raj8mmlTwkdD+v/S/8DxNCMalj
C5VcxkH24T/GG4uOOZ3Vsn7Tlng8ybogQO7SG1mCFAlLqrG5qPo6zQbq4kcp/eeAwxK5Ip0fHk7o
HqS17k+1Rh032hutmi0N2yR+byRcRkWo9MIRpK3OgJHVcJWsy+DCnAxnLucScL4n2t3XSfVTDk/X
ALH3MxqNzIQXG1kQ45HJff+FUtRMHYcbqGvXdsW+LS99/HhLWhun4ikfojeUx6wTJgU8DslIeV/k
zM4RV/tLMn+xg5OEgVCzQaohGuX0EZ5AkdddbwACAT8gc/51IFBUJUdamoOh6d0agAGEA3tFxDCH
aPFu8bbkq0bWBJ2mWlgH1fZsllpfQxh8WPhrcN2a0WwabFdbINsysU8TVG194mrJZOnyQjNT9yc9
/rwTz5MpV181O2hz9y6p3n5j8oVFZD3dSMjP+qFsP8T0lU43mJEXaFcoPZre3YzB8dTVOMx5pBCe
+3OcEYgeg5J6EkgvqIF2ATcRS095UolLpKcufx31vK6LIgisqF1BHEdzDwJRPlcodlMp/xZiHvgi
7exV5Y2BRySpSmUlRqRSbuzin5jFaRCS/faZOqTSR/fDLkgf+8BINsQWyZPpT3jAAJw5S8Wi9F1p
yBG8khnSm2dPBBSCXgi7DBxvBJ6rAT/mH4HemF3zdcigMtIrKu0HIGQOV2DJsg5oWy7aO0fc/BJo
AjgMvTLLJT01qiu4dp/n8TAPfN4WnFUaaXEDbNqi4Nc/PQsKkhHFc2/LdskD7vC/SN0v5877TnMX
87yAy/aMtnpVn5ojKSMgAa3dp2w9+PH8i6zXRnAs90zo3yRTqYvBoGWb8mgeFlAZyixy72wvnX4Q
n3Ij4mu6PoGyR0X6pazxN6zdY/UY/6Ikts4djpmqe9IfTam3Qrz7+mxT8X31NKABlcCC2YRdu1M8
ToSZdQ7F6VyILWs0XxLDVbu9bYdA4IRXti04w3NVpHjUlhD64POFRDOjLa6XV+RBJt2jiZC1uHyT
6vfxvFTrQuhhXzknvVTGR3KVCQwvULepBkvjoWJ5d0ReNRV+CvaBpAM34TnIWNrOxqiQ2WHtKGoM
m3s8Psr4o1m8IZKJk3EoZcTppdeASlPYATatvDx3JeYikbcmTiJsik/2qq4Vk1Hr4T9UMSjZ94vT
xSt3Ct0LA2xggKzaZM9n9Zn0+LloihZ3+DK0uydN1g9toYtty677FyCX0A5qBEl1sioc+L//vQxQ
/jw6cDgZwqoLawomb/Lm8Lh9ayFej9SGyw/ArcuY1suI9KNcv7ntHyKPg5O6FyluQjo8CObsfZYw
DxKDNBKbCjrDZozEjvOSNknD1hKqm6jKKJtDjgWae2TH/917QoZHWBd5faqjjJ+fjWRo+8lVzCDG
04poOGab4Yq7GXnZ23XoHc3PMovp3nT9BL6qLcFVwkzM8JWGtcq6OOJQfizBa6fsKndsigMq/ZaD
dA2XlQxyXQ7g0/Ac65/+SAJbr8HLbjNEZifu/gbEt9dilXfVr0IrbOpCp9h2Nq1THo4eqCBaEGGH
+PUS6+rLo1jBv8LnaE0YPEoY2gf11gJv27DtxEcA6u2NfLAtsJdBn8vKRML1PhjreIIHM39Hf0nk
HuVzOg1yKNqOAARyDcOyrJA40ZYq3MxTTt0f51xK4l41ujlHhXFBneKYV431Nlx07TJU9LwTAz1W
OQGZ28U39xZzuPAPbzpra95Mw12nNq90Sy7F1kPyTOqHxLRT6Lpnt84C63IZz6y1zudFRrzCx+pt
b9USkKOHgBys4nkf+ZpKxiYHjUGx47xI+CREmHDzPZ18mXifDXAXoKr14p5bcCtZ7nEpyX5mFCcq
e8XBS8uSS+//JBzJmlZrkuQtgmhwEjXx7Zv6K0V3uToM3AMULlAfMtyxf4FTVv1aiIv18ZgjhZxf
m3Ca3MbxX3dCxytx+Xhi8jlxA5uX2C9Dxdb+YHsqOUNVYav0N+K5M7AF+EVWDpSizA8XfXNcxmgt
3v4WfhfltRe1aL5Ej5OyOlnH6CBm7D47AZVTLCXaaCZJWN/FexapH/AWif4Wz07dKAhJVUYDJkdN
mFMVKIDGU/oGWIUObYdFl0LflFQqQaE1aLct9C+sbz3GTRrPNP0mlhxblrd3JlWgvocFE+quhleE
plC3+nNlIfpz7Zg0LgPdRIZQ6qxYD0zjUzCyFObum1rs6oGfp35Juuc7etup1tLH1AaJgkdw2Wqr
rSeg1yt8ExgDzpD2oshHJ2/JBenRPBx2Xv0oag0E8F6o1g1IsdYE1+KbB+a3F6EzO3r5WYpsVUJ5
HIyU58zKuqYuVCipncmoO40Hw7HieCHArLFmuk8JxEAlh2z2dmeVM4i3zmkPZCwFO8ZI/y3NfMC/
Hg4A7O+tALQzDrOsHSCkEisGdjjZ83U9r32D/S2Tr2nAMkfy3K9n4oemUTAn/njWLms3UTyH8cDo
9BUDvO3i2S82AZ9Co/r5MQWU7nXKESU9v+c1VWHEXtCOPE1UaGjoBOLt16XBp/gRfmKYZmIT2R+/
44jVSKpKrcHw+Y50pOGLqU+4x49HmyXJifE/TuaNi2vrY4qrGu5v5nfVDcmIR8nyMBMFAfQ8j2MW
67GyBFmqlh8pkZ8MclTtwMzD8Tnl3imo542nMMaEliOABCinjvc+72CXuhLpQ87EVgk5oANTF4AM
8st6U1bE1kEnHiCORiE/2B2O4iaMr6OxDAloYEcCnktgLR2ckp63mQQHX9+qbM0AS8ChZ9rCKa2F
bsWU5lr/eg72SA6jh34dH1x8UWr+widjOjDqKfJfjB9r8THmzazeibr4/CEcozQ6DX2aEhAZ3Mxa
ZcihI7ucPwQaJcdz5phV6Aq6myMDpd3xGctb4exK/9bx4IWwBzGsEiSS2ZzXG84Xw1F3N8SnQD3G
W0OMIoIoax8r/twt+SqpxUoR4KyXTmslFrLr7hXRPOu4wHymmh+2dVvQ+gbcXUv5do2tdIqrELA8
6zCBudiNPiKSsG58XZUXWzK3P1MELW/xGPz4w7FyiVO9bEDGleDdHZA+Qoa0wpx9YM+aGBtEsYzT
9m40i/5FjGhZyVJwAAj2Cl824j1eBcmx+1CYYIgz7a/eTQFV0iDktVOROVnhdpdtkTDGac9dt//J
5WN56GWcjypAMBPWkVpg2XcPb1sXGz4Fyy5fwLTQ686LxKRPOCa7veayVDbvyDjAckHrRwJc1jgi
smpH529hodGBPg6zcONOuMtwQPQZasiz9hwYaoy415+XElIEx771E0QEbuEGKah5SuLYRhxlOv+H
o1/BL+itCWnCXQ/NI12jh9Grn7sul3XFXrb6b+zdlXgtJBEmIgXI16uMllmfAOR+Untdzf2f4dMD
dbcIKaJJorUUAxOGAmsE7uh3nKuwvlzJwVCPursaEap1nynXqJFXH96vFyc7g5HyR7c+UCEvG+Nk
erST8J3ymRbypuqSJ8Rip2I1OytKT09fJD2kvcpZoa0r90+hhK7OgotGqY2tfiGfSj12n1cYliBD
IzWoA87+/a8Ps6ebBPNKK435lA4pvQypH7ZwgkFeVlkHo5by6fXwe6tBwYZQ/2dU6BA/dOjsFjJC
uUFiRUkqD74o7YmwQVyQUUYbzr3PF/jn7FGVbN8sKu12grgVD7baIDTo/5T9mkzdIExKNWkak8oh
SUWjO3Hu8o+4aRQiLWrkPtxnLzptiZ58OvjXMO0BNxtGuWPqORa9OmLYviIzeYVUwFrlyzNA6a30
sc6382nERs6dF+9Pw+jgx1qcRoy4ifBKbmSH//GtSNFRlgIKi1pg8cMEOmottIyJ0DoxCEBY0n4r
oq5iiaFw5IVPZqA/t86Clqi82dB6WEDZYpu6A299k8IYGDoi1gs9tKNROW6S7BdyaA17DDsaIcQw
0yeK7mN5UHM7KOlcFoUvli3Mf0ooBw7PSoAquAiR70gpO2+Isl/xJEm6xEMoAZZh2uTdw/CMFnnm
LbU7L2/xqPz8rYSRU+dP9cMkl/Mb7rJr1F93Xb6thXzHT7V2jz8KxcdCJ9M5HWG6FOMtFPxwWgZg
uB/kaLPDoVjLNjkmXXgNAIxMTfvvk69rlx1SRHk5b30aTNPCQPgZzDSXgWuYM5TEmydqLSB+BM7w
nfNuQ/b01hJ9r1r9x0z8KUDfNOyGeju+EqJoOrloNd3aHtYTNPMmI1YrLN7tv4gtHPnXUtq6oGTR
qHDgS16ydq1C4Gp3u1pOYrlgs7ZBkg2jGIyq94vTy4i6SYwpNGL+TQR3XPbOwjpjUEksXLdfudZ8
tebxo8WpYh5Ybm5WKeL67zp3I0Cy/jLb16AtedVKzTO+J66/kgnHP7f2nHY1NoOeg0D5VeFVVAFQ
6ahu879h7XeyBtat63MFRF1cQW4WsCrfLW08IHzJZ+YWOo1G0whMBTL7yeXjkjYAOwwgtevVqs23
1xbOk4R0u+UZGTaXVzjsXMpSm0yy2PLNF2dmqEdfJiI3XAD2ky1sb0JrYL7fMJa2E7s3nSfpD35n
NVhdrtX+h6ETl2iorg9ut3QORIBmCMEC3d6nqaKq4os3W6x1zGfuPiH2vEmvMJCGxycpq5a3zy4F
2dWBN6/8fiJi3u9fiYP4C2KeygL1LIAL07wbUTcmJc3y6LYtTHOSH4o4Led23kO8gAJipme903lS
Cfiaf+IZLBY8f2F0lrTyK7uea71+7sbCW3kEg7Up+cLTlPb1A9f2+H9gOj/7fq/RIu1p2J3TAjBx
a0cWUteYiSUNBfCV9EjXzzXjjrkiPV+abKo7tdHREg9e6aUwt749zchlUuvXWGQI/DYdFYycEIWb
rYfZSozOy9r7LtpHbss7PA62jG1S7zQ6NwLLaFqxJsrstfAz7BIIjjLilE6HyxdlNRdj5TNlDFSd
4W1jOhhkMEcLDX46Vje0ePShp4zDOUEZAAGoufdfBGDutccZOyRXxAuLkp2+5B0KOo7btTWmImRX
xSrUZNxr5Kz6odDxUg8jH/JQMEjchWnN12pfMAuLST2lxOYhGJcSQ3rtYiSFOMV+noYB4K2CbZm3
8rBfGLDyz3RvfMXZ18Me0itru83oltkG6T5FIP7E+DYtZnMFa1PHdoPfvgaKcEAMaHCTpdRlaNNV
OqKcOrouaU+UNWDjj5DcLxu32v9LA+LLVywnZ5OEUU2K1T8rsu1alKZY4R0PJq5umA14TqiAaq0X
GIRQspbH1bO0uxU/9yJ3bGKF+frn2flEIQnyLiZey7jZe/rlvriuvwIcBNor/k25XA2DloG0ErTt
e719r9PqHQ98p7kdv4wgIGboVbMEUxubdq7HHOh0PgQZzUs0kR7q+K2E+ZBDCe12Gg5k6G6v4bE5
AiqDUWOizbN6pDXJg30Kyd9Yr1QKncjx0pq6Z8FHL9crh6zmeE8nEhrKEMMUEKV6+FlUhLs7sO0a
Ulado8vbaPQkVwqHt/el1Ovg9heA8XnA+t5OU4XYu4YLIzwC2/faChH0bEyG/QjDAdwiAB0iSUns
OKkjeGGnf1N+q4VtwWJVcfSET191Vs79POreeEmtSZN4ZGjjubVbUL4WIYbmg5zR5PC8DdXVTGA4
MQ26gh1uSCNKU3tcFdEmV4eMXJXzpBpPzyt/MgS3QC5VaCoxWRwnKvf/UpTnOED0RJ3sJJvcH1hh
vQDJ9pFFXD4S48TNPiux8w0o0ebRMdv0qIvfsR3RqGF/rlqxMXvci19kvhKO3qt6FcKXt0C+4oZB
K3JjLE66Dva6Go2wq+eqe6+wZNwfrvS4AkZuFVwwq8UM+4hGzr8AQyuU4KoIq/E5SUy+YF8EBNB3
ojXT6aBwb0XEkNtBXV0Rzo+KsPG/XATGkc95vKNfVYMlEFDStblYZ/EeNbkk/enjj4El7olPGl2d
GQZ1iemP8kz/iW5vHI6VuX0VNccCC8HRsA/CpHbpGuf6u08J+0ML3XlZpPaQdevLFY6J8ojH+74X
icj2BjSuChxO0VA/CVJRdm1tkfwG9yMCwE2e7F9p7RwGZY1wUt17dtVx2q5NE3yNNzeE3ARQt4KO
FckokrnXTRdx/UkvnWlHs0ru2zm+HPVfl0BFZt1z8AfX3g+mKYhGfEReD0GQl80VWJ88QHWKHV6V
9vJY1JDtW/fwoxRXZU942og8eV8HiFCNHEpua5Ymc0U9lingnnBubk64i2EkNtaIlRzCyKtwINz0
nJgN1CEcNctIQcmULq4IO4ndWuCSrHDIsHWvouSC9RH7TDgBKNule13RdbRyTNh1nEnjE7CSY7Kd
pTuCBS4m5mRbANqC0L5/t9ZZp7rOqihm/zUV7GpagUvfC5eJ2r3XJDQXOK3mPfxeRCP0bXLApHMY
sm6JXjB52kGw/vINm+SJesj20hej3AGpATqMdZjFkmaCc1uXY+CX+6oZT5i/zFcSRf4YEQ5QMNGk
7qaVMPvGdQGWJIcyggKqc00eeMOiZMC9t44CEsGK0yiB07akmDpIToVmO02OSj6KLHkJouXPY3Lq
uANbVoUPHTnIMfbXS0hRDUUQLb1jKjbaQ1tou4z5dsjC20DkH4HU7r/RTCi6bfxkZzquL6xJW/d8
9EZZXqeU6DDhyQR//0DoruecukazKGpnE/vApXlragvFamZt+7wmBLTEL6CqUNxNOSVLOeaTneMh
2+WqsYuqpwnZYYv7aB6cli7oOkxtb1xUzaO56H4C+7RCFHHvh9irbQUpv+gGUAkM4UxRqXY9xenl
kEfFgcCHX9kyVslwywc31pXBbQEuGAGoT3kFBu0BZAK/8zYxOvks3TqLssHrdmeupzG/M4SyROTp
cvhsxZedqI4H5co003hL3n/7IoTXMyS5zeNxtnKqWsDat7ErKjbRCwqj5uj/U5al0FcK87hbqn2q
vH+8IEwXF+8mf/sGg/C0jtKyHt132ADK6JTAwSr8OM+bV/2OULlP2RX8O5iU0mv3mVy/v+mZ3BaX
royTWB2klNg9ex4fPK8HhhRvrw+nqYFFExYx8f0L8fZRdWhKjDAe8gS6MP08gfNpnhKQdRYH6Nwv
YVeu2dBS1zmwTvJ01E4DCeSqEVLlYShdxjdIZhugtWVl3Q8ji8XClgq0vvVnhzeSzBpEuW45qZ8P
K4riaMGsM+J0O9kBkyyNvDEwfE9ApLYZUABpE7ol4i6xTagF9QWVbTn6KKf3UysOkBCbLZ6CN4t2
O+66FnLJWP4JuZBCFpoLf976WW5p6XPbhKK4q4AYEpRqxnNVAqdTqpIiRJWVz2tA9JxowM+gu1eh
uIzyancSrcrDVOcPmPKVHsAF0tp0+rHxLlkiJ9MwPZPzoib/sp724qXF2gQol+Q1OdtQLwrn5acX
VSbgxMQf1NLpLnprSj9BSV5Ldz8xjYF45pD8FZUsaOru34g0BucBjc++e3f9YP+K9iUXkLqP/hre
2jv9qly6gQ38xuM5qWmLE3xp9kJShb0uouspjb2Mhdnc7YOs6cPG7Uty9T/9CkGk1QGLKx5M/NTz
EpFDKx3pWplqJpZf4L0Fx3A3hpbqT23ATD+IxWUP4SJ8woj87x/O5M8RV6y2rpKelQSxFPCRi9Xs
aUFlzK2xiWlKqso2HMq28OkgenFDu7wLl2MFKG/p4r4rwzZ5+ZL/FweLdHUKoIzDvSxrRSdXAOjV
tiG6hCEDOFODKrgvg5/QyLwV2m4w9pg9jCy07rd3U3H5rB6IkrP2IOsIGmFB1bCcRw61b+mRh53D
uCdL8z3OuxLI1TP6Kw0/HnTjQb8usgYfo+XMQdCmYXMg4TSY7KTDCEa7bcsrq251y5Qq5V2TrQQv
fIkDZRTqU80oInocgM0wh6TmFG0DE9HfqEIS/7D1RJ8OuOS2/1wlFB3+Mfi0pwraCteeNTJUJxUh
hF9L7j8yoxHK4cjpfIQGlBNjA5+LEpRvIQpZK/SACqp3ElWQKM7OHPCo+MpYX/I+zVuOC7dzaMWQ
iBrFthFnYttab1/fW63cfZqpB4XRLRtcmVNf1siQ/AIkg3bp3iuZy64XrGp0R5UOiSNglFzXpIUM
lQZ1sOu2XTf0LhUqff2DO8XwVZg5M1kbAH4iHkCB2OACiRmSpGKy25CR+vrs51RApkhVBkdBe50f
feO/FIzGNtDu6IazzZWyYH8u0bB4a4D+FsRYtvUeGqQKTo1bGG/x5S6fW+RiCMR8k5mtxvt/eb/x
aTygn0w0ZcbhbPPgvd1lyLqNtMSVAsW5CH68/Hh48sZAQGJu30iP3YiYYGJWNUBH3nDocJfeMzPk
/mlsL779nE3wGl3NS0NPDpMWKs+SSXqy/ZZvFa9AMEHKoD4+0PZByRSp1EMoIM8GlR5Tl6192lgF
gxjMLhgbysMIPW8uE42kpcp8yf6MCR32R7dr4YPYxzJeYnEoLvhOD5adQXtWWHZyjLBUe9e05Jwb
bzQGtCl+gDqrvtNRD3MBDbaiCGnZ7uB+MRz5T9jjhd/550Sv/02fh5p4PM6ovRB3LT29cSJA6Yfr
uyBbDQ8sBrpi8+Ch+a3sPu2xzy+RlCUcBZqU0qtyK5mWxVwy4BMdD2zhdGD5sIOxCsodVDe3aGS0
sD5NmvpLF8bmD4COCcRaMzaluYvsEa6OsyjmVxjtLpETxMVrL2YUvGyx+SuCzUPEwir8yavBBh6X
xpDSjmpqXUJHq9U5/DdaAAxAR7vnl5eFbhPz/YmUU3wVpXJwAOQgYK/cvsMXJ9dAB5SZTOWcK/Oq
et1K3eIR7M5KM/lRKgQNHXm3gUDuJtYgWHhawWtPBtfubq23dB2rkufvdGEldqW34rD+7Ouo64cR
xD7J+H+FtdTFUx2BnAFAqFc/nRceIWVjIOei5hERxsclchs/nfbqnAt2eEsIV1Kv9KlGKRV6ChPh
4YG4aW9nQhDoMnemkB41bD9xHeqJZlsjq2eQG05wNpvHeFZNOP55gi9aTGdq7U7C3MbLO6JRpDJR
+zY5w79/xCGjBFrWuGD8iQ7dZUcKj2bXRCh5Lu1prmQuJ1ns6b6+SMWZgOUX/+/dP2q0u8s1f4Dc
PHE2Bg+Fl8vopA3DURN7ckHlwwp6LlCK7m2JrlO2xzUbDcf44TUpGrgrYGIOTM58Dk62k3/6uLnc
iV40MyxhwyKY7wTtsS8lD24QXYEZ4EJ9ptCEWXdaRx9n717l85KqxepnJDurp0qoxHBtr/tku8Gj
JfcG6eluHvTChHP3SdF2Y0C0YZVya8ha25xS1w1VujGf5GszIVpn63ZzFYbS+9aToj/5ucFuuFf7
EnpXaEbgMOcHN6sGvPzN/SHMPmR9l1ZtAQtjDx/6+yoMQdmZxEglENxYgU9LLpF6oo+RSah5uofE
4ZNONwOELfH2pdVcOaRuNipDgr4CE1MePAyg6Ei16XAeZtgJFU0X1ebG+eA2Or/yKDZcxD74CHlG
oCai0eOaXnr0HLDL5ogFqclt23WVTHN4TvPI1J5hE5Yydd7S0vek9Q0iPuqdiExTULKMmjPGpcNn
pDKsSpaiFB1gn81k875ojcWAEgeW/wqJhm0DwO+LByPGOzv+ruajEWOfsVGuKcOuB7cVtVrqrg7m
E//UHuoZanAs0N5OZgGB5LSBf8ZkouyJ9FqZz4iTbk4XB15vreB6DhMZ54/MphD3NnSKHxN7/WF6
e6ORI/cjVpvtjhhIgzC2xSRXmacnOwOpONpUUp30vr/Mm+U8lDkwenbfqhnmaRdzRSzJ17Nt8yzT
bHfk+gJE4gIKNT+MWXFRJJw+JE0R4V6JuRUPUUmGVJWBV0yiQ22Q9RbVdkG3p/o3BRho+OvPEYSH
6IkvAknbff8ckX6YU1AeAQPqgV77JVhopE37ePNYgkz18rYGIXyfZVQkOezfNo132qD2vq3OeS5W
QNVdNUP+hdaGOAmwjj8HbbOnuR1rKGaFQebkXqgabd1cw+MJ3ikCVMDuAw4K4V5K//Xp2sG6YEkq
fCK6TWjyHKLeiQZoAPfxbcrAdR1PNjZdT2yPeT4T5UqLn0r5l5wXluV/I6jF9VbvU3wvq29d6fe8
TWm3sxK4IlKjQn7gNbKNxYR31HHDW8+W5DJVPj9NYxUjUTX2g383Ie7XM+4XMUIvfObDnO77xaCO
m0q8GOvBAgf56gM4r0uuED7oJl4KT7gCIR6W+7FKrAun6+W+IzMfB7v95VhMVX+rl+YQ3z9iEz50
FIGJVbRZZIG/Czi6fBlscIxe1CYgZAnWV0jdsip7LuUVfaF0sTwIXr+bVTgefxiDcjMz1AN9PwDL
O1z7iw69X+mt5ilARTzYNYgANSfo3Xgw70aClgaiOt2IZEvunqmJ0JvZycCKUSEq4nfwcufmhXOy
0JpvilOv4CGfGUzzilVXEbSSHpr/8Mh5L0l8LY6K1ZmzTHoJeq3LH2UjM4K6C7hAYxo2ruQcxHbw
LH40ECbmjvYsfciREgX83lgqKnPvkMHX5YIgQz2aaCem2B6C81THlTIeSTxbKpMRqNN2t4xyKSV+
75/Z/joAAyqK4LOi/20/FyucaJMG9xWQOw5EDATu7EI6tU1ODICL7zYvneYF823o9CesVoKUgDXA
Z3WunqLBWRY2meYq5TS4g2xeqaupFJdQyPeXxUVU2Ue4vaRHFd3fomZmsUNlzZQ4flnmWHjjR7nG
ENjlEPkAgzsd1y4yApOLEw9YMSV+eOCBfhmwulnc8eTGpNhBLA1MGCWFMBM724u6yvtHmp/F3gsL
Te4EIDc3zAQ6Ykjay3VhdEh5yrLtjwIqCZveixlaVs0lYglYyJAJ9crHded86MxPclLOyl5dklZD
7Um96EebLhqWVkUCKqYOu5CxHr0n+3Xaae8OcrgYjb75GaD0Xo/VrSBx9uxzi6z6NZzpbbA1IkwV
bDXUAmO+80JIgC1jx/AvSXnL8OqHj5gZ/VEVr1B6Bk48oo92PknSE8CigAhWMXXp+XbSV222rzwU
ptDh4qtTAvU1Jc0Yz0qT30n/Cr5KzKanoDaPkfx71YpVopCW/vtjOwJskJ21lb+zpa8f+Bh+2GgU
04PnNk5Nb9SUjobhxZFVEpJk401w7vFQ3I5Sqk1p87OaI5JT4tSvc1Jhl5CifReoJ2xD1CQuzZ7K
zIELMEsEihoAz3wrKhpGwPNjJs/Vw6wukQuXIQ/LS94/HdCkhEJJ4bjDHxejhbiu0IhjesPYY7+Q
JSq8AujvATLmD1jr4+VHsUSsqQNNPZH5NDfh6ZkiSACAnRlpmyMZaJkDxgOgf1oWP93pSGvPXws4
K6QR7MPKEETO8cWCQulVoQGpg3Ssp5jmU9WXAues8SWslUIdhh1dmoIgXCHLTt6jf4wh844qT6Ue
kNUEEdu+zZAY8NUEY6RrHLzpwW/0EB3EswcXJS0BLv+Kvcxxo5lKC2io8GrG2U+811NIL1M5+gH7
RS9+0gAGgova2EY3iQG5JIwfh8OjkN8EAf6tp7gxS5z5gwbyA150JdHLOxHkqKPQEv+61NmaACJF
ePzHrk1XzFytXY5aNF3B/RuM9P7aJ0nvVjARgKrvKibpB1DoP8JhKUk5sVk9dMbitwMp34Gc5Mz8
xuG4ENPWrVxi4ZxpgaLWXq3wVaSF/KSAIZYUtv8X9yiZcVPwonqeKxwfQlA5hMX5Dp2TT72pG8cD
IGuI7u346fVGTDCpvsFF2WGKo/qZE9Bw1QjUuKUzayjbWlkZI11++Blv2dB+hQMPyHQH3bMtOAtV
NQxm7hjtxfYaja9vGtLktLZNstUD5X7Fme/C3NEzqMCL3k0F2lDR7eoMVQ/cgYSUmlJqfYyEegea
miHVOQqhGYWn5EebpPFyvvKTY0jw/38aM4A2Q3lwHZ7LGBuRRbrSp8ohiS5CmnaMAoBAMD6ARwn8
IbBVbgi8Ml4TEk/1b59tq18YW3XPrD8eGbFI4zhmXrnBb7MJtsQXnRYYHh9E4aIVUV94L/LKW2Yf
6VmnDldtwxzfRPXXnn+F+X1Asuioal0kx3kkrGs+br+1SD2E1AUsMUIeRYfcj5sN9KNWWeOsrHXd
rMuT8K8jZpJCtxT40NwHabiyaLhNG3fbe/z+cjoJtnLOi9ODyDszKMqlsxR4340fxRFydx3T6IN2
Y9Jdm3npQAbKB6/wnvxXsYYcxsplGbK9brsXg+LEw1Lb58TS76z4no30gKu14QNUP+iVHTznpKCc
QnmDCzaMmfLfNXGx2GSjGl1I/S9G1ssMMKB3e31Voz3jQnefamI76NC7pEynNDl1KUBwWPaXvWjL
49Sb7ol721ngMluQdmEqa8430BTCxyqJyk2hHhIZk2YSya5OtrHwIqS41nkM0r4ur5PsY35EzqUO
6P1sy3lfW2NJksyrbR48XDtR21M19EJpzDHj8JErz68xmEqpxh9m9/0q719CphTgTpfBioRP16Hy
BXgngGTArmN6hKgwTRPkROi0q5Zl+wTQgF6rSJLGwWAEIWHiWK6zZ5e15gyKlWnZVIN9K+VW4lYu
qg5kTTwUY8+FOPqLm/jsmPk/I7lJQ7N63hBZdIULLN2sqdq/1lw5sdtlp+GMrPvgHw/ZPR496684
xdjVDxtU/lV0IzSyoLsamYrpb0HC9FCSsMqSZjtVJHkFQ6Y9CWxFPDxEL3/djWNaQM4F9Qc+B4QH
gfOALDOBYEINNYhaetsTDiLap0tjSkU0ik7H5NrRS5BSIMOClYeqiBluoiIH44LaJR2yeCRr8aBQ
IE9/N0PyoNpoKSzw/ONpCxDaHuqz0fA8wEpn9TMdaMiumbi8MXrwUXVR6I8izNUoT4qdqnfF+PUy
u6wn2Bjr3tCGasxzOo4/zyHE4jkFf6AALR9T1R5oSg1rOmBP8yjvxAZNne8z8W0C2iI8iRUJuHUB
oVI8h9mDLQBuk/Q8FJ2zcOAyHPtGc5BzRjXOOoSDmmpAshyMXF7K0MsVSHe8tj4jsyJJPZJVNfel
su6e36Tehf/6QgUi9DRCMLbISp5uHWKxymwT7UKGvilfh/m00I++HOWoIISHhaIbjREo/YI+CWsR
fnv1wkinTEOFbytcm4iljTjxASXagqamSHah+NspMoCR8ci8sZH32SiwyvmHvpn87fENHpUklN7v
8H3ZE3UHIYanO5tsbdgwFEks/nZOiT5smbn5tg0zzzPkMmIfTBF9lH90egvKLrfpkntrsK9sQvy0
/6nr8j2mAmrxWgnuRSW0vm25os8IoaH/m36dm8g3p2RNAl6Ya+n/mDPJAuGIpsXgRfZHrLfQVNxy
5EXtqWeI5R2mb6xCyUW8ZgvWwu6e44RQ1dQD5mHU+j5bCtAhYQCNIhNPWUxZXQ3tuO1NFs3/QSNz
9s1EWDqQH59qX+xuFTMuszmzdLmhZfR8NNRJ/ekuyxTAOb+Hh5U52B8yHW+q1w4DjsefnOKvKS09
cdSCBYLqU1/USp5xljekPHQtFjecqHoCnaYT0vn8PBxFq0XKEDI9Ag3nAZez3NSPM/QRhZ47BonI
2qHF5oxkDbwIy5MLxTM7TCzGOiG6XiUZBg1ZN+SinH04HYUL8HPD9a6gDkaO1Y/qIuiCcSJ8Kv6g
JKKuhlHESHasjl9krbTXKWkxHVlpWlI6SoOZD4O/VTv5XmLeVWu3a4ciqIt/NS35eP/43zjeJsJF
lMZhswUeJypDDpeuT3z4JE90bdI7IexiV5XdVphOuJB1R2klWUCEBJw/QkwO69cfpnz3uSc88YdH
wq0gFe2JAO3uGORLyg+gMhXQSMSXAwrBLNELqw81yQ5W10PCpGOz2LoYh28YSzUxWE96UtitNaLX
+kNhiJk3CNSi0SN2NEEl9XVZgTyE+fmcVXK3F80Dr91cPz6IuQ98+vcPEi76w6klWCVROVNyr0QI
PBQ40Jv6HAzUPqxf1x4ERv7H1AG9o6T86IeKDnt5/yoPaBgBQQR3QvwAU9iyOW7savdvORyoJ5DY
nXzUUrZznzfXdfSX1dGe/Aja86Xp4Jue1T/dcHrDYf0vui28SpvquU482SJgSC8CAor68PppKQ3v
tHbQRfgx8DKwAIMNTtHDmGOkRssKh1M0jK457eGlMOVV7692Zk6tMpFbCr0m8Lmuur3s7oXf9FCi
atA0+pzAN6OWu9gN8eAcEu9g9csQrdqSMUh2sq1Z1c/A8Du6HDe/C+8R7bPxH9KtLBn0Fi/VvEse
bttYiMVQ0sHpwL3Fv2uZwWYsbycUrl0bqkT4zCiEnXKE5MGXT3j2dO+0kpN7JWwynkb7XlSshnIS
+RPNPftOBcAjmrgckS7tAho1mPgtJxKAf2TMSK7++PC2nwrRGrKd0k87OAoL39xJT0dt4eVCMRD0
lr2i9Mr20Wm85Mjbkn+i4Vq4DFmInoEnuZtb4PFI1eNdTOFvjxgteY8nL7F3/EHLZbpH3zU5opBk
tVilMJ2jkgFakTAPq27g6g2f+DZq2Ji4jcSCh8Zvaat3eRJE6eK69WNJrcmmkpCnMfKkLAZELuoV
/zSYFIbwhVAGF1+WJ5uSdCrQIcikjBDVsb8hb1hkXul603GDo5sk3B5tyGwMn0hEQ/7Dqte+XGrB
UyPJBxtgEObaxOw2rAUv/9yNRfqR9OOu85IZWBvYTwWeN8iHKnLKaUj/+PY/Rw2NJru1EMJZsdWn
xcSBickyE8GI7oaVEUL1Av+MmQRow0j/C/izpB8jPb2jtvhKkjq5qcA/IYW9hQv++jjIouaEeMvU
XiG5M47IUUFqMixWZ9a8i1xccLr5vGgfI5RiC79CqQNBODFKU5xTmuJwz219k0CkMnvq1CW5CC3H
jg+ctug0lkXcz8Ez1lrSGpGz5Yb5onI5j7wuv5b6fj5rBKLzQDNM2WBiY05PgiFlyEnWBFWjVIn1
rguIUanbVStl3HRrXkL1aKGcjoLnYcJDc981dGkAaFrMt+gbYX4+dTu2Lc6/e7giCtiDjesZZOpz
7uN8luIkrjsiNJccMW4/YQ1vnBgLeFQeLWR/l1hzhv9y7yvl7MXrMrlrhqWWeEHjW7Q1lBSxb1sO
BA+hMLqh23/dFXe4fLemd34OURB2wIPZITJTvglVMy0kQ9hzNwanFR1uQD/fAHfNZ3NG0gxyIUGP
kvG6CG35+28g4hraj+NKVpgYotWHCuhIirrk/UdXnXbHhqN2KBN6jEYo7NCvwekrObURvkM/wV1d
PKHsm46jr5WQvna0c5AgXSZkcBozrP9+mZUZ4LmruHhXwpHrkhkRJxCsmarAt4p523A3oeIpju/o
BqzCUTheeVi12HwqozW8xSQKnZG19639ssCx1U+rLTHOkZ+KUi6DAewt7z07yQ2V9pOXXIEZ9kZK
862Un0Wi6jVI9GZS16KOvNspNaCeIiIjchaGMEpKlDO16KdoBNkR7MpiNHO44k9YWiSotKXfmngD
DWP1Hy+nONTmYBB9Ej4PAzEXv0a2/axVqiA+8jsZm1WPN8m9ARgozWWtv9IUOuZYihq+B4ioBKel
5S1NK7UvZjB++nD8u78lqrRZrox9N5XlXRBAZN91OwS5EGU6TkJRVvpDZ6CF/fNyxS6Ky4VQqxrm
j3LOtUoH/sbiGn50RjNFWbuh3T2kuGGB/5FlTFV/JiuwFs7PL4lQOLgSHy12ctFW6NIBJKvMmW4c
C1KWN6tau4XLmX9owFSHJqn+tj6s+gU4lFg7tyAwRPzWSMp1ESsa5mbKmwsZwIojyFFGoNQB3ygd
nnI13Qjc27o/+/Eqks66PSo/vKUg+mJwiL6x7etwdnRHlkJnFeg7yelT73ER+gjJgwE/OM/gDI/R
lr7wT/Ig29iC5xm8rENZr+rk9tfGcaUvl7FpenXYjajABPPcnd6fGjQPzO89hMNBrbhuZBABeDp0
jAex0bcNoI0qKfPocQ9oZAfiaBJnExfuj8JeCTDt6qK+dk+L1k44RN+IU/vJiPd1cIbF3fPhulKz
wW024QtbRPMokOd94VcfAQaN7ZyS6QpuH2VpFVoyEp62WQunePnzfduU+DJ3p7gqYJXb9VitYnWY
G1MfyQgtjgIpN67IRh1LeNko1JOD+4g80M/y2gTHkevhwHWKbehr8+qqEP8WBZpvPI0OQQrnfrEk
lZi5GiekB5HOCSMYPIqjVNEkCWNCoe+JENQG7HWQaEeO+ZJoDYGjdENpplehdDDh/g9TXu/tZqhC
ryfnjnTJtBl8dfNKyAJqTfwjGbv7/lRD5/jRK3uRQ7vJbt8Req+xpoVVt/v3B2BkfWQylipZhFTt
tVoX4uSIS1HTLPDAip4UNPXYQplSm5dcSyE9mnsAn9AWl31YUQ3JlbQhyekR4uobyEjYDG/k9k9v
8naVapkNY12Ufw2LUqx6aoVbVASM2LsVN3LP4Kfj9cMpKz6JyyK+vc7eSAQe2XqqrUUNDzTpHnEU
lA4gkFrBdWnZ/tM8WQ3S99rX+uaxR14nwihctb49+KgAo2uYWhNA2vAfom3LgpQiHeHFYtsr5wTu
xUqO1mjE1D0WII8HZjkarc1Jlw8sL+MqLWnAW3KCk9J2lf241cGR1eV89/7q/41JKoJOwzJD0Cor
K4u8hXtJ+BTrvLWBUZFrs9AvRgbRH/fnHwTghy3jrJl/XwSx40+3Od36pRAjvflNHfD3VaEUkNo+
+JQ8peOwJ2cpVSI1pNnpn1EpNDUNc4cd0hDyh9kT2VoKyARmRPFlHWwUUrCnsjl+6794klzgrHg7
VkBlsg9LlVO996R2pnHuElilCJPAVZR9A7eVmdArhQ5TsOoe++KawEz2VSd+K6pwszcmJEmRmH6Z
OhLLAn6vR6N1an1g6jSWGnibwR+3ratdWTgoLccw8br79dEsPe55N6vMZqezrud2lrjTVvLP3AdU
vQ9C0Hl6aDZOC0mKT8nvwjWQ0vfO1Dcdx2nYJRtDM1NR+97x5HkArHwHDSAT8SHY7Ybtl8G2Adm2
z/Fqq641yG1aAoDwR/rs5XgJCOTkBfqA8ThQ0MQ6Pd8l6WOG+OPSo1bUce4oArsx62S4aUuErhzK
rYGTGdEdfGjm9axNungEIR9B5Xa7zYeQLHOj4lI9PMZmIkTFSSjS1mV6vskgtzEZks2oG5BxpTE0
fUNg4IfV5ZY1+x8K9w6KeT+oGh4gbBC0ODtA4tqKZUQlM3k6RPpWBZp2QeqpDV5O5HnzCp3CaiHZ
RPHbp0aHcKXrF21fTC8NHkEJ8EAdaTVIi78p1+++fA1JpXUes0j+hjGo2mbGMHCMkvbcfDCb24yO
oSEeIa2oGfz97knJ7Vv2RfM5H7al4y2ksoAgxsXqJCnuxbyRWqqE0grRdYAWirs6+KJhg5t5o6ax
avygnBKSyVWLAW1xVqKppk5RivPI+q6UvIWC59jkwci4Z2Jev+Wtz/kTgnl89Om+yC0oFGBa+ECT
cUZJj3Nkrd/CXb6gQG3Sq1omR50rOKoJSuIintXtJCPfCj/9h7UdhGxX9/ZrX51EHkxMI9SBWXnC
kVH2zuuo7Gtvv/gwDOuiTsPq15SxqTNBxilovtdsKKbub1KkX5VcBz+ZYvmQw+aE4NVPkuY4MHv0
FLZ+LfPyTw0DbLZ61LPtgf96t6N0+bgYXbxUJdz/TlrJqO2F2IlLwKCfTpoYrQlm0xEQCMOBFa6V
bY5yqKBSf/5jpeVhZ+sI0TGejSdRRTihgp6o1TUMc5n1HecOdfFVqOxVYtYQyoRaQqxOz532SMZz
IguxU3i3dhBw6uz3rmDNX+Xh090UhmfEzBonyPe0MUVnP/yr2xNFhAIqYQvdoN7Eww9WcLxn3ZYL
OeAveZnmuBG/39KMumBPkaNXMMXOloNay8QQ3C+K21OuJJh8BujAHcFOFAXO/DuxxU8pZUzznN+t
3bUBX7U59r0L40QyGDjpEfMAbwaPfSzGT3wOCJvpD/RU0iMv2XlxRkNjuIOr/+CCjq8EspprBB2A
/hjpAFBkd5nIa03cx7ofq0E9aFphqoIXBJk6o20MOS29TDxIMruYvX+KoAcCvCRUvom2i4CCtrQY
geNPFCncGwUc5O5mG9tEaO8RcSslz8oHDUCofP/pAkwMkDAOUm0/PsWegggtt8PiIbfINEpqdPHc
bTvpe5FYU07/2yfb41Igy4Nvob43SKr1TkNM7e7WC0ikJ/ke4fyDruv10iZsVCTnxn70m08s2gPB
OIfui8wtbq8x9C2hhzQUDW0jXNPz/2/87u/WNX2G+jIN7yHhQCudU9fp7PhTwZUTBxas3b2SP/4B
kRnvv9GqCUvxbjZZbNcdv7TSfNhbLJvI1ldghPBvhkWfYEVyMEzqx+Q/pwmwcedsOLHXGy8gHG4I
GsGREAngZDvrzl3XFRcDACGTtDSkhADsHLENsnRplbOMmPBaH6A2PL1zAmdqjums4Zww29/U09+H
8gTB/8VPtjPE5IuNpR321YZ9sSXXUvDMRrgjczRyJkN6/50C58Qscotr48/90QeyRAey2xXwgO65
uBW2zpBGPN0ifPcFoGJSiaOGRHU7QhJHH4D/z3cTdmtz6UxfrUwd5DXR1WqEJThgaMtQHxEFEKLd
/MV3bRdcU7hTOj3uJ+/PnE4vyvjbsy3h5JnmzC4XUgvfzQcsyYX5d/i6x9j6cTQEqO28VhOhMQEe
l2HmR/OfOC5Tk4prgQ58kKCaL5YGBBy+yGc5F1GM7bSIlLgbDYJATxuD3APQXSMrgsj37n8McUeY
lEfWkxhkqgDB97yR/+ecc2Q5p4f1D5R5Me00Dqfaccfs/fxrupDw4XjHrE/RUG5mUM2rcChLr5S+
+FD4OJWMr9U8hdoZ5RJwyUE7PCHiq7JTSNpD4GByrgPXogOhwEBOCcrlrzi8MzgKaZH9qN4LiG3h
k3rKAjYSuw5EtZGkOFudNZXasQWYCYyA9R4l3MMFXtUj+xIscaOhJnkTJzNJIhQAqBb/MKKzuAXG
xXS+2HCFouD1wOG/uUCG3Ek8/5zEaQRT6cckE5UxrPqNI+4Jjzs6F970IUPpqSfreumNjNAx+FeL
OR8nkYezKNckpiJknHQ5LeFhOtXP9AqHsvGFv0arQs91+7kANNOqZf+u5SoSU0qsQhRCHJDqYXdM
IOpDksLXQm+uq+1rR+SPpEDgr7If7/p+qsq1YeJidbBTAE7dUBIRdET4AnSAy6cqf5w9iXXZwkR+
n1BMDeI3bAdTP5DbCwE5THSH8fCFLOjtZbNv6oIFtCzYdxTP+pfu+OgA3kaTA4jV1w30PqFpYSCA
MuFqLeVh497s5grCZVMdXTxU6GjNEC9weauCBF/y4oSmobkXt6ECEeyQpwc5jbtXlsppzHkaEbhC
ZfASXMLkVimnAVqCtSpY+GDxUUZ+VvXWh3Au96FRE+Mnc3pnqOb/Kpy7VrhivXIA1AgYON3NlRoA
c7DUFJ7dcUtWYrsKfsC/YivMS+SHO846aOytBttmWkZ7DVMLH9tX8u///u7NQ9MeR0eyZHtBQbwj
zXbwD91xhn8O4bHQPQCE5/Z8bMPmIYQvu1BiH33wX8lll8JMTQlO1buY31/JzIg4YHPdLSmvreNb
VQIRjlnpt5m8bhD/cAq904qGmDzHcTtzHhWNhcooIci6dxS2LRGrE2dfncqZnmzpk/haMC6CzsoX
lWynjHbIeaNKqUrl5UooZzoqUcWMLInd3F8ryJPU3Ci2N7SNZ0Cg0229sJFUIK/B8iUQaOh3xXDu
bAmC3VHiokgI8jLdiQBdreJ8k7vJaLaCyIRAEIQS3PdijvnFho8YypASIHz6UlFCpOoqcnGUDmu3
g0uJkg6iXheDGRWAnP+gnw0bInfDQIMERe2XX/nP1KH0v/Sr67fSvsGnSmprLpRcokFJB0vyFc8m
vuivBzH9lKuT+1Ltht8V+ZoI3pv9qjH6s8T/4jYivhSTpiC2AGD5tohLQ+0lr4Cb2Bck+smYI9gu
R/zYwMSNzis2sVKi5NIhiLdQBNlQkX2jp/4Ue9RamZsenNHUr7PwkpZYJYsme2t0cgLYaGZbFLV+
a7UeGy0poahCVr5vqLTor9DoGyxBCETTr66Y7iNi4uZQ4l7KycTkhIfDE6IQ2wC7j1ttZL9CuFUN
6VBOAiwI4Rk4oTHtujJ04er/+E9EA8IYEam/ZxkiVZ5rNSOi2Q11s+9Y3ZSUDQc8CjBy9Edpps7s
huijeixtgSSwxXnEdB4LkbB7RyYzB8NJcAlhiISn5/Qmj37kB8+KvIJDI7THAa/jDfMEN7BX8xq2
+nE9OV2KMJ+ioOnM/9S6Yrjk5Hncmf95xWdLZfgh9qBtZmvOA3JlHT734o3qB6Z/cas61hI6/eVh
6HP0btG5JKkbF6TvT/YhH6A2h1Ud4EJ8AsSMF+RVhNB3Gl10Ghz5X6/VQMLHcqAMup2NskamR03l
xpBfZZKzSFrqyPt/SNJqY7y80Z7typjJVWrswVh63a5Zu7LtAScS84iLEKYYTaBSLQGOtFYUC70W
9QJ9fyxgXkg6L+yav2zhqRIPepSrswT6gxPcKFdQVJAPLotDVcEIWNC05A0rXJiHw1VUGvDMY9eT
LcgIca8gZxp79nv5WTgUQmBl63rynmpB+ozcsvhkM9VNgdo9691TsQhBPfWSjlaA/Mq2XAScEoTX
O8pxKBFM0PzMhRksW3NSlf5S35zJFrfzE78DwWJZRoO2rbRnBmB0e9oi2sEqELkhNze3G7zj4xEr
RNQ/CgAwE0oQue3RaSU6V5PvC6FSf29auQkMjIKX0SnGJv+guS7JxFktHIWDimJti3/QNNW1KrvY
3yBxaiZLxteu+nC4yK50dQhKPA6Acmk3C4WOCtTpMoiQj5tJIceOwKmhprTfaA8lr5KoCuPe+NL0
YRgglU6LP4/xTzh7RMHAPrMgi3HMUVrNL5GEDCzS7zC+sncBYFcWwRWmpoNeLhdx2YCD28R1KZqV
lZASaGayWspjgrZO2tLWs57jYZxdtHrpUNDyQNl9y9isVKWjJJr3iduIVgouYM9/2Kxax7Go5E0C
jBaibRst2Fv1seVOP5Dzvg+54C2+23F4u+EWW3NKxlZiD0gGQPN/r99nrOn/dlpFfVDkrIMe3uXv
rTFY6D0xlYUiMVsQAIYwsB5Rh46nJZbQ4Lyv8mg4CMuZsaD5Vr3rld1quFu0pjXTiWhIg8lGZWza
T/lVPLiNFY58ocsqEHpsSGT90SKR/FYuNhLtSedV0elhgeM4HoSjxTWeJseUZFi8ik+MhhICrHfk
Cz0z23RYhbaqrXqrxU3ok6LPL0MCIAksGa2WBgvuYBCaQR2AXhydiB4gnn0YDQPUx5/0AAOjb7C2
TDINKWsTjOYGKrrqdKG34zYsw27ia8Zz5hZb4+eaX8adXQA7boN0fGalN37JEBN3nsuMiS/lhj5o
D2mKGA9tGpahWkl/8kUvk9sS9vr9fovvd6pn/7D2ahmw4ARHBZIxcXRKFPiozs3g02FFGaRovkup
8FNy7nvuL4GP/sCJSatz6rA+nlwmqYIsnjB23c6t13AZdzD3SbstMv93UaG0K5Fa/Sp38tlEXPFa
q7966gR0+OFC+PnEa8H3K77kgxwlzdg0phkK4dz9aVEfL3zmxbp7VX/MbfdO9ZJAZ9f8Eh9QaCws
VtmK3KHDwxIVgPVmqKODV2U9x/l6AnFy+pNEqOXuP/1/D5peoLlpGPs+gdbBQmRKA7f3H09094aA
UgCuHTB/jAOPwQLhaYF/28PQqCPYShad+YlmAOjxSEOwMiLsEP/qii6cW4EyL1wJ/Jt3zQZ+2CUJ
TrDq1lW1HDbYj4/0U9tpl6C0YUAzaCvj9qGPPJh6th3H9yZMvv9JOBawwektAvVUoBKa1ARrtfir
Dal0FTyh1hh3kVUajyPCjnshMEUvERZOkEuAVuh90ZGoQrMkVIwJDs9H+Z7DNmOt32L18s2I+g+m
Swpwa5m1sJLKMQg+n/U+Gtj+Y0Z87V4UsUaYV+yDr8UkDe0TIXHgJ5yN1u8xJZ0jUGMhrm6eXaGZ
t1tU+JYasbfObboHmIDXWHavPH14QR5OOmAbJKWWC66xZR3w111xspnaqjN4ROBwYB9bcKZeMGAv
2QRwd5S3niMGUVe3E+h7seEruqR9ixNJWQTVx02wUipWhRsAG9hv+GaWECjwI5/9QMgLo3iUOMji
QgM8htCUwmymTDXBockh5ZFPGRE5ObiHz25h9KiLjdnI30ryCJI63tBxpfsJlTFU3K6S24xzSY/m
E3TxA/6i2N4NIW/osIKC3KkNcgIZHccXUt4qcRJ+AVuZXrKHBM8bHkscarv1hM6TkEb8mZ+1t945
9YRbrnVHZxogfQ7LOuuWGjVXYoa9xKkQKq60CAxLA/cWRFIW/gfj1c7fZRFdZB3h5+azDm53c6QM
lSgi0DtPP8QGOMsFRClb0EzvIhk+ByAQ4XVou/Wysw+W4RiLi4T4a6xCrlxkdEv03Hilv5lkzV6G
NyDsCylv1AkNYQ33vvPTv5/YIlp66FLLbadPedV7xz96GqmCznYOLfHR9xxBomD9SFg4wd4w6evb
QkRKSJowsYTzrVbeUiwncCBrXwZs9gIjDrNZEWn0XFo/5C+LRGkBX87lDL8nEzn7Ino8SCtvP98G
8f1NqpZfaAvpObJ2O+8oyW4h+p11VrS7V9BgSAEs9+pqxV5tMJVrYLaatElL/AlT35ADeEQlYND0
qDOVJnwZZ0EX9qe46uDN1cVCHyDLNMjcVMj1FjHohL9ZtemUMRQ1kzSIfyeV/iOk9fZqE92yxijG
MlgtbQrRiYQS46hZpz1/778npciTLQgzrbnClYw058T3Afnvfjm4qaz+d7OGC70BupPonkyJnV3s
ZuD+4L1IwxUEk9DkuQ4eQAdj/kQD01sQ8ydiB/VVQ4Iikgn/jL5QDkCNKAnxePV3LMQZBuwf+JU/
eKJwJyO3sNg2hKlR5PSm1AIhCgng4Cq+yH2HICKKw8DMHTIPIk3TgQCC6zUYBYIkj8q+OUms+p19
+HQnpck3x4/8e9uAk3mRFJpkKGLmGZcRb4mHdFzTPFrbHRG9hEsuAm/BhQ8PJ84Uxb2TtXpOWWPY
NAWvxbPDwugLWUJPBwuYlObUA5RWqDKaw2Vy1NyWaVW6y6NRj62TsTqgArUO75GNnLgkB7Uo8dLL
hnQ4kt8DooWlzXDV1b8NPNQ4CvvZNJMHw0+IFXffau6VOVh+pIr5cPKQrDAZjMG/Kh3dWWJIav7u
YXFL2YpAAbX8gaPN/+zt6iVy/oO5zGbODaryetQGcdwtVXU9FGjbzn7Zt5vLMKs9odfaz9DpcfRD
HIC9bqWi0yzgcS9yBkxhId1/kdkGqf0IbZBUqfafIIyudwDye7REiM0haUxF68UN3fx1bGRz2ZKE
fm5x88VZIHRw8B5m1iMUZ2j+niu489Nta+46/ux4OgGfwfpKvxMPyp3wtY5y3B0idDex+fjHFP30
qTDjNSRafa1mGv+tSqaUKV30WfCQ8M+PXOd4IpSMuZZmqVurRYO4PagI1C4sUEASO6Qh4megxFGX
NGy2mAX3gDFcoLsRVEdy3eZQ9/RQe0EPMgeOBwRkIqMXDhRfBgJAHnYSbB4HZ1k5AWzOxOA4/NG4
LUpbc7nlTPmwr52j2kLjgQn01TQRaDeMmCZKPZbHuUIWFmH9qqYE7xON9/KbzxrPPM0BS6z4yE0L
fKIjpvaWqZTo7Ji/yu96z6QISVrLA1QwsZQchS3DrIYb1ZmYoys9iVouvZp8De4mRs8qLaHCCtvt
0lusxGaOX94DKpgAs+4KFc1dggrLSIsmP9ZNJeZ28oiSM0gNcTySAQ+0ws/Hz7qreueg5tyCnu6z
rIUdhxJTCE1+laUaekmzk3fHk2uAkRAYgqSO5O1O7BOgw5ElsyLuP/FV1sUFXGWCcGpJnSlF0kip
M3KVO+Nt5bbRXo59pUg+aGe07oQbaTpgW2ckq9uJ1q2ArA8b8kZAaiW24/Mw8/0gnBvE+HyBo0KB
xcCtATYGFKvouyaBRqFHWTfInjNPeD2B6PoloHZFWK+u6LXltFL4Q0CAvVPQnaJJYdcqx2bR6sS+
6G9JRiA4+cNp7ks4FqGIQw5eWbaUAhhW3XmWLVKs0mJfK8sYNw3r3N9llU7oLKqw4iuncXdK5OZf
mDOQRbqFneua7M/YxUtm6vOZ6Mk+tF/vxfJBgZktZ1IonfxZh/HalSNJSnwskp6jusjDWlX0muYn
mF2TKU0dQ1lLzMH3hDHj+6LO28brL4Jt/sTvIgxkdIxkH+fc4eZ3V6ap3cwqkxAYUbpQ1YiTqe9G
+1L5fNihOhPa+NoK104Lmj+GpSm++j38XsL01EzyvG+FxNPIWpnMs4OH0Rp3fZzowt9GbcZlvNCH
FOLL9XcxvhNx566gngQ4ogbOdt79FHyf4tTBVbn5FL/+t6RlxgP/InVA2WlxlEdttVybotguGhWv
JuOt2fx9v8hnTjYsj7vBWV3dkjSKxaHP1JVoWRcN3v3soG3TFReEX5POhlc3TTPCYFDjilh6BRdK
f62wpgw2x41bNWBmFM57pPyEwVK8WbATpLA8qjH8qeZHY66sJgPRm+K7a8ugkS9s/rlYh0c90A6J
VFcZCYwRtyRfcTjeDmH/+fnRQQntFKJ6Pkr4JJxFdR6k11r0EXXQ1b8t4rTrpMQx8RdCGeQMCf55
FogEOyYOWPde7rA98cJKMetcGJh+tbPnP83nkNaBe13qJ4c50+fbQYvuJr7lmcLLj5lGUHeDtS1P
4AztPfSJYte5vmRFeT7viMi9T8f+ZxunwXr1k6+ClwsUVZmbticV8pMMI9ix0i6vlLKRyQhxGSa4
pPRIIdy+iqEHT5oFyAvk6HAep9rXSWlk/nZyXszhB/v2VOuHdN2DZPoZYbEsYp34KylN9x8zN00k
btCiCg++kAKjxXFayliApFA4gib4MEMtOxYiUgjyJ2jg7HDFHDrGxwOVvrJTR2yWeKv0Khv4kuwC
8Mk8KdWmlYwKfslE/dMY2IIYINn8X5jnv0GuwvvxQNndJMGv5NJVLmzThEVgNwH8mwvDswqAa8zm
qWBSoEunuLiwNtfOtWqkKHpmfQB2MXmhCy/ptTQ2dPlfjXEh/lAxqWjLHhPQwG50jAplQVtue9pK
T7zof5EyvVWN8pESLpSB7J0ZK6x90UEbxRYzzGNIyj3o1qp+lzE/UZVw12Moz8Yx2w239nFzUJHS
hwqS5J2wmuEhi9CwHHIAIIWg/4n0z4o/lJXp7XgRh9T2RrfqBSsaNCLDBr2hBNQyLs+zG5AlAV5W
TxRKjweoEcthfm6qxq6+hI+C1imlrWHaDCK2QPMgn7clqBTUo5ilRpqFd9qtwxMSRcG5iNORsJ2b
mJ2JwfMKgewK216kety4kasRUZ3AiZNXsra9dJkmHfXtzaPL53sa3xaPLBC3NxmFdH1fJ4iOW3Z4
6lfpbW/+pqNRa/kaxuVAYPKXXupTbtw3ch78wVdO3dd2kQ8zaVo6pvI4aEaUbPGsYeGix7xPcAvM
o88OgWdT1eVW3wuAKObG584unpQt6ePfVRA4OTGgSUtLHKPq8Eb+Kyrsph99UPDUzJMOygrPobSI
Ga9ipc7nfTEWjyfpWiP5Ibo2RdQeE5I6E0akhTkKWtgtnbTJrJGCpBQZmY3MVmaEXKZTpJRIJHCh
pBTlaDUU/IGGSAS5C3VOYnqNIzwjvlb0WHvntNqmDAztWYhd0gWwhC2odytwAX7YkwH4Y8QpP1oz
BXPF3PfDMbqUKonhdxi1JYyojX9oyacmoKIEnxu7i+8hTQUKoIatxSCfw5jT/boJNNhIl0qgc43f
07CDTMf0XLibThX7OBi1bVIFT7/RIevAVRCcnLJ9BtKgHMQxboZ3x07PXbcQ1DgK7+VZTA/sDVwb
MLwvKqyz3KJhMzrhk69q3e87M03wCtzS85eVe3MbNqC4FopFBb3D+MfMsk65IHg3llI2h9BCovx9
643eqJa3PTZiQ900oUcA68hgCGU/BbESvkjg2UDohIwN3jIGrnE0NzwHfzGqnhX5z6IH4olfBD2s
c0r1b6UoGNmZIPbSBPzK4lelO/WWx/+30nS2CKLyB/WNVow7j2LZoo762icvcqNWDTHRgf7s2cH+
7oZsWq8/dG9xJjgzTpRfiGc+4w02aC2JQTjbraseuD2kYYBKaWHeipXuqpdUwLv/vKN3UoLZdW4l
vJAtUsGdV7wbOOWALldJo5yRZ4KzF5b6tA5Ywi7APWjqH+5L7VTRa3XCdcTGzKpQR2H30aAHBcHO
7X6v/tWHWHmjs10ZNJSMby6Yone7T5HRo+wSOFy8/0lUraThDvusxHtL9ekyICwolwtfq5KtXSCM
vadcbga9x+65oIH4NMDT+mXhppjJCRqRzjFqd4lnFOLuHUWc9svANrkKrqH2IKN8VIDdCUM5mSry
0kj7JLZ6xi2XREQQc4pkrdqzvN6k+jqMrUvzgnhH0bHl6GGTJYBfV3d+bNjJhtNF2TndzTBrOCN0
/3MHXO3DlVM0ClB0Ev+gOtU6GGgsZzJbvyqDjhfh6A/aXMyVNmrJn4l8bcBTT7zyz6HCshJNjSGP
5852/W7AccFesk0Wn+qMRAxwJztDY1Ct+d5IcwViZcGI/qyAoBUhqCAWMo07OlLTnn+dmgCKIX5n
O0vYhnzWyUvjcgIBKMpUlnWTy2oBVxGVJnQjKNpzMqqOfF6cqaFOLxh1gKkD7hM9/4F6VRQozRuX
Ifftpl+kUimA0ISDJ2b8CHHxpe9BpaMsH4N/xd+4TdY+ZT3VgIP1JxapGm4OnHvgWY8yZ/cZGr9A
IOGCUurbxgQDdqh8HepK5HnCspgtHlml3awTzUeVDOsieOJ2mXLV8WEwFTQOMYpy69qevR1MkeB7
OWmqFIA/wnTowVMJo5e5sjJb+aTATHquXwkOwMY5NJNwSD9h2IhCgCiB0cSQtH0vUrq5Hf9LH0Cs
dFZ35GvGYya6xAXnoWPVDg5zj8w0VT6BH1i1TvO4THZQG11383OUe0acr+RPaJo/snlh9I03ekA0
ZtZTGOX8Zbv2u/gjiYu59zzr1S9E1W6JgMbgnbv3m2k0f+m5kKqYzLU18nsXKtsm0xt1TCQ0kyvM
CZ8SBYACyVy42VRwegk2sTHUGIkVv/FIIAoGbxR3QqeQyz1AEUcKeYl2LDD4ivjL/WZuKK8Hvlnr
iecGf7VuxLu7HYYcQ8GGiJQi/GAxnWp3CtkqkZ7HWfXxd6MHU+vmveRH+Sj+YnWjM9wZRUP1NdVn
VYWTAnTbVjFnDu0FfSudjn2cH5ZOCdhvvU3A6kYCIVtuJipgf4C06TUsBflEe99V9y1RD/7bygfT
1yAq79VGXJxcjnV5+PrUhbKLQLrKjNuYvOI/YtWaeHHDwZ8JIVsj9oh1zdSE1xm8c30y6gN6ooXS
iXXbQnRAR/UGWR1N6bC2XiwR2/EAQUxHzBItUPPmb9l/9dyzq/0/2fLINxdK7bk4rw85T0M+9Okv
JNzcj4q2vwZKcQdTRtSFtuNjsm3o4OiCCOLGn3E8J1F8bi+fEcOV/WGYbyrMHSAw51QUfCIaIb/+
Ne/J9TE2JefVBzUTcqVUAyalHqdCSNm40wOTvTJCSyzPI7vro08SOPFVqRkSH7CxZYa9Ig6SXitD
wp+mOyBklSHOSbuyZQLYHvPu7pd/36QIfb3QzKQipQYiL+QO5rnxKnUP9XoDDkojHrque+EO7o4Y
C5IwgkhQuPIarBs6QGvIZuGGXz3aEAMcNfoPVrJQuUUxkYTKCXu56F+QmFb3vJTURM/BXyNlOYrh
ajaFjD+JL2BXqmNP9LI82QOHH9mTDHmRH11UVHwrLKH8LtHAaO7NbY34IhrG4N6KXoPB0tZsSfeX
jNEhrwL6d0wIFh6bgq88oNHfIuWVPXn7FvVR/0ogTfBam6lujNMc6caiFAI/ijfZ4eDzgtRZUNcS
u/Esl4i5dlJLK2j6sowCxDtPbzdOvloaN5jFIilVPhCPNgroI3jvZh55ovT8nDjpovqRt9hTvR3f
lnSvAyiVr0fZzJUqJrh3yjj5ho8eTwBGSfS9GUbDIgrKyyAZgtzS6Ur6EtU8lveW9znykHx/BekO
9VnQ3KwEjSeBDPxLjUah3Iy69EvDUT8oP3VPmBfmeJNoltayghLQ6qhciGLwwrotfJL272I49mFm
pErmUOPSGGK+zPtwhMVhw6nwhbHNXdbZUm5Y9SsFDQjbEQb6IwmEoxEqItXeMDRU0zeOL6JEWcPk
AAwYj8w5DKH4zci/36fCbxnr3K6kAUEgV6D9EQW0RmTBLAm4WCv90IUYEg+qQmBcIh9OdQUfwmwZ
ASHP2ucqWahktX/7DmQ42wjYEkBtI5Rs0dJR4bUna3f+5X9MSXNjQ408tHinF4jU5T2jDXRDTnjU
meq1IRpjNSvoB9s3gUXCWlb2Xl1yrKWv0ukx4SXFLrMkhiD6QNoUcanf/4zmmOvP7pLnJY+/JS33
69JIHTCklCgRBcWPh/MtpL7YoEVUCD85wZgd9Xi2oJ9Dn04rBcivPOn0l098mL31bxwFDxKASCqn
6FN4I/PCOQP+ah/xrXOkoJ4NOGOcNK1ZQHzrTp00dLc4Dkh5AgMO4l0OrLO1iEqfk/Un54nc84G2
wkMiss52nfwdTMiPHzSQd92r/1RlXhN2JQ34ifOs+F5GmotSF96TUxFf2J4W0HPZ+QeL6oYzlpW8
888u6uPoB1pYYbuSS0PPAWjVg1s1Dl2M+A7XOGzE0DWDCPIkRUUNJQTk9/iOhTQPNXdMJ+DNy+JY
jUxfQh6h1mSLyS5wqNKCZKxcSBh4RaKAPSuUL30dkuMVz0Dy7Pb0cVstpt1/72XeNOlQt9NhdqkH
SRyEch2GnCgsl8Ff+349WavMkHfaaJGGCvIiUr9RrEUdZqEE0PRe1SDQ19XkyDgaMKtdzWiXYajy
YoO425AcB73yHfy3qiTYNB70TfgwaFv5dMph+jRlzFZJqho8mJmu8d9IKauy3gHyXctWab3Uc7mO
yz+Ah9KZsB1eqPlDoD9VJQgtmGKeKxfEBXE4Cpd7j+cUwctNZip7Y5Ws5EktDUdBTyk20+QpyPM/
6c6UNO7lwmCQHPbavwn/M+Kie0OhmS/fOAks9YZYUFlAmDls2MLh9EZ0w4529TSTwmH7wCGiglAo
NQrWStcB36NX2mWdjFzXS6VqeZSnpdkNaJoK0eWixw/FORlrstAa4raCzsQk09Rwpx4wR+Pch+bc
fqZZvE4Fd9XhXnAAaIRPl5pf+8/Kj5ObCIc5mePw7VIyb5D9RF2eXO4+H9Qkuo7tPGqthYSWoMUc
bvYDpIbFEHwnwEC8wzE++d3l6divUt2osQoowM+2K0vimj620M6NktX/tx1MtLP6h/bdgBxjn5PJ
OdOyDzmeB7aYJuWNhSwIKLDKrQz7MCdriHea+dw3p+aSV/8RwulnaXqueXpgPqP+mihr+UWES+N2
OIGVOD/Tjx2iPjg07I6XZeCVAorbte7+yenOLoSIw+BbRDoko06WooQNZLjNQSPOa2cvCUiUivHh
YGM0SlIoIjMzfODsoLRHzcTZZD7RmGMxsI1MF5FXkMK3gOpvYV84LVS/tYhTLHyAruqjtwAzcH5t
8e90Fva45gUJb47uDsaWRKRWvNafKOoymm3WajOM+wEfmHTjf8UYyDS1qWlzL2bCO4JwupHbXebt
iG8akaN8ZbclXTzQZmkOqP+GtsshgT5+i/rophVvzUdAbNbW3m89zMvEBZEN9Eo17Qcwton56AgM
aHWcKOyldIvTvrmW9EktxsB+e5T+5o59h56IhlDwVPZmpKv5iBX3n7HSqzVWv7GQ79DEEVpMCV3e
7pkxK3Da+ROOVo7jc/IY0iG27Ypwf8OUusdavscNKvhT5kLf9KvkoxXI31fUOl6dicB/NEOH7OtN
qrJfWxk/o/JVGKNb0PGD/UNUw3XNswQsWf5yxPAlF5ieoil9ofcdEaeyV+E9RrJgtn+9OBIbNnaZ
BattntOne+a4Mj8oP5Oh0kh+FJP4WHQ+yUxzkxDmMAXiIQl+xhrYGXV4zb/DALKJyFkv3no9vxwr
r+HyqbmwDyei0eWkyLgiwDICSTI8OpNUqHDD0I+0ZMUw3Unzvcre+AFRJ8HvMeE/b3CGwNRwVXym
eBtBZ/kDE+tNILGN0fGxQvNRFeEdUNn7BQDytl222NvybWwAnNZoNKZJjsGKOTrsOtiqhOmZfymR
JDWdYU8rE4W7Lmuc76LR+3iGYBfy3VzjnzjYQcGd9wXvJUs0nTjC2fglocpp3klgYAB/12vrKsIb
qbYKa4k7p1eiXZbYiW6FK67I8cMgNiXrijReqHit9SdmL4QrAHLiNQSYbDMr7ddJOoVQOzuBhRLZ
FXDx0f6vQE64y6eLXsqvcQbZKZd7DYIPlzFhHvusZvOLPImKDWCFpnMV4XoRgEX7JQO2ycCm6GHJ
MYakVC+lxcehQALMABWwyGm/TP+I7u3cCa+aOSsw3QFY/OKl0peQHp7a0B6c2akBmp1qxP/pVX0y
P3XZ4/6aQg9O1uK6p2nmcgn30YHM9/82/za8824lkMQqKGhgJ0fdzc0JRonBXt38O+Y1XcO5kq7z
wPwQFm1+/HZpJlKOIkvub03P0EOzuGzp6Ns2VShWIy742aSMEbeu+3gikq/RqMjbJ4Lxea62XsDe
SGqrWTPBHg+YFtp3IH3AprvfH6rku/ZGDRNKSZzM2p9/JTukhvHVqgBk7jmA0vq4QX0W1+6kffCE
sESjBDKKI1RiB3OisHoYi5X8G9xR7V0hGdAugOsJhWrwcnB6FP8mfe3Y5sdRfP2N61duLl9bGVf3
rCEJhAyrBtYcMgymYdLvqh5PMf4BK7Hu8o7Ot6OC/O+cUnfF/a/MwAfjuKkpv+ROoyGATfYVKcz9
gFpmuBXhg0W+7q9vOT79PsVZkvM8eheUpEq3W5rxJ3+cVCNEjkH7EK8SFU/xQulSNbKFN85LYIbO
gs8y+lnA0rbKKk7cHxUOKWa/TmJd23RZX6dWZHvkANZ+HVXWHg0rkW2PIK+ZNmRzRc1pRT/zsAuG
nc7KNhvFEOvlw173vg5pPJBrEjGnftWU6WdwlSWVRCa3DcTAUm5pE3m9Z0DfBEejYs/u/uG3adsi
4jJj+tJgjgSXVeahMwXOUwfR5LcAJsJrbykNHLerXA/aw0mccXEGoZZM7L0zpCmAmCoAVMvp65Ix
Ow6kFmOQFSPAyR4jOPlQEKKi1JKpEf8OMx1q6mW6YMTlnobnDL0g+r9xGxd0UFpom4kGpb/ARjvc
+VsYpkUpwIHv9YmKO/xS0UL8WVAkX7knnTO63wSSV25W7MY5EAmHGQJgJRQHumE7axx9cN1RuIZP
6CqMSsKn5pAnRCY+49KkwneNaZUWT7IxwVP7kwfrpmypW0WT7Jj97KeAbMR6E0CrNH3wz8X0eMKd
14859SoJej5cvSmGFkiU7ZqJdWHbko6K73z+5xWhgSTMKc6kTC44AR4aUaXIx/ciIMxfV7OhRqgB
UD19bJWcIvcK8QJDK9D2pEpWRG+R/IviTzPyYBH6s/wbspH/pROHwjsV8TDx5sCC5pjLlY4K7gN8
Tvm12O3a8CHjZmsjLtXmhrtgUOOz4yTSOhld/X2rH5aig8cABFv5rPsjCVpRw38K2fn4B2V0dv0R
xEmTaOb7sVrTtKudyrJyf0VlA1sbHMavtUgnsPOCS+hPhCzy2CmcAo8We1LP4UuARm4p52lDWhwK
0Jj6dxag4Ja7CbT1xTm3UyInfXcz4AOB8S5ZKa8OzJghf2aXD/QVFUUcNda9rUyyRMgj6+bCh812
FHhrmgg/DjsxIB+aF0sJAuQzcafNSmJPlGlqiVzSLLImkgdjxWO5NS8hO0BscDAU6cjMurKn/BeD
T46Kv+cpESdcn6vHRZ7EPbBpKoVa705gW91ih0af/GSABgdJg4yYFlv1CVYzfXGLdJ1EFAtJjdJB
Km7KYz9oAy5ixVPyF1bC9Pee9X0pZ+VWfQqMP0BFgO5rw5JftuSA/7Da1rGmXh5y2uZF+cs3WEDa
dnnS5A1mlTSQktohP1lni0Z1myzO4gHKHYCo0HKmeiN1iaJS/9vgpxdmyVl5qRfDMsXY0VQ+TZ84
+T3pmdb8c66s0JBL6CtJAdLfLfipoCyokVpAkfiuQlR+0NOq4jxD5HROfswO42EPB4wMI++/9Tty
vFRVQQrQk4g6lzUe+gAZFd4+05nO0gpvq6KoVD0FaxtUu6O/Upk4jiOeK70S55HS1l7MLocYuX7v
0gVe/vCFD0qBJlF32TJqSHN/SoRYvTcVe6HYjarS2WZ3J6+n6NTGbASioMJgUF3nEk+eYB7hF14X
H6O/v3HH2ilSw6239PG8yuTA/dxH8LquBvri58V4B38ysPYtFSyPMBpWTsDcMY4dZHXqy3EdcrDw
lHJHGrXb3UnuZ+TO5Gcz46Rk5ER8wbmDcW5kML1nACcR1gYQRT14ARy4ER5hTvCp3nnYi4E698wA
336d+W9iL/LkTJSIXyfhVKMMgNv+cNmJULyaedi+MTW5+G9LS1hGyR1Mx6JgL/W7ToDq17ok6e3b
8cUkSm++nUiumVfWjg6w23I6lTT6lxBlbkHRpbAIrTOQG2WZ/LkZR5aeEgKOaAM8ZEL+vi5+Tbc8
8zfJ0yGzUDnAV5vmxK9Bg5meTfxMUIp6c3o9/A5q58Wh+PXjsUlFC2ZT7Ae0kNvIrccww2ixYW01
RSJA33BDjtoheH175iISlby0r9QODCInWrD/0ASxW9DuqEviDzXivaRoDvSvU3FxMvVbQd4fe/3M
lKBwtAmFdeIWXUX470T6H1c8UAuz/LLzJehp+a4no7K7FGm3+IyrPUL4IOUoxxeOcBgMczbe3GIR
3tC8nYrRTj7H7h/f5KzY3u89g4on1YI9Pr0wp4PSgPQBvaqvPFU6VQfiqTykY7GWgMoYo7fRgx+5
Tvk15DyA5VqwAIKYnMF6YrtnzjE6wURRNRK6hQ2xROfYCsjeYySfcyp19pIo3OczK0/G0vWP4G0O
ZGZ8sdznnrG7C1dsRbl10Szu6Wr8Uq0vmYtKoynTSUy9at5Z3O0ZbZjsq+2rbiRh6U2tZybhuzvu
7YB+wB2vBiJjallIeGIDwu7121cpWKCqexVRL+v2tPGZl3gXyUB2aN8WClnBm+F248+DrjvqMGGQ
utyW+qIh8jkg6sHd5zya9F41ZWzPITRewHtCinaO7gbmlUmVnUbUwby5OBpCg3A+PulXSFi1vMqE
NQkJbE1dZ7e07aSeMl2TSqQFvYDKyDLo5DgVo6LWRNenJAJbB6y6bRl5HUcuhce7Fl7YDGUU/Cpz
cti7nJLxnvxMf40Aktr3buS+7XDhz7/pZf5CR4Ch4okcUmhCpDwqcPV2b4t7JauodOXMIcbXG8Wr
O0z5uLy1Uf4L1btjpS1XF5fKk4POg0ww3BlPAeLTq+QjWrmMvCAJrb9bil2//gtTr//Hiv201Vaj
kSIxJnR+VsDvAM1XFqK/AjEMIyn7/ZnMPRtE/7YqqVC2lw3tDtnFLXNSpgk6N7Efk+vpzhNMwEeS
c8TuplmD7Ayqs9nHDtWjjpAcgyAR3Be9ooR0ruxA2S5r3dFqEn1vKrMI8Rx9aE6kYht3/J06MFFT
ajddBJL9VeNGDib10jylBLufyp1VBsfbSOCo/SnaR4GiPLiJ8xdsYSiwHiK/rDBZlWw7PZrkV9c9
Xq50HNLf/M1wG+9r1PO+FEtZDS4Y2Kd4eLB3XrmNG8liextbs8B4dAAlSxteagkOJPUZtCygu+I1
RFUBWix7OmYthTObQRsUuCGAEZS6pMuJmysIwnB53WQk9BqJGgdafsPKyNbYHUJzZnm9pqGFC6w6
IcI+D/WKkleubga1jcSa4CAlvIFgF0WLnVx83Vqkmt68iftiQJ4Zo30kKt/2bMRhbPQbO1Dd6Apf
kSimM0H+bB2PmZZY58Mc57L+7IVnmOu7cbFtv9/K+c50+X1nrRpQDyGKXtSWDyGUSTcbd5+b1c6r
YrpHBHLBb+LqqdM7C0FQJGJdVlqnCmiCVuLKPNR8kY4BWywwcOYPnTDV30o7OIOZ/XoZOnNTR0/G
BzzaqYWH9L3Cup8uTRli13pFoyxT26IIR9FxR8tR2s4u6+jwSuvjU2DFMMbU8DST9QGu686bwmm8
SYxbHafPQaGka+MlM6dq13k9XX/NR14feVVJ8rSds+CYmJajKmcmLDKXnEkgL7qu2xSB4Q4wxW7G
7Xg1Q4Zh0WWNJ4ltlBEQtAZUNRDJYsoPQCeGiqMsQj4gX5/bqh39+FlAp8/+9wFa2j0vx13IoiQf
rTf01J3LZ9NjTFewOjNcOc3i35MKW2NY+r/NM+WXLBgWVCV8LUYzBhBkZMjXl9VxPKE+auaj4GTi
elobFweB5ezFvKwncpgCMyQD5SSHfSh9XXZjlBE+DtQjhBsS+C0smZaz7+LPq0mQ6hI0/lRBBn9W
CizjXo4MSkty5+kFPpqlW5R95la9MtLoBVZCkdBkKKcpivTQ7OEErUYJg6MCwSkfdLdDgYpgl1FI
wXtLBCqEUptgC9Jf9TLwQC91yHx5o+k6dl98klC1jjp2TlXpfJt70tflezkYrp/gPVtOAB606E/L
Q3wDRKmjhvTUGOVaHQiU4VnDycnPgfqTGG2vMv9rMj7QBKhLqNgnvGpu8qkzWY46EvFjFfIFsCj3
Dd0yvAK7UmvusXkBZygpsxMA2pGwZmaOgoKcwj+ifu3dtXgHfompTGjEXiV14Ikady9HbsS5uvGJ
6jIZZxhmx1wtdyvarEhSRWNPcZd7QQlZh1gJnsJOUohuZcO5crTix/RM7SHtkI4SFdpmEgXwCKWC
XXrSY9YWj6YCb5qcmtmsLa+yFau2UZ5ywO8xxEXfYIDgWA4SkbtTCiOEPGp4+PBqhS9+1X8ftvhp
iiWEH8bRAyBniTQp2c8493xcNgcT+WqD71YNsEZ+8tISfwRkVn+1bUOrZko5rdWaXNfZAEAFmNFg
NWp290Fs42jVE6kPjxXgmXtwpe11ia5x3OJHeDherLQkDdPjje9bjTPgdGcRw1i0sn4rNnVhu2nV
Vlt5Q7mqb9U43BzdDo4oIDs7iK0SzFvSI6GlYqIm8NvSZzWp6VnqHZCPgHLxUyfy0i3ay65HDeGC
2nmlGJoZS+cixaXJklJ896CKUXSVSg2eiu6bvXYrTsZSiNsYBlxg8CZZo7xC5u2LkETTYaCPaeQR
MROXgQZfSxIiUYSmdEVI5SAxuX5in6ggappvZ4SSVPmPQqZaIf8UgtJMUXHD/uO13QVHqI3AFOUc
L03VBN+M1et8owRsyA2DwPoNKTe/ylIdk4yN2zADAuJfEVWUjIDpQTbzk7z9cqdc2sdhrXCjAqco
rhTSDufUvfZEJ25CXYv+HvZYFemO9uRmjb13sFDEb1VRxF606aKrt4Emagb8mZSdR+CUzW96Atza
14i9uCOcplOSQ5imGMLbUvGbVg8Eq75SrB5Aoprr8vZ2oopWNu0vq+qpoo/UAaJ6fUFMPhKI74YF
Ewoe5eH8dqWwZjerZIEcb+4e1ZQxucoRHq6JfltSaL2RgV55JWidDhcWXenNECee7Gi5cKa4Y/0c
NVtjdJwoVWUcBrTxOBqySZU1smEJvLCtkqVD5IX7C6EfMUQuCy8rvu0sIBRP4pS7CaSRnRH6rESv
HO2kAF+aBYATHTg63lULZwc2fszc8zQc5I35jDisZZfRDii2XwXashGCSaUSF20sh81hNhuitdUG
7W2EtxCjXzb9OiZORBpepHP7ohht8jV2piHX3idl9BaElaAfArIVLNxASc1sLcsgPnTYIE2+EizZ
5ITjFAPDoHEjUx3r/YVnn0sL5OkDFQXrpdtrgHiuRppW1tLx1VBnxjAgXiL4fjV/4IktYGCeTh/q
xDkecpG6hNQhjd4UkJVy2p1+Q5eNwPQgwK+RZ6eJEzl1B8qLaFeA1Qti5+5ok0Lgr1z/Jm0QXRDJ
fMD9SeoJDE4dRQvPBSN6AaWE2o3O2PjFIcCtEMJqEdQtTfVJPDw6/BAVfxwU9WUP1eA9v9T1c5eI
fwhuZRsRBaULzwuQQwirZlJEWS6MCLcmOxK5Rw6mnGOuRY+22Eev6EM0FCH44FNLMTWETUZ6W3xh
bkNMzdHZodz21Bq4od+czokQrBtMk6aKNZJlQ3e6jKPVi035RSPVeXrRp7rFuUi58uISGTlJXY0b
OuOkt89iILW5G5sMC0Eoj1j6ldvkn4dgijIYgxuxNU8omKoAwOBhOGdMDgykPTKuoxDiTp4g3CCq
7zczcFpDBTyxTaNF1IZZ99FCHsIx68RQMmPMASm3Gz/EKVhzbFYoVz0Q2fOW8njMK8MwitObUu56
wKkBOvdeurjU01N8BfDM2uqa0zyoiDRnoYfFo8TKOt9OzlMPSiyg1d/e7Mar6ne8bdZ4/ytb/v2e
1KKPZ7cvEYXVAx6i6tj0bqjWYp2KlNFqJNTZ+8yvbyj6s50wOGmwryLVAqKPQMNusECRzYEtO84f
AbqRXPyUvrfycZB3g8FRfRb/5dfmfTjVb6XIGjDS1NgGVxvHIsr2Kb/rOsNZDXIynpvWrDRqAtQB
Hk3kZK9Oatq+pce0rei2neKBKpoPTvlaWKnTK5Rwd2uPEiuYVgdZX70WTCvVMxETXuZQiAKVNLTK
jHUKrpdsuklkOBN45UGYcjaPw0RrvKd/c/JMBbaVkoHCrPhvv4f2+Gah73bWBWnX/mBWVq4X1KvE
IKRIkwyTGxvqotsOyVmC21LTXEJmgtMW3oOMEC6HcAmSME+9sisYVorxHNk0pH3jCtoPp9vLHIgS
YMw2ZJu5fsICFdox2n9lTdo6xwlqplck2EVkPji7B0kbHQpjOAWSqS8Bj22BlhAMNeqmXYADCIaQ
gYCZ/EeeTSag4ltD8AK7gusYWB0f26DtmTckUxqMJJg+5bJJcSyJ/G9zXfHUf2Ic4Uvo4Zok4hQ3
wQ2scJPD4l9kgvmG79GrCohVGY3cr/7cHPox8V5hn83zk8SgwRrs3ccLAwImcSI4JAUz7I4qEQFN
/VJH80guKoSsbZERpoqGVnVZXG+7TatJ9twJL3yOKJ7D6+cKujryiSEbeKEIJUqvXZngqknKvTmE
utp+Ej8PKgnvOW+GTxU3LLqZPZt20Jdbmr0q9FiP7wSmugMz7cq4n8EvnTj2aqxl8JsSxnGDzsnx
da14aZYD3M3hnZjuy0tje4gnK9VRPnjDOj6o7lamn01jYtpEe9e8xBE8UGCui9LQzQ61wa75mS/p
37yxH5goOYZ/P9AJBc6m7Bprq0q1bafQbd9jwZQi73Klw6z0yRpYk+2shGBm3+qKTJvb6EW68XnD
FRHnxvpYV4JsJlJQPcb5dBqF6IIlUpxkJ0TADxOLFwW6P8doYZ0Io8ARhjg+KnBTkvX5eSbNknBe
oWWmpsAWyh53eVspvjRedv/NG5hK7EXIPhy9LT4Fs9osuCsOunk9aI+JZ/355+uDr6AjZeIfHFeN
apzxQ5k+vMmJ7zjS7GwXlMNPYq4/FkkmZjUbV3pNx+AP1KoG1/6wQt8lArOVhEPvmpUYJ8bfX8sX
OpYFFF5L4QNx1QSi39t4mAEQjxyaF67E1Pv0+67c6UDIHntiFKde8vJHwLV0wG87hhIKklgfAOwf
fA5450Mkwf8OlC9qx0Xi+dbs2xMDWJmDVBIVzHqVzASHJUR6HT3jeXIkZemb2nHm117Q71I6dVEh
2HzRzyRo826l9OGsmXgl8BDBBbWyJCkFftz2yvHZ8JjJWhODRQz5Vv85aXR+XrvRYf3rOpGjwh1U
t/SpsKVSH+zGBwzeRJnLFDLEZO79RLCcfdplMKTX/fT5Z7zTT5oqVG/LOSqwkXBkTUucb4hQ5hMK
bX3EOxsUfnFW7HqJ2eAnGeC25feqR8+hX11/cAE+Oc0apA40AShMF/J1XD66BICY4L0Elyjk++yY
Gbtg9ajqlP3Wmi8m+ObqLCBSFKWQk48+Ig/LQ7kTc/H+fqZsO9heoq7XVVXj4U82Qa9rDwa34liL
rcFC3Vs0uZExlm+IYXQhi4AuteuKEGJtQ4MkrcGcnZTbUzVtj0XvandoL/oH5WDQQNxibsZckANZ
vjmLMbn9DBUhoeobnu40Ud8Bl5Lb2CoxdUcrE0J5M31Tb3OY7NspCsS3B1E3jUysd+2J74Xk1d6X
HGXT2QM2qQqtgcWrP9EsegNWgNGYRDJS15sABlQT92md7lTiP5CGvHYt5eCNGBjfigtqmkWKPunN
usjAi+MuQPwWWUqeFnjaPr5eYLLJNGyX3Jj0HXkQIyudsxjymLQMxx7xtuS9CDTbz2izbzWP2JqA
thr9DunMiId8FEV5pEonfD6JXJUDEgBPVJhlaYYHc74p1gY+1ZUzNFg9lpjYH8PGkFD/ttKk6DxT
Xy/ojIjb2C+Atm/Owy6pby+nj4/iSOjlk8YOVylFAUnMwW+gPO/4Q0EynuIQjOCgXoBZAlwZo56P
wAvd3EtJ11Zi5t9q9/bG5qVzq9RgURO6UoqmgSVGztTBRUOkbrJm4RjF4RD2RPqlifI011wtB8/P
MHmfqvjQqtFQeg2XLdfM71WHPvykLt1mSx2lHQIe3USsus3mTjfgr53hxvAeLOxmpXz0TeDe9D7f
OOnXynsLZwnCkd16d4JH0tlzA07mKxoRs3E01V+nydLUKBesZNq0renNkAhGzUcnrs5G7sZnqHEs
nbmA+FtGQM8P+m2faWqPP+8ILIZIEBpaBDMK/N3VBrfSvDFlGlWNYpUwUygy2xjETAnjOURf760e
MUyE1PcJgkMwy8R6LX8/g7X0Sstd+VSSCO6jnVIXdY7+fYtQDFI8Q5xBRaI0B1Ch0aC6q+/w/l/j
fY19hwcRBmxTcZ0srvbK/hTHspz/dv20+PG6yiCcrPE5HXHwyI3NyAUy0e2amzZHv2GwuAkjnl5c
jgo7R5YfRvwOOwK44pLVhT5y9W7VIsCpRuN1LUzZOOtJwURSRM2919+6njxDQZmmRPubfoD2KU1B
W9hqlpQInGLtS6mykRWh2eUZHkgafyukbPasMPDQfHOOKvgdmgFd6JhZJuqL2aJYDK8Y/gyVYmoT
lZOqbjQmhggzsr5rJWsO2ge6V7Iifr7VetkwMIUn5Ji3tmlEp2mwmDb1lyXqFGWdV6B53xyzWNzZ
9zzV/R29Qcqya1VVVRYHPEIil0hYBnAvDY3n3fBg/NiSfMLyvmNn69SVT2ByiAv0DXrF47N7VGw+
cMClp8XzeP3yAzYmqgDKfBTicm0ebTc0D5CY5HsUX7YrFhcStly1EJRzu6ngHG4VBTxhS3vIbTsE
Ofva29KIyjnDjeKd7cKxK9XJGUbmZu6cpaBHR7Q9U76vZgPv4GYQpkd+0Q0sHGJd33iYAW0i7R1c
AhSXw0Qz14aGmUaAz0ccZU8pVsSVjS/Dq83f4zc/6E+gfVemgPId2O56g86QzvKpsHyea9s+NdlE
De6cHJvH+GCMw81ugktn9jJlkUbv5etdoA1hnDrRMhUPHt5lySnshje9hDm7+aLAoIuZSru0AvEM
JGNyJVliWhK5YKS3FfMCUdp/Ox+3Vcgj7XCR1jdhZ2uSDtYAnGvGj8d1+kuV5cItOB74zAv6vL/W
U+6UFZdM4Q6fU0sMzX/lAWmEg3MOZ6qTjpBYj+FwIWi6Jz8KLgD+0n8YRgsVJFKEgSscyV2z9oz6
3ZS9B+XGms0dszIVWLa8cu0SYKpY3BIPixZi2zhqKoSqQqQDzVB/cVBE5OjDBY4jmk4h7n+loMzr
lt6nSjCoK79u+Oz/WWCoNhJUSUPCppd9eN+HNvAw+zzDiJcDNPPvLsbQIfJn3eLfsGMKJPhxEWhy
Sz6gIhfpz+LpWO16noCnowOW6o54f0RuEjpf4rnRVUp52ZCBo11NqIUNtTl2tnqBaCPrU/NpEAUp
DDNfKCty/8rpkNYMOjVKC14fxUdLtNx4pnRFFIUdEOtOlz15ara9UCKF0RE6DJdVrFfGMfIOi9Y0
q+pf91//p0x9MSUJAxYzD16+hd5gptmkCzaxYK7gVVPuFbzaED9nieWkPFEbatefrhWOOnsM06Zg
sseIsOMtIHALINZWiTsb+fSII2+kgMMajGHIGw8qR0bpjQYV446Ifrybh1sK5OCO/xC70GM/5VXb
ipeynUi6tUiiub5yZeeF2xGqyOuxHwgb83+NDWneSln7E/osM3bWDCshS4WZBM64dekzzOmouE+G
vN//4+tXV/2sP9ig9gMsf70IgVirGYpCyrSIYDkiqI0A3O1wvlHMkx/5iHEztPhHFVv+RMzFpKNK
NHNVAZg+gDRkDmH799BgjvGBetEjnb6Dw0sLTmy+H5kfSR+ueeQBT7PNbnEtSsQw/pTc9xP8rzK7
pNdmTHLf4V35khd03crfNXWFe6JVw3bMSDJRMOvdLcW5MualJeapvDzm/5Wmf7cNA8vTfRrmU4f4
p3q+2dybRMra4x0KpxgP+P4EqQ0OwVke3p4CV04MtT6VY1vhlfNthU/XAppeN6SMd8LOsHGmk6H8
V6y2+hPjevSKZuun6bjMcCGXBkN35NdYImren2C6AnuXByjEXV306Mw6iCJaVB5y/X/OqHrE5MHF
H1GNdijTxwKeEorKiiewMx3UUVwGsrDFO/T8iUJuDZaE3KjE0xCgHKcTZgDcCiJ1Zzv5EKZ3flGB
W9FAJLMpXKq430nBiOMHhSXK6YlxMuutEB1dIvo1NUTTYAH94BTh4i3jgZfO3ma6Qc9GzOqjL8At
69jV3zyzsb4aV82wzGPYvEKYFl7CR+7DPTA5E+OdaqvrfXKA81Gg5IaAWNzy2TVe3J0892afh2Oq
MDVEZV2cflJyjtwfNd3ghBmWT8MmjSyX2hPIGe+PTHGaRh1bvmzcnzp78Gpw1SmkAi5MgTh40pHJ
+CnpRwXvFHbrifMonDlImrJmTKY3oH8cz3QFBf6SqTmHDg3vQPcrSode/nNHzNanMxJv/xKLSjji
OqTbeAAmbkrSU30Lhkh5XldjX63RVoGOJ+pi/cElNskeYIkcVlI3dl8P848KWx+uTm8E77w6IZ0x
gTVliGMdKb0MyjEdhChp1X4U7LNZ5FdGUUsBdDsPFKgYMLaTB2UoDcTPa2UxLA4aFUzEDtZ+kSTK
3sjZvIQVP/c2fbP++O7BodH+DwO0ugRvQXENySs4nBWSsbAdxm/xusgYJjfD91YGjbcgPxDkmrRz
n54Ezr+UMM4BnRf+fo0w3GJY1QuNt1ogCBzmRbl8MfMMhzE/17pDhI5NPade3P1LtoSxkDBepiQ6
HQi+RneRbK3L+S05mp5z7FXzbtiUQaTfDaKscfhA7c9AZGfecXh2cer2kclq4FgBdWfyJE6Adj17
MrSg0vcbgq65nxS8rHhkQArIFhr031g5/s3Z9fwQWz8R3yY10+44nW2pMa6yVwvyI7+rU2ou1uwz
XC8bTNHlOCVHmtcATGN7+Vb2e2/VQYN+MVAKvd+VAMOzIV8dY6e87/dbwv3WdVYYfJiphxFrli4Q
wNTsTen26HnW8PQ37TjwXFbHT8VEtANwS0HyCXV6RZOIiQbDjODQhYWj2vPRrIGSBWo44m0NITYO
9DVuZQuEC5L4TGx6XYdRClt4Y3hhlqFb/elMxjhFCUA+AAF/YzZz/ij+N6FUwIdQX4CiEA4InVdD
DyGlYL8wzkBheCM6+OmdfpOuEXVOhP+dijJAUaw19pZxQ+XsFTWpJ6A4rww02mUlaj2tmqhV7b9n
wfHAhTpVcx6JEXI4NQIjzs4Eb39W5j6cG7bLCsoMMiUWaNQoP1lTMdS+Y4P56QzFEMz4HCW1QA2q
V4PFMWS/ZP018GNE8BFJRaCQI8qud5K8I6q4EoT6g2Zp5ZWSQjDAQ73CXcY9xF9DvTodGxNj0OJS
OD2dYcnabrA6QjIur2lrOKGcTPH/VmJjkp87dlCKyWX4cz/9NgzYBfxiNfHMimkJxGb2vvpbZF2H
bOVjbfFpKBfXK2LnNUZCwAJaIcx3MexEmtYD+zr5yy+dYoPC0tbDc49D7cLunNFFoW25BY46rlfG
si7igLvWi2sgD1hS2FV3g5laIAY9akUxWLAZDXTRVQUn47k49+vkdTms7WPVaS2myfoSbok6vChj
+5pvgE1cBkhe3i1Y96BRLQTqnZ/s7PxRn4uGe3qtEIXYcLXAaMLu0Q0b+4wFDAIayBCC8AQITZf5
Lv+9a3nE+kHniUg/v0pYs9wTvRU8RP6HrFMugvM4X8jgC0f3CnG8jQRL4udaog355tyl4Mv7yLOh
7h664l7+nm4+A794vKoKEbKtVbL7mTjWf3dEEFZXl5KGTVlyA4xqg2HRBwhLL7ZA7NwokpshijwO
o2AF56NESWGVQNQCDWiNCeIH32YGjHCxF4wRum1CWtcCf1zyu7+fGh6rZL2j2KoBHUoDAM+bn1+E
xFb6WVW5UQTJdSWCliiTmLSwDyJ+7IGEcbBBrA0YGsj0NZyvmVnOlfM5/tB8ZqCCfmoWNDVkWvCG
HkhYOkC/yG7wqpEmHiB38arkmUsN9eTZv88apDWzdS7T1IR0iPg0U7QdHK8FI7mC0N/LFDGJS0bX
nSCR8Q7mt2e8i/53P4IGZP59UsYy3b5lW8idSeg1T/+DGMU5AcJh2SBGmaHP9/liMQBd4I10idXu
0UXsbD+lDJq7F1REIcISpJAf76m5+ju+4Ors+udrMBLTil87htmn24gHtBkKvA+bQ5Q/t6So1g2C
PAmhX9TGCDi6hBWcSkwJESgmKyawSWdcp2T+A5znPQNMsTUiq/Z+NxoJakZy5LzU5IOEjVV8OsEb
InFVM6CSNiPSXfJwpGcpSRMvImQR/7aaciom3DYDgtcZuUznKehL4xsN9v4NuC4cR69xEipXQiOM
RP4yJW+HS0DMUpeuesszz7njkKeR80ayWG6Swx3yNa22AZkAOYuHyzxXnbK4gox+ramXAdBL7rQ0
lqqcCqMPbEclXm5OdQyS65M0eoZncLwGDz+U0x8e/8ODgwi5e8nWPcEXoiWWuOvm2b8bfmisxJ0H
V58AfUSvAiwOs4rjL5OslVhFQponsu8GGqry0Tvvs2MPfUwmPUzHxPpvZxl/+uWSh1If803+bsqK
vZWyrXdtFS7xTlBZucfHw+8ub38dm2eiSL/xgjhrCAxp3cVR0jWtsLZnPeSwge/pugV7d6qJlDYu
eRfAij1NIYBtTUVH2pSpi6XiFtNRtF7lbbWS5nFYcHkI8KazfBATd7zp7OLPIHY2v3YIXJJ1IG+H
mpoNZO5Eff04OUyPoXc/oU1KFG6Vm+WupvNkvGPkTSq9f+b1AfFY+xwTuCKyHNcN5QKK+hUOPNd6
mausywCbt1KifLu/pdU/JS9PxmFtQdFyl+gmxzvIamYYaKbgdYa2ziHK0IJfO7TcrJkPvrZCqlic
EfeUHUkMLoFb9uJaEhYtGZnxucK22yb8UsfBetKF99pTwpLbeKknwOnJ1pllvHIAluHLNsPi7a/s
SZdDLFRT1F2Qx4eembi8qwnxNIA+qPC4dgLIYIILLB184WClY+H+Lwu3yt5XYv4oQhMsCinl4nS1
f/z+NGPajQHAqp+9yrGm0oSIGPzF2oBOCBZKszbuaeIOECHqqjjcfnaNGzHAaiSgYVgoyW3vMXfI
GITTwRttW+IFwGP7CsH0cf4XbMMUENCgM8D5wt1x5Rhf2d/7R5VjzpBIQV1MvONimbYhTD6AXFXy
G6F0VORFgKwCgtUxjAm7Idc1Cd5R46ciolmP8TYY9cbI13u0gw/b/zlsR1SNjpQKWpPPvihu1U/X
oB7wMVHmyyHRD802UJ9+1w6T6yjyx4LaD6JkqroEKc9TRCE6qLlCCOG/ErNBQzqJqpYTSI7rwCFN
kthwhxKq3oKQKPqmm40G2Qhmo7SlM4d4tzH+dONyGOfm3yB89t72bfMYsQkGItFpdcOHBMk0OVVR
EW1h6BfO+Yf4WoWfopNc815074hpjZo1lAkfRohnCWMEFM2m9McOiviM/JsB72yAoe+NxDZfFPVM
NQVZlLWv8xNJju4Ac5UBqFAqAo/NJReJY7MZgRUqpkOAmRWX3+l/TieFdOQDyaE+kbCqM3BaZTdP
C8JwFqbHozpsehlcqi1b2Bfur1Q0G7srJ/hdbr5KI4PzKgY9Hz0NttNuyFDlE0/cg689w5tWwGRE
ObBOU8XKAi0v46UafQQhspkurCA8XvijURpxE0Yzdc9e0ZkfJjZgRDXRHJ0PUoMcv3grWXmj7hTq
V9mbM4pKWsHSEaAuqy1o6d7bqQqpd40Ehq7q5IaYb1qhfVTNY899pehsM2WsLReJFyRqUpZf7FQt
ow33YqF3Kj71KxCdQgTCQ/hrx3Uz6RXyk1ZTNbic4eZXXFZh1nAWvoGKgGDgNUzfC+GZ9s5VgrfU
uHPsOg1ufyg7X21559THnQhfg+nxgdiDEUhHdDSe8U/cRMFsQSFGDNabFPhW+R9kzTTcpwUViixu
8A+knf69bEjI2rUT0P8X9EwpP39tnHFVD1urABzlyW95OqQmGDY7X2wfQTw+NgWMWLBTYCLVIbjM
u98Vln0ksX5C2x4Q4V5LkcTFc8bQdU7tSdJYHtIkiUzEn8tP+xuS18KtVb9xLZpEiHrF0Ckdk2Nz
N4uM+oWjUuxvdINobCdiJF+bywy7QM4ADoqL0JrPNJy67/V1uT1y0rwbJb0eGqPyzt4kIy/xllk/
FKGU5QxrFAfe0t2wZrIPZjqlbM9Nx0X3kvWIoa/YXNqMXhFiypwfC7qKQFssn1lUIKJudINpXzHm
zq9pcQPlDkjjI22gWFY6FuMvaQY4x06Y7ts/T6txkXxc0C/BtZnPJifyBPUih2/6KUrFuBLeVOou
7dHlaFrAPDGe1cfGUlk2/IaHO6q4sRSxt+UmE78lllBR5Fatzggtin6gswpsdnsZTXcGAOwPpGxf
cBosL7bWEfnYVJMCsV8PU0kdlT684sVvY7GZ7Uin436KZ+9DJ6nMzX1CQIst2LTfj4IodrMUxkZt
JHFY0Fl5drTCdx6lcR4kxNUHZAEa/SVaGK9H3VOXwvQMp1UrwlJ6AO1zNHlYZClUllIXcRdky0oE
jOfbMrfGi4V7o9BM2ewXGzxHJd6gwjgnDkQOeOk3ZLWMISxWjBkWjZIcTCbIikRjQW4DnWPHMle0
qnQIVypHDFqU9eRnSle051h2HzQUDfMOQ7gnfUebmZch3VbjA6XEm5/Ub7vxsM5LJOfgQV9N6dvB
X3iTSJzhLHXr/x1U6Poz9KvNNqPBGP+L10V56MJzoNBsQ9vP1ITdURzx8+cJjB7osd0Exprda5eM
nKum2vNfr997v6VDUavqiiFkCDFUKpdlxSJ0yka+GNKbKTreGhE5hhdVTac92+yz7v1kwzoumzgY
QiLKeKgIW/WDVvM3dTI4rCBbf5s0iXS4FuaKiEnvfppP6lOAcY2Qhq8NEIdj1vMuxLevx2mLK0Oc
isHbcp/6oRMfXHKMOn4HdPOQhx90ZewPrEnwjcJRi9ALcCfDYOisUgwkoGRLej7LTEJ+wkyb7v/F
1X5xPTYbYzqbnR8X9ASnN5Xl2JyKK5BgzXalUuF5zhbzri8ddNIxf94zovKeMoMyZWkeBv6AWRc2
V2tsdAr+QOpGVI7zZVPaHN89+AquumeSDWq8adtrSxIMY5ePmK8vXIU5MNr3/0de3VGkmNSUTuYK
uA/zRB7WgSVFd5o9B2STzCGfs+zuwBraPAacYGsZzdSyw3jbBZHIiBZiJ8oahpvhVnIcFMDI2ngr
3ESccRQHxnNigWg/PEwxpwdpIm/O3AYQCzlytWzhwWiZWvCi/PmuaT/rMcinf/69Xs5g4EqWVoZM
VwXZohK0Sz5a5WBfJWCq1XqKlO/kbwSXUl3t6A4Sdy299oXxg7D/eJqFbAh19ZUdL48SKGOfm45D
vV6pg1wKHj4GFwUvbtyRNYxNE2CZci7i+WZKK9lOEwKGRhsaaG9w93KuqlPSBgvbUJRsRRlOSoM6
UNldG9lhMDwwVndA11jZtFD59aTctarlHOdcFzUCGdjj6/mW2G1cEB+3RXGNQGFAe+ilS5FGQnvX
+R/WhqJCcZJfacO+EriXe3Tgj97xnrgmtA4p630nS8ZImJmnVKlqKSpX/eTB7GljVz3R6RbieZ/w
7wdpP1u/toF5By1jBjzTvFfZL7hiSkHRYjOuZZ6zC3m+t4YQvmFwNPaz+W/DVXq5sYTtA5hn+vHn
IlnEv+WgFrm0cxrSDxWYexs1OzqyT1veAU2HCFU6arK+0NZRNerR1KwXzE1YUBWNFLHTBdbICd0t
8Qdjbp9mDKySNGTAsmmp3JABX5rjqh+MnMYyKC3dm1SBL4ZStu26v8HbBcw+tntZVqeXVZizW/Jt
JmeMVYLgQRbRMdboqG1ClwPz7EUba8yhp6DDB9roWXB5tst+bk5MYV7ZGLW/x/+P16iY68GLgLVc
CjqDN8O7ZWv+Fw6/C9G2LckhvLR41Vz6Ij9pTHyyB3hqw+HHC9Bb/MO44ZZ8nFYVa5eM0tkphR43
SboTsVU8S5JBjiNq+EUr5OMSXhVbkO0AINlyiWN1TJSzLTxLCWRT2MGakPIEoTynxN2beQyZ2QF7
PzFQ1L1rSzWWiD4WJm9t/tXUNVp73RYRss1vzSLbcobVouSoRjhH8uoPSDXZzgRwvIIMCmmQB+KQ
6T79W8HpsypC12lzdNzzzi8/+c0fx4lhgx4DYoNjj5Lb9nfrSFQ5OX9+jJiiBD4bH8BpdSDBb8wU
KpNHLvPx8aQJM7uR1tFtV8LWM+Udoazj/5s42rBbIUgtJCSC5QmDl3RDOD3DguvjgrdVaYgHYK02
S0xZ4BEvA2COjJGP1Aj27uSxycPevm2NC9UU1QCOEZj8/I5Mh3o4+4Ubnusmk5b2wpFHx+ivHksB
ImlSAsub9M2FCDBr4GHnDSkuWyqcmHgtd9aiIBTcO4h7+uXgMAUQk/KeyYqJrahMyCdxmrTAn6bl
bmLBpZ77qQV3upERD56qQH6jUs/pb5eUKBSJRlFjhC8L8iwhpCOlNqloCTGeiKxiyQK7GooPOc5B
IfjE7aYDX5vZrgpSnnjLrqVpJ2b8IcqKszKotIJ5bQCrYPrGnEaWpZJ+CLnEHAJJx070Rakn0dZG
XAKDNPZMpUqnFl/7ExrZpmgS1FeejwM7EVR32ejn3cjT6fDoT78bvhWw04RRRoiLaYJS/4z2nLG3
7uVl/wqlxWc/6/zDPS6wnSD/G0ES0/0tv3LJq7R7DtD5YIGL9o1RULR2zcLGna52rjmeykBTzDLx
Z9XydKoomIyOpC/IMHWTB4joK5qmLKDydIxiXmfY/vpdMptwLjw1U62cfTAHlNDSEZj+EMf0zAQ4
aLGcOuBDaKGvhf2MjRJnXjNbl+yBsbOSFR/3ZpH42vZhgCBjBdz376CyKXB86S7a2FPH46pkuThv
pHECg+UBhfMisH1f4XXdpuA0+mBwY9GZmlvgwPuq4KiIQSSJVDLqThz8ut6tfx5jleBOzykB1QDZ
ecVwRiBHk/h0ZadCsFmEgUSxFUz+tgN7+gpuD6F11D7Ncxj1Ao50l8qKVw+tlqdyJ6QUh8aQhwbH
UA47Utv6Z1PB7iE2+lmGKAFCTAd5HESqqUOAga6AiblvbvheQpiXSeA/b0+ETTEh+ahovxg5m7I0
nbTd/4rl3JtKYe9MspcivWL3w3bEiOO1h/TARbpu8n+dLPFwxgHmCEmcP1QoKtDwRj0T7tEmct/U
DGVkqpjnHQmgb/YW77lGdDMtufc1iXOSkNZxYqWMRqdh0Fm90qr3MTLyfroD8d7PVuphAj7ahDEI
/gzSz74Wt8uyfPePWhNp81RBRMV7Hy6nbMi3Qrc7IPZ70/ke2EIjMlwbwYdPnVZHJqB/Gd1mWKfa
9IXosHYZ7AXABp0k8LDnKm/n+cXDHsaxThUVsITnbM3hJEvULAKZd2zgIZtg2W8C505NNz18wy80
MlGXs8U+dPraJHoFROABX1NXPP7Q5P/UYrHl85OD7Wsv7TwKDxsSFGpvtrIbk/vgtTFu3tYEww6C
/HBJ9KcBYQZb4O2zLvtu6awHQTZe0sp+c2D7FJ3qawgRQB7bRu/Qsdw8/EahyV9tQ++nQiEElRtE
4JNdaS0ZpxZmGhMqM3NfN5Vp3rjMdAAkFSeCJ78bNVv4EkxO2JWvSwP71z43yo1LplT0sTl7j0J6
NRT6XCKCrCHZMueTVc35tTNpmSa03IJ00KPuXdvyvzjzlicqhFfKcxb2V3vw1RCzjs+iLDL7ckgV
Cg10rfmvm2qJCekqtyxQ8kAmdOKy4r9jbZ89W03lVTy72LDMUlFbArqOYXXYXIECzm5dFDro3EvE
HnashWXkV/qUuwWKr34cWehvreP6yIclDxyuUZDMDqTlCe/1yDeNyUadD1kCoEXMNeqlBG3Q9ufU
P5hpoFEbkNMHKf3pvb7Ddw4Cn2V5riweNMw2jx04eMkq/pS2E4r1gGMZsiCkRCfe0G3d7mj1jNc0
+cOpaPKNYED8/XCSXpLXhpKw5RL0cs0EKFs4oVBkJg1AbBRQv7FQshd8/9zUmOBAUy3N4YbEqQQe
47P/Le4F5WEcWlW7oMcIBZ18z6Qvdttsh3GMLGYVZ1g5GALmHeeTwB6+FX1ljS1oUW7VUawklAab
r4B+fb1p//OG9iY4HRluZQj8RLE58tpiDW8ywHFF4Rrem8s7fnqXs8G5WZZ2ysYQeLJPRZihB/aV
Ny4/i5FHwU/43FI5gMfKr8h+4ITALSHPrgYgjZw7qGKpNdxeqbfzpoM/dPccZp0hqBb4ksNV38bY
12MlUvBI9FcTIVOyhUWa58Qd6A/hhyvXodZn33q9grhrQCEVt9Su1y+41YsOzNYIDQVeOXr/4Qs0
p3gNG8pqDFCGI7kaa9SaGp/XjqQqDUL/mePROfVRYcQHJoyT9rQ2jm0n68dw3bIEA4f/eTGYLqyu
x0MOfCWrybrFV92m6tpBAEhoj6U32PMt54LWX6BtqeriPLpwsUw/4RMNkPArnyvbBp995ZLtUuU9
YlzmMgrkmM1ROBOF18Y4MeWOxSTGlPrHlvBi2JqdOQ4Y04gMzeq5k4sobrVFH8MGNnNp9q1tRYEg
1s/GJ0/5xopJ7Mja7KNwsxkeNyBmsObYUJ7+2r9/SGKqE+9syjvtUORT7zjCmhYjrje8dazGz3Ot
h5xlkgQsuelx7bXb650hJqkrU7jcZCs0YCMu7UzblO9yEeF/BLR1suxQ3k/YVXYeJs1BJxj9x9gg
Vp/1H7XvmbN0MncrprOIiwkSOXxXUwFdwoeHcqbfJ3Ks5R2ddyUbLF5Hd8W8h1f/81edc5IG63Zo
BMWjyMx6NpBufxxD5x2T+cCCbDFjuZkdkok4pJgds6Bmup6qrWnV4xISyyNGYzG1w4elv7Pq9x4C
6XRP+30yFtLKs+dHmXU549W1ny3kPpmnobdwCIhzCwrbhAkdC3D7ueVO7+77QYk5RvTzo18AAais
avY4TxVJqrxwAfSm/Rr9zPpgOSa/5YH6zZiUu0Ixr5a5hgf/mOW/yF/p4HRMMIw+HCtz3mIIR1Qf
OPLwXV8oRbNOe6coxQHfJbn+Yituw8THcrsG1tjnf3hTNVY6IopE0F2KveOXQLZMLEx8/MgTTFTR
nIJ938eHSh/GSH41cnfxxE7wCynQRg/Q024OniHVQrzuvBpe6f1nD5UF4EyVB8mT1v5XwzYBUmfl
YALg39IP38hmDSRfGWBOMAXuPjb2wIhMY9UKfdqU5ZsVa/eJNu2p2wUSg1Hj+Cx5ozwwKsk6IGLM
rfhSGEqai0jdWY0KIby9B4vbCXMMySpKohJn/kyseyTKZ29sayt1oKE6M0hm+NQTFwj2fbscJYKI
7D/q0SlBaEy34JD97FXZnmiwUJmtsf0p+hMAA0C57p54QK+Cx9DKYfdGQRL4MtMXXGSP4HN5AH9n
Gl+Cq/0SGjoam0ab4Djl5pgZC4y2BdYQm760+gWeBuNJGHqTSr7ANHLyB3UXN1sPaDk4mbfAa18z
S6pYpzZlruB7Bpxm28H+Sf2zQqYYnFM/y2Fa0LhXPoWPKofBisWsD+r0eG2vrgreoBwYQA9llVwN
NnOYgSZC3pt7mlmnZJdBcEVRbj8Bj0Q9Z9Xji/+mIVrAVXEmuMC/tyBQKv+dr5/cCq9c2QEazZvy
OUJ2Zgi3iju7iI8W9HNWmbADrI0WH7eoEPIj6r1p93QiUiKxmWLD3dpNzIxKSYYtqjt2ioY+qo7D
ZtwCOlb0HGt6bZtpNOzGcrc1jzSX4q2fFp9RJ1VoFIsGJg10C/DeJTg9RiXIE0WrNadXbrSDEitK
VFxQQvjPKu25on4MfdFGr4Y0+5x/XhXrcvKgDogr37vDoE58DL7RoHHNwhSNhYkK4+lt3VIyVoJu
fF5R7gbgsena7k6bL89tLyKCMDfDjMzgr9WLXr8W9r6fjwYuWAh6j+XrAfWcf7dQlweH2QRBSTVv
cjoSWqqLeAjEl05xvaE0knSI+6fdQb/VM8k00OMo7GcjraQm7dGgP2CU6NLAHHVuQxMsehy73T+9
iFw9mLLHTxg7wmplBFyHyyp0TDIYOeRVY7lNX6+GwtNaJOKwZtC2zgSXmjm/GHE6D9p1n5MEouhH
SPN5O/11Wmfs9iZDLh8ARuXNM33HONMGGJPgJfUrrshqhTkoEcR1eb1azUr8MBLBcKPFmP9AlANn
yQd4ouXh4IAh9SrDUY/V/dlz3+TMFe+iHIQ+k+m30o4e6KvODAywsllQYOq/EL2YUvQ7ta/hY+gv
ahXi3yNQGrkWnlle1dOZTWhusyphk56xhURdzLnZkhsNBZhFVBQPGFELTBJgVJwUGkv1cUFmgIuw
NzOMn4mny63gEYumFuPjwAjlRhZwbmoPYf1lYxwePYKggEzZwrLwgaMiuTbxq5a+OvLqAT9MbnOQ
QfHwyihhwst6sjApnRvhrhpj/x33IQpnXo4cabu1D+wDVNXU9jPTEF130ijdzOsI57HZlQ8Ev6Nj
uyu8u/MIlZKzmS+NlYberb2Ug9y1HbieO/DkddamEEG82i3f9WG1Oas2691T3EQ991zv9BYd9XKV
6Rp5lMdBwubLRywwhoi83OWtR7WkgLt+NaZLQSWNbEZfzz0QnMCP5e1yT/3ZiZbEyS+5jxmx2ZRK
9MxJMfr2E/5O6O34/aQ8fI8K6HgEZ+LGdIl0q4XzPVpxi9QWbGnzSTy7Ym6C1Um42qDELYR/Qj27
jfQOVTtjlFUko0klK+BjQXexvMubWClEbAEHNTaYgn/13zcRlQ/FJXzhIL6kfqlpyNrRzpNi05uV
6BX+Hbig3Rztv2+Np0UXpCinWvFwFB1hRxPVzl38XRfb+mdgkmxUyzQQG2YjBHEcintoqyLRE8rb
dXFLGJHMcwNmLRvMCCrh7jIz+v25FNTLK3oReX5gW2rCEIHT6QJE5LeJyeDXUMTkaQdk+9IIYYhT
xA2TGpt6LSsTRxFNGr5SoT9N3eF+bZJ2bOPPbI7mzWV97Yd39osp5DT/1W2GRDJWmKEDLEHLHFLa
ezrLN+49aoEJVEfcm/EukcjM+KGnpzo3IBLa/qv2O+UfkKU9LVJoD74JyK4e9b1WhJ54jypleG87
7wD9AnU2VMQWTbGgHhT1KQesCUuAceMjYh92Bjv9/i8DLavaJa2V8q5uwbDYJXKym1R81YGOMriT
IVsqD9vX6yRJENstcnd3eYkVAgG6Xce9OJxwDLhkUenxBFkyrRQFM13B/C3coKQ/3rclSFbha/lu
kUNgIMHxd04H4YsSPT7zImEwPUT6v49NEikz1riVNu7a2mZFBOI/wpkmxhG2KaiJIg3Ua+aMS5V2
gZ2TIjW7N1d5bPdckn+nNWgqIENK/tfDzAOx7PsdWoaYsHZBp9wxFjggYGjQFvkoCGF+cSBWZWFH
4lUzj0nVHEnPTryEC+wePhUO/r523q6hEHzqfZv4SQuJsgTiAMyQ7JaIDkRG3VfXA6F9ZKO70nyp
yB4OWAuflVgn/U6oZEiOEeDZVBzWZfFcYfZ9LMwsqGAk9Zci3I4fJJFnFqb547lyGLgo/6SNc+Tv
i1+AxM+2aaDGPXJKWdBOo6ShyL9LfWY+5PxCaPXUshcCV4namYb0vZW54Un9Ts9ffrmVzMur91oK
mI1u6C8KBk86+SfSdnHeg7Uw3WBsd1gwUNJVkDH/YB2JcdLZitlUqe3A626n6bn6XVbOhsxm9uET
q05KfZU226g+DiiDeg6PkkwObg4KZ5PPd0g7alJ/a3B+V9AHXg/28++8oFcCGQSTBSanm58haQOk
mLoBCsqnq7qFFvaF8GNKjO0Tq/g2kQyk/Zb4peSm9djd1MOaG/aGkb7hY2+kvyRQCeCCaZN9nYfu
IpEbd4yvj9O2dcjvaijq+9w0Pot3treL7JewLrkGWpG9yhAvDtP+OPw9cw12z60wC98F+ahXobvV
4xxONceTe1xt9eFZJe7d1v1QjPv2VfYy9c+oUDrABirJA0AR7Wok3YbcjrPCFoHv6N26NfczV9xe
4dYynlcW3j/RwM3nFBHQir2HJ4KOmjBxiUkwdLNBWmAsptyPinraoj4dKUeyn/yn1CcG+wUgeaaG
mqoBdiX+3nHEfXM3+R1pyPWWViKeriJaoexf43K4wEfEQ2lhubAkcn6n3OL+mPYgAm3ubFT9BxJG
uZYDuMgXXvNFF65U5CCtECDUko13gacVxvnF4UTEOPJtm8ncZbo8kfCkA4QlNAbTCy3q9fnRwHNR
Fwy8I+5cSCjjIdRxrlsQ86PPNgVsK+p2W4humPdDiGuRHWLCOlrQRQsPzcB0HWTrAaV9nCPjvHLn
qfnAqxcQTcB5ineZtqLrFAlzQJmRzcfJJyXISYZ1cmzFre0sT7URNRK1SYBM54kzK1Q0QXsw5iYK
DKUK70nPm0e6wrMQiLshoH8dJRRhOzKLsFDddXzj2pJBt8irFI7vaWduyTkMPmvutkQH9WHIya/v
RA+7jKMwVY+gPFWx2H2UvCyW0F/OoKa9FJ942y+CejwaBXsNdgXWhbYL2SKhor16tIR0ZKzs6C7y
lDvuZY0oeAwBBbQvM0y2v9g/Fl+mO7seC6BaY8Dv2ksOBoi5QhaqDSEnTuGgLjyoK4MqhjxzMXKL
kA6X7Gnjp2uDpc0QgqpNp6ikgCsIjqARpveAvKRrvejKcLt3LNTEPsIsHK1prIRLKxpK5dC8j8Q6
BOL7JbIwur72yBA+AUzPG4V0fWZaIveWXTVU+xG7gbWkEL23w2twY4rNEscYb7CCh5JTG6r0g8+F
F4n8JyHUdhpG0i9O1efDG+NlA1znPl/iBcq1aKDsrc6Kb3zcxcr9tRpSMFNAvzEz+jlwfUQxp9sE
Rm39lhEz7rd5xBE+cbf/6ukECmnkZLVaJCI2WwfTI54hnXmaIzK0cP2X9Bkw9r6XBHcgCVRWUrrz
7wMpASOXYk7EoIR8KWFqjS7Vtzf45brKaI/aQXnQTP7pwvPua3Gqbqi8pvJpFJ7ufyd2plzAp1Kg
pPeF2J0ryqmuOn0kHTnfDgKVmVT1up9bagxJulpQx57IYZfS6+Pyp46sGvMq2ofKGToQ4nStJ6U1
0FqT3BPlPqcDEHJBqVHiyapH5cmmrI5e7GNw2Vl3sF9gtCTl/kIbRLRuPgmZFxs/Hh98iCWs1hYy
LKd3MX3bJ5FCXSuSv4mlaf09pLhW1fMQXMeSq44GFfyOF+ldxErCOZ2dc07hxl4IJ+1tdy2ETjnt
ddV/sCNdJsvgNVSun0oCaRIfb+CSUZhfctZ2zP2py+QDtcYGNfZkAGYgS9CE+U9CfgPvI9qoSdFQ
TvH6L1M4F7QWazW9OIPPVoR9aaMbRlnovDSMBUcY7Q5kgHEnrG+M2fPlbVgWipO5QZl3KWennlT4
GKTYJUlXpf5EcG3UqTp/1rLNzHxxrHs/f0K9wEwIvW3jTiLJl3eGOVqhuvryML8U1ilCLg/YLuNB
8HSAM8RtUGSPtLTPOEh/R240TrNqGqzVkUjrTd+J6LQl+r/q4M+h4gPQHlnUr6T0SNAiW+eWeGX/
FfBFLe8JtkWOe7U3bARBEPwhmf1/F8MEWY0tSi8ArIA/h/u2ZKEztA0PdfI0zjWlrPQb5nY+2APw
JXRPelnKyOsU0FuTOUGMBuYgOQmhOeHnrC0MQcYtWcBhTHdCyJbXpnPkOs1ECqy3fCbyRJYHyrYg
HaC+SVOUje5Nc/sbKReo0mAFwVEa5vnN48bqx8Eb9zNRsgHmlQQgOQRtPPIkdHGVnZYeHOrI40nt
VCXgO5kAfbvM/b4p3wjM4ZP3PaHQdgyU1NXrjAVPbjFth9qNLgxJ1YH+rIm9JWJKtSngQFDESwfQ
wQSRjNIE7WpPiYoMHDKu9yvIdqDLVmhzEKlwr+9As+T5JHaeHEDRl54TL8hyw3DFL2uoPtYHm/8u
op00g+f3skRcb9+sTAjpOqrynZ5dSQmRrD7qQDKoWfB0FkJ3BhMdl3dqGKF0buGs5y8AI0olxEhs
ILtd3C/8/nwv6h57RUq5rRDiFfsw9V0QS2yKkbq8quCOJ4jFjp+tE2+kd72hMJfqu3myqx5rQZeg
6Nv+EE8LHQpKkTr3hAJJCBSjVPJJ3h+aOUNHzoXUgBhZljW2j68W59GGFR7pTdKKA819qz0iTweh
yroCsBkLrAIYl4OkFrEMGE9Jg96B3WilrCCa2QlnQw+akz2j7tfRofOdPBJ/yIRBeA4+GE5Qe9+X
wgKXuLe9yhVl4Bn9lAPUJ47SCdLWSsZZFzh4cY3Og0eDThwQaK/oOjhjPZdrvI0pbk/v1ojmyFrN
Sc7Z40B3pLV02qgAtXOCdoX3PzVQnOIrH9CKL52GVGZRLo5oiXG+VLio02TkMUSrk4PpE61IPw8K
DB6OX3gU99nrDkBTjqQE4zRUGv7QtD+aARd7Ahkoybp3LWqYRYQOYzLzz/QtpLKKJEZtoTwFb6Ab
jieN1GVjIQjSNit2LmfQPNaq2TwTtmzHkf3lujlP9rNBeY7bJZS06FjMyDmBIHrvvf39/dWlYmOz
YaBDwJwsB35WowlVqfJH+B6pL71vndMmN7qbrBAwEPmAd8YNr/lvVue0iZXcKP6S7KjtqJL/VdD4
S1TyHUOJE0esDpGkd4Mi+wZUdz2Wlnw0b+K/LYH6DekQlhKxBwUV0cMgc4dpkkjNPPFQghYI0zUZ
I/kcuKGnXc31LZxfzsu/u9n5cuBq9VXg9x59OSZWuOhHfgYRmJdkBOz1rO0uBT2pLKHvFAXwVOWz
/xvS4gWF7RrPPfiIi3M54gWmXceWdvGx3SRIjGHgV0Cb17xUcw+5HuQtC5uQAwNfBI1nX/c5++Y7
s7ATxSOif7uELVfp1+zxCIviAuHFl2oLb+8VUEhLTJZ5wN5Uore6JYEhxpz+WRlg40PJS1OF2z69
tLb+PAqEjnAUCYHch71bipW3+6L9MWp+gJYR+flYxnqTgExBN47GypiGAkvsdFxgeL3OkakyF8w1
czM3A4XJrYqqfe8K+GCkCXayG/FqChdKjtu7UEMK29PUahlKk3imuCqZYy1BhrAs1ZbI7W68I4sk
FnJNtbg8hiKZ2ScxRzAF+Oji0E173K0uPC8lDZbA87lvxz3yOTKXtcYMjUjHwLE5ZBQ53MnbSaAR
XBJsrrixPrNJ+LuoTigG3FzaaGr+T1cCGni21lVWd9Blr9/eikFlhAxUpgEMeoZqwxoBm4ZdBz20
evHL6PbAm1U6ATQXjd2d9ZNa4c9XXaR0d23MvVnukIl42VcaW1b40MoBAE0U+i3NPbwNRXzyjS5u
ZvX+twrwkwgNBBqyZhDM8Va9zZuP84v0myiarTzo7vKn6mQoYA81TOxfNy4QOodhEQfoGDboVBXI
SNHTCACpg38njZzg1HKmtpxgm3Nk68oV9hP8TLur23zPT0UIzujFQ+tDH5+glas/zdZCwas9I2k5
zQueIXPZP8n0IORR+1GvQceiHooGDFMWLTUqXnBxOtduXuMbgtw/dbTbTlePlLUvG5n9ts2/P/W/
XiUpwy+vFBDaEG6U0PJAcxSAMkIMn8M9X5tDjGIsDZTRqJjmKrcQnKVWJya9+XITIh6qKdPzibVZ
3OY7wN7JLKE3ChMuk6VoGHFUDFvinyrg9902V8LsmcAtl1lkagBfkq5tSY0ZmEwwlB0CRIwpQ6X9
5kX8vK+5fIVI8zsT8MziGscfzzHpYR18ccVwEf6zT/OMvzMSwP4BphoM0h1RqicD4WbI2IDiKMsY
ue/WP25qqgMgvfgxB3zn8uq5g+CWTSJHFJsGdMVJFX10DU6Qy255fJ00kDSXuSuqnAWIhj97vdpu
83lWIikgNjDJ7Pl9vtJQmHgllnqYL2BpxUqZsrlDvQo/jZ7GL9iA2WWvhjvJfhn4xG7atGrif74J
b+JwdG4EavjGJdGR+aC9tftt4dCLv+IZmKR/S/LqWAtuWRTVOoSU5piNXXA91FvIlDerJFNa4Krh
qc4oYaqdtWNv4hzGqNROzbYGu8lowjmjrHq68t128xLZN3S/wJF3EXeJ0E2mU72Fqi46UEbD2Xy5
dpyKWMZQnXLJ2vuoQK2vvO4j9iJZnRYpxI9NGaqFE+CLvEp/ATmc0T+KL+mdcTve6V/N5xsqWp3P
GU46jJk28KrahHUHVf1GUTCCt3HFGU1madJ64zxAN+N15LajOr0963Z83PjRrDLjzjlmglSp/gzH
luP7HeS44ylpIv1lqCs8O4EdPSCM2JF9ug8SBa+7ofj9P5TzFeZjaEXHbTUWVTvKk9/MPw5TaIqJ
8KVyruaNiIuFcX0Q17eBJym5d/OK+1AHcj0ia17LbMW/jfD0WfxktukvbrfpYOfC2Cy+FlkuoHZG
fGRmpxuUJspdfAcYyDAgCU6Htg7vvPQF64fnsyi7dKfE5WMlyDBbmBhqV9camZQksNgE5K+mHJ+3
1p+Th79JaM4cSfk4Hu/Wsi1o+K9SncT8trgcm8WFG9UoYNLyZX7LlAdk7CzAzxTsW4/9BNiFXdCd
BxB6aU7NToou9pxxFlydpSReNn3ih+qA4rTK7ctXOfgF+YuQIOWzaN471jY4pkFC1KXWBcPmtHjP
98ZGT2HA8mpaVxtVRythPjuV0YAV7pSFXNBlcc98TCTXCfOii60UKyA6t7mQ/apLGAoFAwIiLLrq
8pNu+O1xpFPf+emhDg5NLX8ltz8g4TncB9HHRm+NPzjPz8yKcELJqI/Gp+85eX2SwAYlqaSYWg3a
KZtB8Dgow7kczqHTu3zgXkejBb2zlW02fZ/WR4p8LGL+ltI2pbAFZbnrwcDsCXGocXLe97gi+g88
u04Q/NzTfNiQBUAZ1Qh4/dKrq6bqwZJDr2Bg29744CheEpLx5xdgAr2L26CuNN4Yu5z/41lwRmHF
eMT5RyCYNAj1VRj81nmjiyHsZlxwj3QG8SwNe6ZBIKpRARGgxnFnEWdKkG+O5ILo4X71WrQFBXTF
uwQKvItIbaUeQMuFjGkmCIKiZ55NpORKerFjY8BwblzjfMGleSp9Es2KmMrI20iAmm+BI+zpVFYf
n6mOlhUT17NgVwWZdRpGsWfxUmYPxz814y2oxvKJhKb6U45H5N/H38e4CBtSm0g4g3YhTej8amZF
WKtRUHBno6QvMq/13ONChEU2++o1PD64y/a22FdhZ3cSVbZlXtWVbhyXARrGU+zWZfkABAJCmsRQ
5jXM/0eNKF3pqtDzGqrVrYdcYCTer0wBgKgP6bKe4lc0WC6ofcwPqyfxTEpiPbz32Ag08K0lRp24
bhloriZFyRe/CGRa11lpRT5GgQJDkTGFFH6n+GRvg0J6x8Yob8EEIofNooCYUtQh/WPmX0Lfdjp7
agfm7LV5HxsGp9eB7W3WHHVSY/1W2Ud6zfZz4ZZYNRVoV0ef1pmGx8fTV6vjR6KjXO+s7DHInuPQ
eYDfIZLNtBPziL5sWXlmPmjUccvWATTWUjhUFpeBpPhYkXNvBiqUtJpa2r4nwp14PjA5G6+g5/C6
Ur1JAkR3Xez0LNfhvXQ/DlAz+u364L6ur02KHOgAJeny4iMo9Tb1mqreaWrAZZhwUg5OHETYDph8
X3ondj4qGdYbvQKpoDRgWexa5xLoxqvYL5diYZOkKifX+dt/E8ESA8SfJo6ZwOyMawu4ILBGW/t9
mI8DESx7jvzPwdeluKwup8Ku99k4es8sDi443wb+kVGgCihleMkBeFyQcPOEpNkE7i+80wQ6YPk1
6REMKmJ2Qhy7SGP6SiSjnDhUZs1nSAFDdFmbagxbWLnL+ldgfMfB4Arv7SJxbNmdgPsvwhrZYzyz
WgWyuUHnVFTm1+DZGGnVoUNHmhPhlvcZXMrfPstPNnWd5zpUIQGQWi+M+4jeibx19CE2BBrdKDtf
dnIBbLwC/ACePoo5wPWRbNROffXTrGMLSvXIq6mozWIAtxcaNWq5I8USwesxC/CnM2cvj9DeC1qg
iwZlAcb1MhXnjI/nBGA4ww9uaHXaGTZN0wSiiNrgyOK0r041aos80ctSPLAWRTlwwXqA90j3I5yK
BeHDPq9XTO/bD/aGAsywcewf5fQEj2KCAws6dFrvJrB5KziaI/oo7HJCeIXaSvDAn/6UlIpktqcJ
3RmEUUM8HPQ665BUbTqD+2MlUO7f9m9Uypy+VNqFjToWB1l7AvRrkNUzUr+BbqCtbJaThC1F5ckN
hRcUzGWj9fCfgXtOLCJWtzGDQ+cZQLAAvQA17MLbMtP5UuW3MQayawe5SBZSl6wjqGIRDvjUraq+
p7q05U9wSzPIVlAwFHJrMdkrpUPUVaPi6OiCoZZdfAEeGPlKLlHqP/En21TqROPxHoWeHWP0Qonl
JINEFI/xcVO9zG/vPxyPKhJlpD/57s5g9WmJFvVaXaCPo7+zHxYVRbxuDsMBXgDVPsxhGpmirlKv
W/xKOB5kLw2M8szbHrKhlMZwUwhrnqRG2fK0JiaGwOBDoNigzSo7PE57xQSfRmcaD9Lao+wG4M1N
60r6oL7FEBWyhu9go2mJFu+NFOHFkPkNSASiZny0DnDl5mKkmhuWDAKJNxyGiGiKrClf0bV/GbzJ
SGhlaEtZMFre0oq2dpGa0pThhgy0yx6mG0+th9xCVc1hSWUxhnDKQZwjfX4D7J756zIdhWfkgAgN
pQfdT2b157xEw/NXC6dvO7aS6dJJ6T8FCvpVwByoCRSG26L7lSh7VFRJ1UfOkE8hIgcWzCdtIowo
AS+7pfF34IoMniy34GAjV5abCC4OODq+Wpid672/bzoI3LPDWGl9gJoiZcWz38bE4xn2EgQPNSex
QXVzVkQ5+qEC1l/K3jSM+9UHEsM6+Rj3xgfDYiXSB+5ejSDUJEwApNDzuHnkWD6eJO/GJz/NStmz
6/lIyc4CkjEtgVBGsRyFawzle4M+bBSdWHYch2J3gBAVzbRZnCw1rD70L1O4oV7YJaKpZIKZvBQH
YdtwHIxVusuCRKtvVIfqk6lf8NxO02c+wi9L9ug9uy025Y8cYaxiFblFGhTIjoefw3oKsl+9F/di
NsuCZnSwqW6pwsU0dzsEY3bEHuVmmnx0pXgfuBL1yXK0PV3016K13dSVkW5hDgeVp0zO/yLgC5gt
NmZb48To75UCfPu5XBWMeCZO5AFdqVQNCprVP5L1HGRQbjBFtcV8lLRdlNnMEBZDfDw6gTL5BwcI
Pb/uW/eKYhvoRKFW4+Xwdqs3h1M1UaMN5J+pl8L5gHHhMiNAcIPcwFXPYARFb6QyQIGQQofdpMdt
9zlVYjhnBZ/IPvSGCluFkzkTTKsT9bXnmzJkksSBxz2yZ0Uac01CwloChFEB/e/zI+0eVhRmk/o4
WQDu60GG+Ho7Xocn8KAtQvF49e9pvam5V1sTLFm76fsDvVZ0EmbPBZ1rjRWkA04ugdICUHvWbIIn
zMugNXEwk9Fcx7qYjkEUVR7Q+QfZScjWUP3DjZFRQc+M8bB3/miiuswcH809HBfR7gDD/l/M8ktC
3c9ujTzJXYFYHrtmmyVyrsgEODmEyzpSg5UPJaoMhyIDRYHMCFded3+9dHmtvmmknEkZPBDiEbQY
E1vC0o2Prni0dDj4qFnU7UAw2e5c4BAODi1+nbslrB+MEc8Pvp+S9unejYPvFn4QnlH09KZsoKsB
mZKe0u2o9cbliyB3fPacUnz6tvyFdJVauMVnSrDN6N4S7JrYrAxDE7rjQGIoqb8bkhB7GPlRLX24
TP9RzG+XvJFSNGl1ca7NHTAaufRCel3qtmRaQmClzJ+GNtD30iOmmnZQEtxXt09cvgvVnm9aD8su
KO1iEHLvN8sTSJ+0OoY/jscIOJoK6eCGmYizMMeT4Reg7fCPENKO4d5VTklIJSWEwIRgohQ0378+
tuZLb8FnQ0ejnj0yLOrgb4xFeSrqR9MKkRZn05lLk7yYaV+o6NDDec7Cpw4BKF+VN8+m01oXx+B3
6vLvqd43i9gOenKZBh2gmqCZg0GGwLSRNWpGIPOAoka4TID+RN4SIBGwoUnPysXgORpx6jSIAvNW
FoBI1x7tCEDa2EdS+Ty9xtK8XeeC/9paUGa4dmuf62N91Tdo2PGTz5o+YabfrHin6uu7MzWKujw2
sX9PNO/9R9iNZuVBuw5VnoxwKmZaAwBArU4SA8Lz088eN9rbkmXAC30Hjdiu7yH0RFdaqA/TLfgP
HZDJB9FnB49+OVYxERcqDs6gCI/hkPYty3h67B4+VG6XuV48Ahv4XFmxVZtWpy0AJYr3a3pdgUxD
wdUttqeFOVili9VFTk1dm2bRtLcX74x8YttrtCAuzfq7SjyvvVsbN0/WFs80UN3dI4qAfAtp3zeh
pNhcrJcpVmK/sQmU9S7JCm996jJSohYey6bUBKspryoqJvrvOXf7C7yWfMokxpAdiRtpR6VVvt2E
jznd2JuaGkKa+nywyt3wlfkTs3AbOrJHywTLkLRdVv/tk9yeZ5/cNgCxZdQ+muWeVi9sRUggGscP
iZoE9D2O/cD7LQN51Jl1bn8xjTVGR8Z1oFQxs45QKIp7Jdc3qN9yyj3GhLtgMbaiaL2DOrbxe4W0
LGgQ1TISj4rbp2TIQ4BMT+fU2MPXxmPz8RPnb+7GCQt6DN80GNYHBVN0X5F9LdPVHW0t8lzutoD8
QzjAtut6p2od6JCaRB5Jgui/Uu7/eVeYtWnKSB9WOiBqXH6ONPw+oOUYkpPLIFn8+/jSlChYOfKa
NbKyOVXWgPQnC5nUrNrLWjsnjE5JVatl7XcrFMUrJTSzXCgUBcoGCDC8Fd+cdZt+tEIX5xt4QHlZ
3VRybqE90N0GOPKfxJw1F+dCA/H0OwIm4kfsMqhEalpJ6PFj43C3Bul9wfM2Y9H4yrx+DE2b0pAz
u26rSyAADvTPvdXq64NCuf8OMR0U7PEETuX84etpsl9fwGr32cEff/VcZ95QPzJWBtVkeBQSFVjf
RBHtr2Eqe89lDHvfcXKAiooARZTI1Wq6OjyO0jg1rIUL2QEUr740wLKLjym2bxYyxMPz0NIuTEv7
8I9z6V4cHjx+pPkUnkIDgiEEEraNGh3y8b+Nrs+l+L8B+Y5bONl0EI/nF3TrmgzL28A+lQ4bwMQa
46vWS9cno6rV9nRvvqxeQ7Zsz+vsFRuz6+qdEb/DYEK6AeO198DbdHRrkl9mB03NTFWSgkoqOIBZ
AN0e6rzIm0AD3t/mZ3qByd5kUoauJ0JmhwVy2Lulaj4yk7AlApLQWcimN/xbqUNFL+9psRBKNrRP
6QLEqHQ5OFUT09D0JWQTYTJ04CzHx1QAGjS5ogz0yGKQirXnl4dZknVRw3OrMKaDz1NwxhEoqtM7
ukqn5u0GGp0h6PchkJb8gyZxoJpl2qkhwLr97k2bm+aTfOSu4AJg98hSXiajbJsJUy7t+uXyAt+G
qliwfbt6ghC2Gi7YZf2o5XPuaR5o/kXnJkst4aAaTrM+nt6OEBIEU77mJKMN4bneW3meCpjbRxHN
xqlRp9ID11WVrNSMS6Ej8/Yd17TaEUUnVmG6QCBKvwgsgDsta4mvQILmU2ylYN/hfCjEtnLLFzmr
6aJVbqbKDyklKG/eRqVQsPX9bfEL6RlYUP99vxJjpcPIti8nK7lXor9tqXZqcrXUeW5t5GHerM0g
1DRgRx1lhY/tTITyFqXR1kr16DgAXnrKgm0MhhBYTdnhFgPSf2nuShr5tLyYtbc8Za/ykSNRyiZk
U/QEZdFWFAm972YOqx/RniBGRWPZEiOiZZCIEMNsEwrF65RsuBz8fMBvJch6lYbmVbtFi+R9LFp9
3yXwlCz9DPrVTA/zhYY97NZO+uZkpp9YbIvD344JB0w7kZALBxMKiM8VS1w3o2HfVFCuTgKsXrpS
4dJGeUKoCcBhSOqNEj5iSM3KvUEx0Bf5q1H/3Vdqd/Q2MkFLtVDaWqXSB6S38VCv0dkDevPsLXOy
aMCszLhJFg3Na7oDp2djV/cRM2YjOVuugJ7QCZjkpCfA2rfd/Okp9PZXedFRUmqNH/zSthk4Oqid
KwKnASTH32rmWTnYHRwFPYMydud09IA2FVVkul8NSNi6wn+EIu5wLJGwBuROV9AI9++e5N0lp+3q
eVdbyQmabZk/ihWSORxtY6ow/OyWpxAHS6HUv5LgZVR5lKVW4zElZMAfv/sVFD3vBW2JNz07KrlD
7/JPGCNBZ+mv/IcD1kjpisQQoXRdgR1fdqc2zdFDuP9WU/XDUwPGLY4FSdc9LffAgo9d4IH8rI+o
o+bHyJrescvKOpKYrMcYNzDLgDxF+pO8IovhDdZG5Mvwn4VU7NmVyqiNqmCzPAwbnDd5xs8wuDA9
/NkNxKdNbBqTgjVAMsN2fxzLmvijxWmtRhpLRVDj01Kv5U+Me4BV/YtrkLavd2rBYsnFfWoUm4pa
DLt393tw4VVO76eMxagfTfHLVSq/ewkhswihToCfe44g7AeZFrIy4/HWZ0AEbrVlBSY0vFFuLJy4
HKE2U43TG64/NClQYZiI584sWJnwoKGooGifIX8OEnVtYQZHNO6JjlP8snRcYAj3ecDWyhL7CUgR
P/hAmZmSguuVxUZ8M0h1LQYs5CeSr5r5SaAr6xX8iNjLnVsi8VuCs21lxhqvOZ4pysanoWmoF3wG
BT1Z+Uq2EB9gdbKvAIg1k2EWmMSG1Taoucyp9373Lrt99EUg02hpaK2hPCeZRmMxmSvHXOCC3UZa
RfYgZB3POs4pdrhz/PfE+H9DmkuB+wcvFTGqN13hZrcZD2+XHVe1HJYH/jyR7yZal2w+vMQQYZkG
4kAIdqn5enYO5PPO9kJZk6JnGmWwpDgbcQuBjUvMSq4nR1ae+hFuM+x90+vjFUPdqpk55z7wLZUj
YX6fD/cSh41DdVG78nuJrNW9MLbDlHF3aXbjoaH57+OxB9iDxFpwW3H8qukqCE9dlqhM+KJHDVgL
8liiKf/Yn3CyH8QG+eOvy4KUfxRrw/VQe7n3IRI0qPyCpGoZ67d6Pf/6qCt4SsajxkhR3JfCrLil
cbJAdfbFL0mES2z4UNikcDsit75ad55krYORt82QXJBzS1tkTZ8ajgq+ghPrp+VZD8q178Eprl4D
TzQxng6dze3c/7ysJDKCiQY2UJHOQ55V7gKt9R7yTBBHLhEOUqIJBh/0jYPny7iEvyxrGVUj8qYC
BBoOcJ9lHeB1Eb4Vttqj2IBMZ5ODddertDWFaQOfdlBj5mh3OLkyngNqfg+QWenh9QuXHNbHn5oK
3bRzKznVmnoX62Ec2areuEnEomfJYSSoSmtQt9X3SjAoWnzfxsXkTfSuW9lW4Zq3ERN369DIRX9O
2bGm3hpeQnnJip0vEK6fkqwB99rLmdf9c3RqUzE79G3sSv69CYfGMn5dOsw/+P/gO31rdEDJV3mH
P+3UJKOEVu+ZDG/TqCn+TDllJVh7vrHKqx7xdndr4oDbfoorOVGR9XSwbMPG14f8wZXLvxwIwXBt
h8y1MpCw7XA0WGJc0SH7vH0ecuYJbEzrZhzOFoYeFWymOtmZARau10KFNTsZ4w68aDUcQXwxPBtR
aSGOgTUYgMGbCz2qDgeWCJ4ONXcsuIwjyZTSwOpK31yRoiH3aoQooAR1CbcoVVaP186CXyaaHa0C
OYmKbYnhN8kb+JNsvkHE3GpREWKcVo9rPepfYV+7fRRDpHU9ODB8hiN945uGYIQhsRxitql0/KKk
WUzEq8+6KbAe8m6G57Ft/q+gAWad5jZZvEvuEIPEtOerzFTWriK3EMeLz5K1cKCcLiB1K2x5CS3I
uXYD1F6COgv0GEeM9unCmGoo6cqQx0+pSZNhY3WhAi//KbwPI5AtXPntPwE/OMPQ7Hp1rVSKuTcT
en6T30QpifwIhypKAp2aoyZU22+33o1GuiIq03hoW/T0XVKHw/IJEGmbe7c/BICN6E69qcRWqvXf
keHpwN6idI0tegy+ZLpR9h7VDW3FSw0rSQoTF6IX2DctPKfY4B6zC/1A2v0Othe9/ciwpnBtcY6k
thU94wIxK5R9NtjY9A/xKvPQzFeZBlmB5lkacLJ96GKpYkFX7bp2FQtvyDqLTNqWvAzPx5USDA1N
O60ZT5gN/bejmLN/ULs1LyAIeTSGdjfXIfA4hLgtCIS08VLr2er01N+7q7/TGjQCliuZvbKPWKt+
W2a7XhryFTd+b6DSenSrVPxddVRz5Y7vAucYFz2Cs/42Dth7LBgFXmIbfY+O2qLXrPEpXbBX8XEW
lR6YiMkmr3UdGeIYyPAQcIiG9FoHd+fJEDk934y3MlewSftI4XCKl4cmjZejpLK3fi25ethnEhgI
m0x8SnrXF62VIK0jP8I5WPQ887yGeq5JiwrfoypKYQ+22VBpG7pI2XgsFPEl3yeZbqa3vqGoQKnH
lxAMBH1kt+1058uKhe7TwFlFkgFgV7r5viSpKkeTe8Zbu8sSlBfWbQWaZKEqjWCJFz8iKWNfviil
RLIrcBpZxMR9JvHXAvrI+xVCjeJXLY4ipIvVDyHcaVIcGx9F6cUO1lp9gd9FK1TCtE8+M5OkEOUF
Q4f/e2n18fR34gwTKsH8WUd8UqJRERmeer0OEPmFf5QU8iU1wXZSahneqgnzhgbAzFDAqJ3pg0cK
CsImps8kluts5qQ6CUVyPrZxY0CtaP/eTNjDzQ6Wxr7nyYoTEuuKNM3e1SGBnGifgYBhkBTtRy/m
454rVp8wjISZVc2ohWqtmPN07wZij4K73/Wgtwc5AZ4XMCYDcXN/O96KrVQLxL7IT63S2zJ4FDoe
feQ3+Z/9m/N6zEKwDwrHXAo62cgGciJzuzpGv2ATSuFDWeexT9D2GhfT0IKMJRH+AqgaLQUG1SnT
xM6kpmvgWo3HmXTZNT41PrI57piq2W+8TpWdwtrqjUh1AV8SeYR7b0/rbBHX29f04ACdbuaBKUmp
FvVW0ME3ZPQEegRphZ/MwDF/s+JEAIkS8lsxCC6Od5NYkDhkmQDS1z7kneDUZb3aoVki7IUhHvkG
kqs0Q62ifVkJPKpzLeMhELRL8t7o7QujlUjIKNHtK+drvi4FkEJgZrQnQEltoLStHmTe9goaQwiJ
ArtV3/oJ08rV34wy3Br5uy9i0pNGNvgx/YzSU6xv2W6sRad3jiF1visBvCBAQhps/Kvlutfx7JxW
vQee47gshkvZFu+5YB98LOFBsG+0I3J931q0yen+7zwSgisv9HRBcQnq+ENgTn8oBgPU8GNcdkNq
6AasiQuni62/sOeThtqNPmZZUwX/pL9aTLpE+IvqGVCJpgQsREGxUlT+Svd8UZq98xWYntv3pOHF
+U9s6SLU+CmI3sz2uw7T8VdoM4Q+8kkPHEMOuiJxynPSpl/+vjXvr1biDYu+fsQiECMx/okTmzpw
VDaUBzczlCOIxjtqzyrVGrrUNk4SWEsGdhwcQ0+vRjDDfXi83S+/OKqZu4f0smodtEkO65eADQxd
f71ClYf81xsGCqNUI825DidvqEyf5Knr18eroQ64S1E3eEBE3bVMzrCTyMylyB7kOMpGGcEAFD4X
dZO21219ip9Cnk4z4MfFUfKiCRH8Aa3tAiDHhq2C8K51eTTRC1Kyq3zMRH8XTd4UsQNXKWMXWj3g
sJ+At6d0b/jUzz2B6uf9cYcunMEIs1Nd6NQ8lom7TjasPXNVV7TiE8JAygBHxoTLhvkYDAeCYw8z
BjEjPxiectmnClHRRpWbOOCyxyqTFaFqeefb81SRhQ6IkWhLoT3xwTOPetEWcbyhttatfYEXYQBb
hPbTmF8CqbuZYlrmMzvfmZ3zqtORDBf1AZsWgrjv5ZgLs5NsPq3rfg6LoduOQLZuNDIgHZsmNaHf
mVzrj8D2+8fC4kkq1WJUtFgtr2BREwuGlTqTQc266Le0r+AJREbF7B9f1oz98HjoWMxUKlsxEyT8
L3G+42GUgIWvcR5WmVsOOXzTPhwwtL2WV55/C6LWFLJHtAAsnUrsipT1Hx4X6EUs/h472y9PNmNI
7yH1OMDDrcUgXoT/NNjfhcetoRZ3FbsiSTUKPR00SN3e5cI+uvZ64j+zdT0dwDig+mnX2xXeYi+v
NlsgIyAQbTLsFX9NCUcTqHITbzNO4hWKkBV7250wutjADU3PSrlQx51ioNDBlICR+7RlHz3pXWHO
5LlLW5iY3Wa1bsgJ3PzbWHwcHhp+oQyIiq6GH+VhYulSmJ4wPEll3ZJe8qDpz/d0cCVMfgtYUFlo
7e82yiIuP47CKmOPQFzvefKC4nDNie2GqappIDprv9eusFG4mdSW6U09dg/NGBaSBdAtYRVa1h5E
u+vNubUKOvuPeQ+YjATw70optrL7ZNu5/2NctyPjvzHoBz/kW3PDLC9zkPWYRFharCjtyTPqdY/g
ZtndO7UwuATDCqMPeO2S2cLcz/VYgQ2A14d3O7UAWkOzDIG2dZOG6CU3iDAcPjHatZKzGmk03tra
NZvAQx5V6RToqKYm66oYYvKMLyeXeGghwb8oi9kWQ+Q51izzPcUwT4gmWqYcfMp1Q6FUgkxQ/d0h
lKxyYSxSyPjJ1wdQhzMBDwd9q4kc5+syPmJBUWVtWflLxC2sGahcgx9CPtuau4IdzBHPY1DEOxL5
zbLfZcyJ52CP5iGRL0T4QjvvSQAfcbPX/kkEW+m7DxPhHKKFzBEvaVW6lwHDsM1EhhULOb3gdw6z
LVFVk7pqrf35njcL+UGPf5fZ6ntDjMMHlPp60nSPfwfL31sQqk6fgvltZ0uxdtT6HlzACieVTEmE
mYzU9NYoZlWwMiVx8iK59elui8ChPxXdf+42BRMruclYWZoaflPHs7CP9idTN1djekMZElNIoosK
O0cwey/KZbS+fmix6iJdv3zBWTlhY4IVZleXpY4pgheBaR+scnjop4kfJHaIrNg1U20bjxb2CR+C
t7bgUW32RHCzO9plNghBjvQoVEgLi90RAX3+qrJjFaYv29hsIqukKMGToKhz5j9ptQ1ygwApBDLp
O6dI0g/Sno/aRH89RNFQjrPvW+plFn6PlYOZwJPwlwvZuLxm7dkMlvJ9OHHDn7R1bKY9ZE/4YsLy
7FIkYKNp71cnrC6UaY4YMuPViNZzPWhteXdI/pObeFqLM73FWea4GHuD2y5Pu0zT/077Ip8RpFXJ
JnA/wF+mQdTNDaRv6om8YlwV76Api/EmLvEUT3Uv+HV5X6SGa8uYTkBzVAi74ocFuZndfRZhJaER
tG0h63Gl/NNfTWqHemhPHER3bZd/YeH0TT4U7JnhIJEChwkoUjN7TnlnWnjlEiN7tKlfF3Mj+UXq
ma8KCsCyKxnIdZK2akF+ydyXkqs3FxaZjUu54Bgw/0EWQa6SYrEFT8sPBdfGpUlDZm92XoMQfrxe
DCgJ85JTRu37af4iCeDaTCLZSYz/zOpJlIjp6F9LKd6mU7tVoNMMr6PYPDdqYxiQmWz7mrogBZWW
fTsENuGiT+41C9BQt+nULpT6ihSoIT00UN+rCAjgUGDoRjDLsMaOjerMTiOwgS1Y0ruIY5WP2vqO
JhL1+ch6c6SV/TcduQIbsKJAkykE0dquSEvhlhjk3U1qIxgDYoG255C8AdsdJHKx+ZDH1KM6hTjY
iFcK1vsmYZrhj+QM937rKvIQd5ywsXUrVGdIzy7uI0AAj3/7JH14Y3WeYrhiE3EpZM8MELa9sG0K
4UzzxrVGwnkOc8org1qvOECcfhCd+S9yVITME+eLlJLUIFBhdGiH4R209oXq9TVFI+glEbO2Nx/H
Zu4PuatnXq1IvZu3BVqBA7jtvDDAUFB3EnBFjzKdmYat00IS4yeK7JjsDMrqWvi9TP7GMOncWmBm
lawGu8exCkJ95mvkZJfQv8Fvj9p2oio2Et2bijNjo+n3++X0oZV/a6BA1Ptc+9c/PMV/+o59LLR6
66d0kZRDz2850flqn23j7uFc4kmRF0ZWNrFRzTcVIob+ThVeZL2U7FJexE2gRKBMAKgtJYcTAWyV
rw0TyWCitTnJ3ZlDxaZK+pxzysD0bgSrdfdyAjBmRIeJSe3eq66NmcGwVAom/J+0ig+zHBpwRwy6
ocYaN7aA3QgDtr5RCU8reiZYAWEcPP3ctSmbNmV+yGnF4fBuxqyUcTiGmtM4rF60Tua3tE6/KBVG
kNNr1+Idt+cxoJqcB5a875m5pXwY39Qy0ITNTmSwPKQhVLHowdvNcfjQMn0ZrCaHfZgYvJqR3uw6
eH7z/yyCxAncWTixUlov/3YE02iBeDy5eb9xMak6Flk1poRm2r3fEAOyD+pTx/QQKQTNH3pdB7dv
RBCKMKBeABnCX5AWO4yHTx+kRX2CwpnrTObdQ2PYwBmkIimGh4q61NBFXkN5dbjbuwDoVY+7Kqe/
cN7a50bvAoieEqm9/qFU/4TH07rxzor4haioYB89Mh1uUDHHhsN6Wcwon2iyQjQAyWaVQ00xCROS
QjXQP37pkVNDv1gOe70aYw3MzBnmp9ZCLzg2/adzdrU2zGuQI3ERUJsMTMbnQSAK4By7/bnMkC2i
+5w/MC7lFsytcmuEeW3nFCU3S0MaD0YvVyQ93/MqgkAD5yw5PW0QLoJlfYGa9Y8VHEmuMhJKo5dW
khaIylW1ZnBYW+ZGza+tH3SE3MWyoRAN+S0uXDwvIGx+uZ9LRHV+1OZ+HtxUWRn+rtQOy119JttY
jTX/BYsA9RJzOwEgjKgKw+C0oYPj5oOeo0FSO2q+dDW3ESaMRfuUxkwvYRSnUnMSWMkMi12Pcdyb
pzOWNKAc6dsHtfCnRka+77cBPJdhRXfVy7e5GNEt73Fc4AUSv6aOttMfnmxuN3inU0jOa45RX8Ts
35TICh0lVaPKnXqSUs+K/dljE6ECmpDZtJzFvs8jLPzqE+3ouAuTfbcdbaA+NqRKhUra3rW/ENlo
GEfqQQDIbMbnH00gCOmjzxbDfS7PfuaaLK/2rPctYEwhm4syTTyw6WPeWn7qytpamfD94ApzrDwW
l0/i9bM+7zQimxtFTg592pdAwMbvzS8Mua8tA6xhf/7bAaQd1MbLfspWqkIpES4mz7mQslmWrWQ4
tFVoCXlfnJ52Q1BBvR6+zifOn8dr/IOccyw3GIxuyQQFmAr4lIfxMGYZwvKDbwqu2Zxb6dgrzdVX
fLDpQp7/4mzt8vdc2qNra9ounz4SHujORI1LK8SzN80cr1B3i6oCRvDG9DM4OilTq3no/f+v0rAV
R5909nhwT2b+N6FzWo86efC/gal4jv4b3KUBUTumIVrJnDG7sIvKF3Gns81hXWXuWqgLVglBu58F
VnJt8jP4XBy0qbpdPHPEIi621yHDpI+iMrucxi5ovUGeOjNK574zyhjJHwdi+Ud0bcejzI5KruNI
3Nc53rPuaxKxs0k8VMv3Bi2pLAHC+aUFBB0mvI3wFZpr2emGV66RHiMBQPfL97/IEWOCBXbJmk0P
F4sWyBdmtWxZ7Abslj4k7+DzjdLYS63j8NavP5EDz35Q2iGRMhZPR84QFtRtvjwIzVbGzsD+y7tq
81RfkGuNnS3/2ytVPptVY3u6/Ke7FH5BCEBd7FnUQ4iEsjl/3ce9JjTX/H+fxJT9BxvK6ZwdPAgV
T7tc1f0DQ0Cpcyo2XsMJTHI/+747yJ1vP8CKr0gkHMtZAYLTN4HHF0q9dc/nsxlGAHJQvmJXFphV
yf0LXW0zFKQ+1Bt03U6+61NUxqNcXP6jqSCQNk16ryQYmkYax0MmsqfORmVaLAUbxqzW5xyqpOmI
e38DE8XsxQHdTzZ0325uisVwT2TPoA0xqkThSSYlPNyxfgfhTUfp0lM/sdXluSiYqdd3L1XtGxyU
NHQJwE/0nojvy08CzvvZNt7ygy7dGXhuq1g0fcoJ55v6kCWxvKvbkxuN6R3m0wX2+uS7HuNtoGb6
TiwUYEeQwILtv5HqGsoSqNYRVzXp8H7ejfsEgUo7ECbxw7xcxRwO36pTOOZXIv891VGSwqBUKe+R
gB6BqBpwR7eS42N45rQ6tv7+PpWTeuUy/bIJX4olO6GAzs6BG/ITB/d0H9uPQ9u8V962RcLIYIRj
CKrf+lqkzKzSUl5yt36mwjPn7iVH6osEZiSZEy2QZvR6G1VIKubq5ZbMIu/nUcil5zqwO8dLPFi1
x/jOt3I2nTABpYOOcQugCIA2LE67i2YXt6iOpuQ9CqERKZNvCdI535aKTNByYofc7zl3sCSoACi5
tXrwKk2v/0Nfv3qPdzrDO+Ln8djkna90H8RUDVYCeeYBPXXWh8MgowTsW/jIjvJx9ROlok0hEEfB
INy0NTcWjK/KVQnMkzIUURHRlcD2sJ/SIpx6nfqY6gaPFmRdZmive1dY8EyMSWa3RTNrYcAp8eng
egfwJ0VDHQNEIXcIb8qH5rXDbIwESJBGnFeSPl2bafwIKK3NN09WuL5j9KqiHV6EIRTI59n/N7pi
f2o5r151zzdeFv+EW0vzXB9fP45T+6dWMdAiuXENcOqNdZFGJqRYffLRBkhago4m5/vKF9h7BypQ
zdOFuc+THbZhLCXpQN/IQbY8tZ4vb8tT24BLmMuW32G87F68sudg2b4ZvUArNZGhYWpNTaWh0lVs
9VxE3hZnTHP0RIoOuKiREoLFyj1PEkXdsYNYqhj9fotTiidQPApqD5fTMhwJDOLhbrtaJZl/vggv
dkCofDj9XpJKOLjgUBuQV8uvqzs9qRC5fhPXS2/ECei+cUTyOMoi4nGA3xoHMMxvzcHyS/WGaQ9/
mrMKWfCfJ3nnBOMccW5vVIhEi/o7uKgd2AkmcAUh063ynJQ35LCCcyeRPmyjHLNjGDKT0FeCGRbB
n4Z2y1UqTrqw5u60WlAGIE4tTMOhfyg3L54rdfkpOSNBLQQoS7hAj1DmGW1WQEU5fbryE/BR7UqK
5ww2OjV9oYQplzGeMucYobB2MfTk1W3miFmryDFpBINJOWuA4lD/7iK7zWYrpNkzoTHTlJfrrXie
DFov+kopxadd0NWCcJmdj0vcDHv5MDtGNouCK5aJK59EHJTBnyvn4V4+r9uGsQCq58dcGOdmfbhj
YqqyPV2b2nXJ/z4zW+iWPA9qpGoHMiEzrrsFIBmcAfVz8vqYPGWAjJulS8/XyyAp10URO8k15MCd
1obgGeXxXegky8UQCERqRb5Qm1oRbejNTr1+YAirGUO4OGwh/FloEMDZrZAaq4noIOArTRldLBp9
gSQtTm+UJk3bx/r9ui5n0m+D659hMhl80DtHUYHnX2KfQ3/YmSyCZ0OoEVeRBDm6ZB8ODRcgomhQ
MoRJBN5HrzhCUX6eEhIKVrVGnPnd41ZFWLFO+qC6p23UJKPMRj/NWmdfV7ttNAgloSEGHltUKpcU
GyOkbDsUxPjN3fBpLZpZsBwMkE5w77qdC62DlvhFRDilJ5HucOClHfKUctSnEPxGTWtfyizzgXXi
MdDbOcOm+e0KAzqkgIa1qm5baKeSe0p38kxPUP+xzCYxThRPPLb7vUCI0YxRwP5AyGZB168/mPE9
7mAxaoDmG5nJNWbmq1KW/zMDwGNv4s/yUyRh244E4LLMuJUm8LrneoDiUVffijRvJBLR6w9vB6wd
URoYxTscoaVppHkRJJ2RbtFDB4ZxS/tpHSDxG9mErOORaDE8XSbIlkTI/cQkJ7n4GmqwA4dN6vjr
HWxCbTy296O6yhpyqUViDf0mqRwG2srFgpDsXZo+M2Q+ppJMmcNTSZ47tojrKbtyD8rlDrljNMJO
/QAUjsTd7BWwjATyp1ur7rHrPRJvEz8mtXaZqUwzwyNBEE2yEuyEE5Gwf5ZRTvcpGeuojTqvYbsx
YPIYwIHWD+kvVNqbub4wCT8iWZLWEcU4jI+2qFQ6b0tgvsMh8zkfq+ZZqouPVA0ElMgf1U/VhLGK
WzAi5SFpC3LsLDRVZDnOnREMgu9OI0nPgQaNS4V3H2a0s3tnLs+TeFn68CUbCGCKd243tGlNuIUe
JXloHp0gCGeAFdPMEjoo8sDPad74di8WA1Fybf7xlLoCxWZOko9V8uFgcq+FibCc6B2CK51tmRFn
SJau2qlxFawwl+P91aXjbMkEhnzthRnU8FSsD7L8v0ReWRp0h8oOXCbfGzOzkRQkdmojUCJ2Mpt4
rQvLIojMnETv86aqBVP52/Aj/4X/NZ8m8S4eOnERUQLWB9mhHCrEJDYGTkhQDUWBS7hgJWIbA4nd
VSo3Xsx4L7njKcCAmFo9jKALpL8euoFXXMvfWoBZzSuh8+26eqjooXtwKFTeQIlrpjAbo6Ta12g7
0nCJ3trNrSNFNNaSTpjIRQfsOuw/zGySIQLJpViEqfO/8KXTllARCm3o/4W+eBCE5EQJVfGmXH9x
p0NImzYuWy5hen9yvufZJBeTtNOiXBL4Q2CFvrnzUVXbnVTiguBMHqtdyJooWZPxVUIeb1Jg0e2R
zcDC8UHHCMDUJpT85DSYotOPAqYZ0Izb9JFj8j16hfwKZarMrSEA5RkoFuk/F5cOVPh1RvXWfSUp
FJff75MUQGNLTBMdV4ox+rjVkOx9eXKvj7P/G02tJ7HI5icc2qHvFUg0rpAubuNjd1SVRj5FTSp0
jZ8LMbO3Vzv792XO2beIZf9gYxJxbGRAp9l3k4Nu9eJteLf2BDph0SmZKEfBBhgzvjCfFF6cjoyM
uLWT1+f863Mjn/xofIQSNj8UotcorxwZ/ICYHRBJvkZF1WKuZcBRlvuDCnZI7JLeToEQKUwOV79T
rilDBaw/ui/dynVkEsP8PxExqLlJL3qFZJ/Sh4hOBAnxFNqCx3h8ong+iI/II5S6fIHQfMx9cAnO
kDJ9r99m/Vbry2a/jBQPveYhsj9hzF5vg4ub9dJT5LVrLrNyrNUP8GSNHepX8LO+EOoNV/NV1GaW
dTMcHHCCQIwE8HyrEnLklxcaYazSr28Qze6D6vbZJL+bkSgQQpzuGQKsJNrQ6jeFNUj9NuVBuRfj
xdONVNukye7YnXszhIvMF4/WS1jOvR+wB9N0DnxxWFfl26mVYhqNuPRdhKWnHsZT+4GIIqfUhEiq
IUJgRJQ5NKyPx12bt6VdPJGj85AipJBz6icCMBxxcuD2gi1F/U4ULglTS2aVWek+4BZZx82aQlq9
hvnL9DmsQ+G7px6CqVOQTrFzif63Zc38nDAxUnIHrIEIMMQWKGh+sKrYu64vbNSkeffz0prqpyEn
TVx5YVX24QM68/iKK6iVrkRCcHXCfQRpOKUQLWeX9zKk4HtzBtyhWYoD3S9vTFJ5HmDuYM4f8GKp
1WndgymqTcRqM3+IiJFEpnGY+NuqjNd4uo6PyYBpmflWAfCkkPMVi3rPbCrpWDw6fgnwz76OKakw
BjbpDQhi9lGr7S2MT6Bbv9qci3TUpUJMQgtmPwQgqaKkFbbMku6Sm3gZRAhtoMMWO946wxA7L3yT
aIfom8sAZHpkry5BMX78dP9ITCLYxe+Tw7B/jg431Jo+vtRuztua7cr4ZpeNfthtaS8M/ntBXAHY
fMJRCHn560Il41RyWRyZex9FHjYXVBwgUdLfiKOVLB0RxBIeck3/B4wvaI/6hSwQM8l5fMfVzyDq
PG28MEZVnEbTS8Nr88dDj8w0eZcmnq4LOgYV8nNqoUkccroeGCTZ8SmghMglBA6lV/Mr/hS4RrfT
QsVNqSvsRvgRkw1tgWO2Kd6lXm3xIcWNzMfxeUmXvxsIiPmxvZh++G0sM5ab2EjSjiyWZhMpRCFS
Q01i096IFIqXNEDEXq8rKrGyzVuAtEbJTn0hFv30ip/LbOm+JLi2MFw1tbuAF5LTcznzdeFpyQhP
glDSqIQaUtXqWPnlADfPMt40LIFdvWva69yA65UYZ+IRcjUlhTqskkIIaIVk/WSjiG5tS7K5r5O0
xDkj10eApnQszBZU1v78godvSyeL78xhxMDg2cekicdvMDv2OYBSWFz2zVJAPP1+5wnvIS3NuIux
n+QYiJ8xhTqztarvTMkBDcaXR7LWGQFlUzuj42yn5Kc9s0xV9VJq7ZOFkWQ/yBKxHq3Z8AJODjCn
b8fzqbhxkU89WhOhY04dCk84m2RPLt+vmWgv+OrlRGRws5LuCkCgMGvceEP3KBp9f3Szx18yFYbq
vrmSVhKKBBdTxZnSqx0cUvYakC6fExiCq7HpjQC+Fe/0frZpBFD5Gxly374qApl29MaoPbVWY4+f
TUlvsV1wvEmatchEL4pZc5BrUxpXZg3BYzwr4NFKhXpHGJ9U36OUeQ+qB8P9xTFinD1MdwHbMufK
mzooqD3aBp0t17uhE1LkHIUScdn0oQdyBLm1lGa0l4A4mCn6z5PTXMj9pCo3Uc29IRYERtSNlTWs
QwQiyZRLCwv0WkDoH3wiqnLU81qT5Eyb35mRBb8MQAhvC0ncXCmjkr9qWCUkNGUPvmdCAtdltx62
w7xZTpDhebsUAfhhVyASp9qg8qltYd3uKgiiNscet8Vy9PiVvjG05AOmPy3oTLKo5BLn8fNajvZi
jNLLGk6dOg1PhMYc1pTr26bcsfrnD14e5Ju9JJ5qZYywEJ5XSSJmpQuaj/MZSX3FJ5tt4PLfPwrQ
e9ItlduHvZpwa2NkigOv9S/FiNH5OO3byB+6NiwNCa+WPCOpJc7H3RHV5usdKrV2r7CMFZ8ohac7
CN7pa+9ceEb8cnq8M2mXU/oi/3cz2SvjrZUtnrMC/63mAs5C4EgndR8v9PMICQoFyiN464aBE5s0
dKVAOvKOJmm6SxVhQrV5K/zYzW9FXUv08fVjLS4ynQ95B7Sd0VX2sqPewnHNQrDJQqPVmlR+XgVM
tHMnsM9nijKXx6yohLJGaAz33UvxvJs6rUovW2X1t6lJfbkP+o8Pw4nDVDGM90KXCs6NeUFPVpMY
rn5fcTCW+k2Q38VYtGZP4CqkbT5hpBon/K54hKZoV6D8IGeZjTu3o5ZwvE5DnZr4H8rfsL6z8ig+
qhHPU0ieqcN+QfvJTUn67Py0HdICiz1lQNWsk43wb7PC+UsmZ/UR5NLAbY2eBNXixb6snPttFm7O
OhT/nEpHCtr26wUfa7s3QH6UrbDrFSertj4tkOyZKvFlkStDNtmZMYBRNnHW/xuvBQIUiWn/hbO2
kIgvUWXlvWemFh3aIQijr3uD5LxDR6pdw7Viiu3VD3OFphrh4L+qG6hpII+fwKDqlislH6MKwxnD
wAfUJWwmwi5pBQuiC9KucA8eLzDBYyiEXpBTr0Be16qc/ffyWAZhNjD56xFa8u8zG0daZg4SN/PT
fE/MXY7R+kokg/yQProNO/b56QpYd2DhcJAMgou66+upm/nDEfmyhdNgQXAwq+cvGoi6dbFnzBH1
aBUediLYraZBw0a5Sqs6QC7ug7a0wvVe7GgenbE2pUUKG24keRFkghB279v6izR5ddxoZaQIKQTj
ivnFpeVknoVZ5+WyN1dM3ANUNX1/JzGJHQbuqdN2T8+K3Uoiai7E13/25c0Q3H3jZEX1zSIZSMSf
4WZsyzZ9RYh995FrIZkWOrw1HhWu23lrOoVclfFbFir7QeT4hHz7gYAlofxcI4GSoNpjV77a6TlG
wP+IRD6DppitSNE3VJ6DmNgG9HqOUhld9jb28dIcib/IeD6EqLSGdBsWAJ/YM1PcqYRzd+0jgH/3
40tSDlvi6y2nINXP+sVQlbdZWpFql4MrU2tqCYXr2i7Sb263rfuSD8gN//wfC01Kft2dRKX+cuot
Y0uaPOHOhR+h2wJZX76XWo6WVWFBFq2EhU+i92CyNJ2Dbrc+gvyYOzAwJKlJrWVzm9fyynPtc1hg
yzVYurG574Q4YNd/ZhTHdjuxcA49QwDpqhJQSwVC8MLfaWlgvqZQMbqijNN5WKAZRD18ZNW4tXgP
/TWpB1FiJ1UahJq+hHZhXpAaDLOF1Y1AjhxU5/dVxpqJp81Kxpf28f5vTDU5Mp1JOTnTJ/ecLZHa
+TmVuLKVZZ2Ldr4e1GosDxhLKSc77SH0z5k0TuwtBJudI1dkU9zS1rzt7qVLyON/8ynajsjQhF5U
WW9OikqLrFM4EhziN4JmIy1saeD/ylarq15Q2Jf0pW4FRptafkwM2Qvy5i8fU6J3Pn/qJvzmTjUU
seh7nOzml8nbPROu8+qtr1x3yLGDqE3xyOgXGTUBIolBTsBPNBplXpkwqb1tUQsoZipg0jGEMCth
/XSF6sPyO59ZlmrotAGfCfU1soV9A78os12o91bUqXlBC2fQzbZ/gCBvI5YzpZcMEQKZE8czZRTs
CZkwcVmEyBIQFTvnRB6xrwnXsdnKt3XofMnTzKpJioyUSelIis8uH/bLi4DLN9LZr+SCANNXvXeG
TM4FUMBqBIlpN1KHwDEHlsOnmSCBfl/npYyQs0sGKkycq9mMdQj/U+sexL1ej/a0UYlZgSwUNAhp
c7S3IK02nXtVz0lVSFkjv5c1xRTVcH3+Calo1ckCvMe0pb0fQ/QMopUJXhJCgX9Nbb9ySm7s65PX
DrFBD6DNCE5dy/XHAgoztb/i82O4EtAf1xZbcg6VO8N4zOf3wCF/QLXYfLhzQZj8LDm5LIMGjULS
/aMn0f74U4tiV5mS1XFS5n5mcfQu8zaDsUBmD3IgrdLlHlPQUCzZFeiCcpW/3eTh0HUJFo1jmRhN
RyobW2uEWz37r81f/LRaHhxYjydlZlW+6P+7ZM35UPfS5vW7IhYina6gVnM1yasdztVboGYj+SrW
O3/xaFE6ymWAhJodJmx4hwnpZ4jwY9f8L5TktWkfZGaSxc2nMwpMmPqt4w3GDBr726+ex0/FjF/M
EJklLYXYr0omlau9e4nLfmbzqeBfoDC46H7Z7/Vtq0C2NuZRJ3PVTOX4VfTeKw8Y5HW+xmNH3yIy
MDHHAzR5m0GwYvUIhi81Q4IxWm7wUrXjL5e8SkIGO4dTKtwG53yMTiWIbqC0dLzBFnLBKFeEPLO8
D+2U1ib6AQ+cxjVnAbzYdDyppEaaUnZ1lPE8etrfgRKceSUAw9bUislIiDwHCrFMfBl4NsfXNIS4
Bwsein2362lB6y7hEa5zXQpKy0i8QTz9fUQmISnBp8mpRDunl/V4z36F53xL+vD+8UniYUwP3pFg
xltCny6f0L4Jek7bU2zVvB0NzGtIbtDZv/dLeo8iV+LEaEt9oheZrjzKwSq6FH5iWBY35eBp5lt/
E1wG6iQDhfw/JLCVqQcv5ijSK2Oma2T0EtkNfndFcSuFXzwGD5Wze1IzTaT9aJ5qtalY4baUJFWp
WHCG8e55F1T2MVwki11j/Fic+iR86iLJU/ciunmSo6LSs2CNYSYAQYqW24UpPNB250xN/8j7AuMI
Y8gjdS8ulD1ZqD4836q1sVdgUUn+OgGdT/p3FISsAbX91+qqnP/VzUOZ46QI4BYoUEE0BQFVI4rN
kcnzX35W0MZ5H+78CttBo7PXjdC/Cx2VMgOF9tzhIiMJI0T9HhMA21N/ygQlFKOvVm2BZXMJkcuU
5pLijm98OHGfusy8pLDIdjEmGTSIL0hpX9ZFrQarJJThhFr+JPmC36plWTeoMqo8mD7LSZIMra+b
nfeMvYbXvNc0QGe4RWI8ZQk4b2l3l0IvNoS6qmdrtUVXgbW6ABt1rgwDcC5KfgeCcHPp3uHC1hGH
XtgY1oKkyv/grEUGeOABrYS5trEbdwxW0mCBkUG/IKzcy4CCdnds9lDUmIAu9gZO5Ww8cc/b/eGH
17OcEy3jmewoqcF95tEwps/oFH1Hg/555ybTCnkD8Quhu9BHZa4v4ufwvbwOHsQ0NIyX28Cqm+xe
WLT8Lgwzk9ywty0CrZ8wLWA0DsXlozujGzPFSVqh9l3Icmas6NdenTOe9z2Nvjlua4T289J91ZVo
zLaJMONOgA+Pc3AGbT4yPuTb1SkZXUyM8zH6G6jp3Bi2zyyb5DUuVCjosgz2hCkSLadEZROPXNAc
LrILXPfSZv8Y6h41ZFQAq4ms5inaP7dyDYGIV3AzRhTfxiVqmj0Q59DrHqv5tQIpswQAjkjOcMbx
dI/nZyXk7fKzpW586rwiBVe1GoYrrL3h9qrW+IexRf5ks7rFZcVX4kxjl1EkrTV2WC8NQSJCkADX
Om1bZq7HSEHIsiAccgwl0KhBurXSN+0wZRI3GLmROM1p92o3BYwZQd9QbVEl6Siu2whN9oyLGMUW
IDGtqSFEUufoHgQhrDlsnj7sypZV52dZcbMcdd0wzvO5rKSJ5KvNrtXoZ5NFtpKfcH+pnYMoxdZ5
YTPY73euFZIGyXeHSvMR62/zBcuwaz4lrGmwv5K0LjD0XZ8NUPGyiHqs8cZHEhxsbAJdpZX/WGqj
u7msULajs6J70VLlPWico+H1DNPegqrOIexlX9e5I0sKmd7ShxEy9AQIjVVyof0/Px82Ccbzabsb
0HuBKeyohEr9+21NnPewqrWwoOUhm1353EtMVf4kBLVjAYwRNRY/r5Sq1YVMzEsKr3G3R6zNEjOv
OGWHoG9LLBuh3zDWEiSYE5N3DhD2zlYnMEEHO4VLUuEBxGyzHKDrCFHCHwLEeO0Ya+Q4Mj4/gyUP
BWIHViOHJwTd/BLTuieW/tLLS2hkl9K+J3DcjmRXf9/um7PHtMRj65SPiaHAbVj2QU3j5cYu7UCE
RDR7jTUzqx0ekoBEUShKVDKsqvX5Zq83lHsfo5flnrQvjm4KMj4cb1Oqi6xClTSpx2ur6mPHS77W
xNfP384Ya8h2I8Y09xdjmQtc6VDcFGz5ImgjZ12sAtb7vhtk6+DVdSwC214PO0WLEuzKlFxvcPvm
vKIIv8gsHwydzf7X7kjlYpJnV507cRrS7t1On9NH1H6V1E5nMwMULvg5FA0u11XK6PVGJY7r04a9
bwvOI9CJIVh1+AhQDgyFX0IZN7YJ+g6FboSOOsfs8q17pYKcysXOnYFOjXiHkMkLNTuNqv1cuvno
mEIazWVh0W42KhJ9AaFADbWvhN1YLbflMHdBqWf7G5mt5c72ROaSS/8XpUm/I09dTu14s1t5eKw9
2R+NNOZi6xogK79v/fKF8Huk42oC8fnYzkEeecZtZT7ZIsN7W/4bgZjHbnGMhmwwr2N1ZPB+1Nx3
ae3+3zTYiPwP1YOvTnAly/XVSk93vOH/Kja5olYtC5fUGY23vcOIIzpi105c68PjTzeKlLpOGHUz
kXaBU/hIvW65ZbAp0bygvJn6SvHcalpjzAIRuESjZO2ccv4wHS2ZvMXDS7DBSKY2cNSYYDtR+NkC
aqgnKwECYd/BFC+nQGLRlvbn8CzvX7Reu95WoqSBolpUmyQY9lYVpiwJ3+MauR7HV1mJUgc1KNmL
/6AftfUxIdH/gRW+Fyknw7k8TLD3N1es0098CKTHMYlEiPhlWEWu4UuuBPpBI+YGdrE9vmRsUx9M
ZCFZkHHDdJkYxCBoZryGDy2zWLXiJlGk2tQGBkm/Xbp9Qmag4NNw30u0bBrShzpi9J07qtJfJq6Q
H3ZBtWTA76+s0P903VGbx9Mn+YVN6F0RfAr92XUxCek7/dpNsjAga3BoBZonATnuYL6nvH0qeiwN
IznIHBKrEL4F4DUE+zBkjSlqFug8V4WoFT9zetjPWECyXf0oMLOHDqfSzRCx2mVr+1bwNaeFuu5G
l2Gfi7jntuY5XoehpQLaXCz39/w3evY3JndXuo67jxngYce0+/B1/6wE3euY7Rn5vRj9ngmqsVG+
IMdYlCyRxxixlGNXJo4tgKhDaffQ24OqphcrnSWuH5qTsPPGojEBMoDZDfRAP47shf9tXVNgGrd0
pAqLNLdNnYljVSezh4acEc5+NH0QBgKiBCDn4uFbjW9tp6KE7gJK93byMrEUaiXG+tA9zfN0cLrl
q65Vaoqw3oe95xMOwwt+BlYN1PKRcuSP3IECjOG7WBO5btVD7tLxTGhEJ1VywRxmeQcrvk0MMWB0
QnZDtALSsDkSdFGjty/QlWwXs7/sS6kEvQJyTSW9igkl8Es3kGybTrSgRFFCgUk0IE0F7rtacDIM
6KGG8QNNxHOp5lSlhKogh5zWeTaDNKDkwqzja6U2HGAWBGzgpDjx0Ez9ky0/nE7aJWruxmTEMkrY
jwlo+JnPDR0ZE/NjxrpvWQ0FWvmzmHTaT4GtmxfRHezbgYtqT+MFN6eqFnCQTTYEJvTp6MhbXJ1g
ByIMD0NNny25WtY/+TXk3HxVr2pzM8vmA8nxUAx1RUhWqYhHoP++TF/OEYdodBm87xmpg6wXEM6i
g0e2wg+O5hqSSz1mi1360+Ps8uiHgd0zAPj0X/CN5Al5m06r6Ko+5QRgLUMYK4zWnQWpa2JxKvsY
pXp4SBQIkmzSrZH0s3vkm4hxqSUfbCM/AaM9fqALn2FM++TGpkOLjQUJ4xlJCon8iLvcaN8PnGr/
7RhgakfY94bpLgTa403TKOccgfCkmqUUIOD0ajrunGaFhqBeU+numWBFcijBBnGCaInB3l9YiUOb
e8NnR77vqADGJ+pZ2c+sg3yTN9RraBBEoqC2ObykBEmXzQ4Rnpb+4Z7LCrJ6IkRpaav2x9TnLeYB
w3SWKhGmPsfxIiZMntAw7+LC1TD0k9BaFzeJZ/FUjwfF7sVm91giSvba7ey63ABtuwqEkTBORzIC
6vApwxX/wrFo40mRt6QkeRWPxVmhTlmtAv0nE54rCKc48Acqhdb8/6Nyu6mZ3tgOo8BhYyrjg7UK
2EhWzn+5ivs0h+ofGIQfcpVA3NI0l65/eaIYl09ssPigU2FWSWSB20AppF2KKmBU96JjV+YiPOsP
10ep0njKNST1Q3ksn+mlAByInQfoymSvU36nBTAuR6sJJwvpCMammKrTXirCvnnrn9wTG7PksivL
MLRsP+uXfM/B3KNfmIvVoVxnrnAFxm46s222WA8Rx0nWNRgBxPk1/IolPr19ahVIg6gyTPO96LhN
ALEkX3OYOOgbpThCGQkt3ilZGSwVOeVjBm7XJkuYu8c+gOSLkC2hs1804F3AxDggZPXGBu6FAWnd
l/myKsnCIf1MMCIs6K9WU74PwaRln3KfsXvojrYx5bNH6u6knkXKQDOVyneVAdunqbd4T2foGbii
a48QiME4XmFClUajQQnkYe9MINrQy19jmSvSLfGqIPbGmjp21fmtnZRyCT8pF+qzBc0TDG/WuHCX
LnddJYujG5z+P1hoLqmMivR2S7qryRPjgXApn7xp3KGW24e/pEjnGw+8ooMGHgJiVKapnr2d9Q7E
X73swX+6KmnG8Mb8EFqPLbZ2T6pts8IJEZtY+bjZxiB5pudLM0ueezI4ROqH+HrO4iFKMQNkEL0L
N9qicD7sbRozw80uu4DCrzI8/R2LG4VKTg8DoIEwbU2OogVVW7QP8S0JE39q1QdOsm2+bTjP3+Iw
Sra7G1ivuZhns+gO/tjFiqOvfSCqLKVIf1b80kVw3nKm/26kzCU4WIzSrj1QTuHsXEO2d3B8Ey3R
rrzNArVCQQ+gA7xhTn7YQ2Nm9ApiyINOWMFkhzVoNQDDLXJXmyXlEBn5TmjegZ9tsKGDn3NdgBzO
PRJUh7f2qvvJ8b//xyo7bmeWIQuqm9oEbBcFeQOEoDgQJuzS36Ebbp9epXxbULr7DCcJROwg9UQX
Wj2ZngbUToKG2tCOVCT3SsbZFJihn34FwSP+syELqQsztrKaQd0+8xPedW4DIotm2uiEJ/Kqf32g
xGPmR6I1LxE3mxYiPQjZJf7rMgGJQdoLkKypFhbUhkxeXi8cIZLxOJomTV7gBZr39oiYH3YBTHMa
60AIZwdygT00SDKMC1WL6Mr817fUinq5Efz6l8LOWf3uHQ8DLQdhfLgM0zMpUGWo2fAUpluawbbn
pSi3tSn+UrWn5a5T4FUpYMdj5K5n1njzMRWlk1q+CbRCMRXltUmnLVcp1gLnBY2OlfrcP8XBZabk
Fytv1cIg/153lzP0MC9fZLnM2Y7VJWSRAOWG/ayV4MFw5W87/63PHiakDaCGI1lndyJvuxKdAHZV
MHU/MrTSjSEnJAM9dweG/FDPGBIyuqyjpKKW37Jk4dQS+ymjjau8ct7ATDCCaEf8rb3OS9glEP7M
jMyXW7ihU4g216rRZHVoIjrZoijcKUzwDbsf9qW8GQx3OB/maI4IgcPBCcehyjUz//sxZCX0zRRZ
W5FtO3fUs2udbU1DAGl8KUoQPnopHILxh+6MSkMfrCTNX9Te/tmcvALG33CqKW0vro8faUqEaTgO
JcoTPgIw4YkAjQiUl2FXPAU4p+wG1fOs64pftxjQbFJ0CeDF/q55pzHxe4Saj7HZ/Rfinjo7FOZm
HJbhpb1Baoq2FnCVwPYvSnYaCqAR2S7nTeuUC1CdEBzwQawRGbstDUukpwHgLtFG6c6yTIpMoyZC
t1qbUPXZInCebkvrZZ2atEdvoTj9tlDEsRt6V/WcGPApNeWeVWpJxscNLS1Fk8BF96PNfg3uY51Q
oGc2DFfz80uJVOSQTXRqVRxEMcB9sE+KFy5ctR19JEyIMN65iS6AjFUuLYW0iP/xs5fj86dMKvfA
A4RqgSOAAPmGHRXOITDHBfuIIGImOpTiRBwcWCRITRFMycN1U+KJTmEGqqNJodC9TvtZkR7NlM77
+CR9tWeOTSrpatvSl7680K0ZkSbqIDnFi6zM6EVqWTWmQEvo2Bs3z9ZBW1Wdcb53kqMQCXWvKXn4
Hkqd4sE7NQnT1y+uL5mELTU94oX4DCErawrKUmPN1+9EggQmh6KQwwCZWu52o9N87+LcFYgiZ0SS
ruXR9+HI2kfyN9+stMXUXj9j2nqkSfaFFCBjJ/f4tusZGNHQ2o1bgEPuoAfrhyzpZZLviLe2P/9A
Lgl1sBFTMh8gYV+bYv43RIFVfaypzGVHxQ1gtVZgsyUyVaghixAZ1TLEhNbnVrN/8OugrctVKZoB
qwpbD6nySUYheF+VVrNIgzLmVwkR+nGyw9ZCU5fHlMnaJaAZm8mwWiPqbaCYxcFNtrr08CyoaJ+I
qeUc5ZpGjsWzyMnoKR4g6CXU9nUoJnkGGd1fhQRFLLgbSlJVP1iyYI998lDR7kgOrcgdqet5laZy
ONJZTu16BnjQ7T715ALitfq9TRyl9HSUfkMreMm4rPJJokUxFbwZyOiDrTPKUSYLHVjpiY6reMDp
1c4QOvcsfAb7CLZmTtKZPKCQZJ7ux6FnzIIv7ahMgUDrDhy2oMa9DitcsrXr4V/ny1vBFN6F+NLv
V9eFgGhOQo5PlkH+QrkAU9Q/OBglibg+Fa+y9Ccsq0Ktv/S2q8MzSddCmYwoHRs2vHJBAavfYZCG
fJO2T/CWqn4N0s7s08j5ApHyYPPcaqMoNau4ACeVTG7KqKMAjUnftc4iUtg4gHX3Td0YDGNikfFw
1vZPncOCzS4UISPGe63Wrgn/l++y0OaNtJBC3TPbfbzTLO8poJVyU9NLiHIGcKIxAOTpuiQ7HfKv
WvlZhiCgG4j+TXM1RtM5vfIU6MbxVSuj+Y6dvmb5JeufZPdarCyr21Bu4JAV1WWKKigSsqyAoIOB
MQqL5EH0YlKvStor6O6+/ai6SZqCiruVK2n/emrdt74cdDij4eFqBai3RHNMepVKghYN7cKtE0Fi
6kldSF6O3SKVz6/LI1n3c2oeDcJLbihN4tFt4X3aDfDzqNxhRUf51vdCUdtPNlwA/ZMxRVQSvB8I
UZAI8FNp3pRMhpnav7JvHZOZa6MXMpLjlBPShMRuq03o8vDdhLmQ+iIyum7zuKqvnedLTthP8/iO
ulAj1Y90VAFvHZA8VENK8iCb91V8b360KhVQy6mQ3UYDIvPr+w4qLiVH2Cxyw7Dou3botnXyurPw
OVVflRDTgGDgvl5eVSnQGUlKlEBT2U0zwJf7fq2DVRjNbw5J8HDPx1m5Q+pfCtc3c5qb7fC25uO3
Lrwn5iaiNapfb/Kg738O4VG+8zTvB8z43AtZ9eTx8FkgbHqe5jXk9NzxLvbeKvrAgANPDs0JcO+z
xTE3V3WR+lIpWYJVsgYUK63x15PKNa1R0hXmtzxkPLtK3cCBuP5x5pOzl2Fbv83fBaWtWe27xKn0
58tDKAXKZlNugjgUv4lOKKkZbVObYilhUTWjGCkbyBmO12LihRyfcSDWfghKb70H41WRKpFl6qvE
TM1mFiFqPt8LoRVrBujDRYXiZbLBwm+vlr5jT1D607ntMcdGiooh8lc0Nu2Vk3OaBcCKJhWN8To1
wO+GdUwVlWCGzgYeBQIsE5RueNoF1BMacLr81CoAXFjSuasBWOpVuqEhn69BcEeN/WQWabvBXs1x
OURyM4z7KJc4FIRKmCch1AwftAgl4ofrPuLjk/pLBZD9e3jK+V6whQim/QE9kLmF+0YFYoitghxi
ynMk8KYvptEOcMd02ZZ/M+r+TNjA8Bt2IYDQoGoNb4QwriXOYYw4q1fz2EjuR81gEoQArwr8Iofk
bO84M7BMn6qo1eOs9y35AfEoD3vHAFiL3lyO+56UDj20uVfOYi6VnTSIzN+fqaonzL6Rhf6DNd8c
aMNRiV2GGQenDkkiCY1e0XkSuRVV9P0ByFD0qHbBy7r+DqBcV9vmnSYI5UCE6xrz9hBAO4mdjuoP
pwUUnsO42KT3I4CpCWsZw57FkVQ9343GwUUY1yQEPnKHbtgaQ6zDWl45w90EWEd1ZhiyNzuRPIHU
qBDa3YC7/A6VPZGMab2GiIls15HOAogK+I+q3xWm2u7SOjrSEh+3NFrs3JI+b84FyQ9AwKAHtyuj
64DlQOpmVyXFfEfBN/kdda0RogPs4/C+f5u6acWBJvpMYy5/E0TTgjH84ylFQeRUrJmSA9nsW/h2
xT4Wnh/tTk5BeajyZILuYaPbXyRy5llAvASzwBTPsV2hBIZquKqSQvwDhmp0VPqURYDvK6Dd9EZo
floWM3m2KwIyfYZ0J5st8BqmccJIa1Nz8RH52jiDK6ilTG1pGz7s9+PuRM3dqswXQxbngEVFiBSd
SzkWArLVT55WNxIUuF1O1c46xs42bF9HnFVhjTG9ZDrlq9oGQLBex1eOKYPAyM4zTnVx62sz3wcI
gy020vi2RrO1AbGAjgExO1SNYKJElG3/tCvIjwYUSdwu5YHm4TVz5moES9KKl4fv5AX0VDP8fM8Q
MaA+KYksDALDut5xQSIzuEnximgWhs+seNeGU52lbI6azdN1sZlh+ewJuZAvylLclX9pr7rNZfbW
Fs1g7xPVNgCjD6mwHDXkXMMZclHNz11pQD32/DWcdbCgG1v86jJi8NBuRsFofoJ9hEexuEfzlzVa
ZkjWvvCz+fL4cxflPEtJT649F6f30lixQcrM8BYBcLyKksx6NOQ3MF8E0O8bGfKYPnA+K1OSimcR
iWWQen8M9SEmJzxdLLnQRkUg5X9o/62paZrBBX5/83pVRmDp4seNNKcAXi4AQMeA0vxZ8EkavxCm
Tt6VH/I7uITvy96SUCLGjYa7tRRZczsUUUsMKbQkkDa86i+bq9sl6wc6KgH7AmWO1o7ZfUXauW3r
1MaYq4QUl/Q4pMu5OJBcXq3rlLbZElYMYbLYATSnAwP0DNSPR7ceaNmifcPU6Tbkmq0E7ZgVVZ/a
m2JQG30Bibq+0RX08eVj6p8ZsmHcJkcBHpcGvfJUeIShsi7kl82LGDnjW3C635Sj7UNkqvmhycwx
AD81mCg1arJI3lJFbj0KkH2S2myQEFhgyLMov2cSNoWuxiD/e3JbCcJCsS0GlMn5fkwf8sMd+7wy
7B5jX8EzukHsbXeaVepUkL9XDR4cljQs+c+rc6eY/cNSRJLn2VDctx0N4sppVsHYCZd/ZW+wI9w5
lxypNhT1GmQjcxBR+Z4Nu/g/2T2tGtIBREmtIJsH4umXmR/CQfJf92HGSup1ankE0TV+Ce1yxVQQ
u/GHGPpcVFAAe6mTID2xWjuqrPLvZl196kNj4VoXt4RUqXhLZh2dsvbj4xkEEs38mxM5dCQdtYFa
OgxJsi+HfqGDz0snKGHRPHcQT6I6WtsZJA17AD5c9wkzFHPtT8/4O9MRbXAMM1WnGUnU9FbvHQyn
aueolX6y0SlzXm51gGPob4Ddg5HSEINoVFzJ1yExOipcuNIplartsWIgZmLFBe70qjcU8VZMNzQv
Z+y3hQl5XNsV3A5iyo3h/BUaG8bg+UZecqHosjqYQgUiCqHeXw6+CwgW7+gMWVeEOM2pHnwOkNVn
lp+bMo9GwflaK23/oI+g7B/BFL3+vL2oxA0xQptnfMdOng8yp4PmZDvnrTZGxjNcPaQq3Ka4JRda
XGOF7Qc+2JOsszj6Xl+igYsj7sO69Yi+R45xEb5TOQ7pl6pksR7EWwRc+HzP60LS5aF2VtnYFk0l
lPOG0NkeddBCMj/LiNd88eE/fKuUp+jlYstibUk/cuue7eHVfxwemXL7S0MAni4bW3Rw7ZgnZqgm
lTA0HriamSaLRHaR1deRnQUcGgi79y5wJkG43rLxEsOzi57hGb4nl70q/yKjzxh/iuM9bDqUSZRK
lrC5DvSD4qW1dPZdyibPvgYTZ6YmMxpK36SlmUKGWHqkjaAU6rKFvDwS26LFO41bBiCBN4gM8Nl4
Y6/8XBaJ8kiY5jHbueHcv0vJ6g82L5D4Cfd95XpKEfHGJQy1sR3XFaegzHgYBfvw8jg49ooVrKgf
oZ14/lhto3qePDFyvie0UIJ9fFeH67EejXe7XtAXt3hJlA9KXeQh9i5exOM8L7w9BZTdVU8gW04g
xKdEs5ePW9y18jhKYV0tC7VAJENw1K7MT38oeiIqpN1d6GHU067Bgc+UI6Ybx0UpECcWN22CzYLE
JLyIz8AJCscoCO6Kh36ynUozj1EOPScltUjQCyq3gXd3Gm75nwkq2FWeEGUmWsQAlEZ1NBowWc8c
cwZT2MIbu2vekfsw7p9Wnmwap5NwIHjcV7PrrVy0RCGAwIfzIoaS7PJ3xYh1FgYVcD8uMqmiMk/6
vB/tKMEJjr5VPQuq++XQsFp5An4gJXA0YASmxsbf7cH/1n5ahiyBt8O5mcZdxPZEu9BtgEHIPbhm
hH+v+3gd0VZSj8UKiQHkQKaSkJ8aKmMI1XGXSJO5iYyxl0Vjghxnfh8uf4+mqnN23KHLvRHFDunn
2jxq5T6BqbruEBE+S1KBxEobv2HXNtdM4LT1mxpUuTx6vc9Qyrt7UjokLj/Qs87llCGUiaC9tV0m
K5wlX5SMW1xQ3xnSLl3IyheF9FUpmNHxMZpw6p7Kvg/ILC8VGT0zLsZ8AymAaAhZ5xQinhzs51Bu
FLzFZGhXpQNBghDbdbKN7rwjNVjh5zDmYO9fZZTOxC3nNzrDMLJ58K2KUfgXs80zNufAW/oyT62/
2DEfGhZtGoqXl9NJnXu4u9dufB9nsJb6bWbgwWHBvLy38X33i7smSUejoSEiueUtNoCCMq1RCV1i
3gGpTWKdwcOSgHvtzO0ppg/I/xDBcEo596VvcdsOkzynCbZ9Cmt5gWIqFqpOBvCJHpcVLh0I+Bms
+wiyINkyLAao3Ubhc+G1XVfy5eRPKAJqXDFPoZ++TJWF2Mx4tjB1qqzCHzLDKvsYyn/gT3XEZKOc
qKiptzXkie6kIasrHr10X0o9EU+u0JQNxc6vGmhw3EjkL5X1rursy1B7ldzVJVxPqPXfjsfpTcyO
MhD/6ieZlVyeGk2eQ9Win42F3GtQgcBQcS5EfYazNZ7v6yqx2BpmAJ6J33dbdyT6g2lGY+VuRf5K
fwIegcKtAM0scE09E7hFGgm/0izNGJOaUIlUgJY7w69yJx0twqQRNCyAu/rEVCC2+gX7PqMyAs2q
+Pjm2yjWrgG6+uQWFL+/8fIvHYk60bBNESbsVix6QNSVNxBHhoy+f5vf6JyuAI9ZKp8SqIT2Ksdl
QMZnDYyhtvQm6sNKGOFDuhXsffOyaPj1ILENTARQAVAzK9boSViBxomfT0TmAkLc4VwA8lucJVQD
uuz4prniNK2vv96CLIZzlvWf4Qoy+jK3ZzdAbN+FpoYEh7589N+sdSI+uHn84KM4XNwPCgsch1OP
uvNN/PObvtri7fIhC3OCXnKTVKkUEfMWSssymB5NpHn0m8AXYFaFExp+KB1aE0o88se5dxryHV3D
ycio2nVOcI4cISHmTdKcNh72ntcxGmCMf7oRB7i24JVANhokAlribYA64Z9lmmFGmaaw0CK/jtmP
/9NiyGgWTslTb++iqIoYrYwkJRpYz1eINXaWJ+ZKZe5xFyzXPT4UZtXhFc29LDM564yMWvuXtasL
naYwxyWO/09UcfDP6pKUiVNPMgKQ2/8hydjW/+zLi4ZVgSleBlK2kBewDCq4J9709FSWEUB0SxuM
G5Spd6ywSpM1ngoOevaDKrrUwJ37O62tiBQ4ZOUap9Lfxlqo8ugyJTAR1h7wpl+o1L9QsUiOV2jQ
ltiY62R+F3CInCM4GP7ABuB44R0iTbt25fLLfmGYSUTReF9ylacrHDEtPVlodRQOAlwGkYK7Ival
fpsHkGY05h9iGbDpgYMHovHNc31zfMXUjWzDQWnVAA3YB3B4203WUracKCHRRMoO4vEdM3VeL7Nl
ZEy7Jzio1GXsAl6m3HxDNfyVIGDQYgY/SQnfxG6EOxUfCRpWmHX7j/9+KTRZwZbC9y3XGAWLo+aj
oRTBzRUl6uybNgW4HuHisGKF/XAI9krU7o9ZMw4GSFwCzUt26U4WuKVUKL5QCAt4YxVupJcAE3e7
ZRZc16BMxAYX3WSz1jWH/HB4NcxM9MihZxucqAvHrXxAw3kuNuJRbsTRsIhsceHZowAX7nQkG4wh
HlB8LtCju0KK6gwxAzvfGD/ji8f5SsnoOn1L2T8w2Vshf/LQKQm0qyMgJ9bn9okq+nf17MAXNo85
ur4XWb8JTk8oYSMdEQuHFwD3pbf6OsB5SXfj0q6bEekFAJLqRAx3V5f+kgAs/j9kw3LTaFBoXMJ3
ltHxfHeSC6coSi6F9iJ98kFaH+OdgdM8Mc48w1X2GCN9yH7pUU+qByZBp7zZaaHhUNyRiw7mnnd6
CQio6LYF6rhA8MQhiS7TEh2Q06VRu1OipAcyOZJE/m9E6/n5sGpETax1yalNOa0H0JX5WSmpYNfy
SOrUv9Cj/6NaITFMFOOoeY/Jde4wkQEJ3u2rGXPjnSkAvWXxUfY2Y/JZQI8HQXGPm5Jbn0EyzDxw
N1/8e7E6yT2VRaF762TdU7vrleCZ98KBuTZVDjWzinoy+ja+5FWG73um+cdub5cerBQ68gBZS9Na
DNME7vMOer6197roHdSeySGE1p26bdohCm00Z/eNsOK832lE7Hyrpf1xE4kdDYuWR0sxnxkSiA+U
4LXNEuu802bkwKlQAmfAlctLEc2zCJPRmHxuFQIBjxpEoc6yVzqcgG0Y8wIhkYtOfc6Nn32tjz23
NMaDwjMRTP17XZBKVOz1ArAiPVMgGq7kxzz9HnN/i8yFswsVvtcoTQzIBj6n789Ux1WmTrQ2/nFA
y2ukwVcP/ba+T3IiBxhMvsaoGLJX/PoZTEGbjV6YkTuvLgI9rGn+pP5pCZMiypX9uxzOddCb9bpN
B8lhf8fPkiE9A0JzPpFtjEXci9ackq9m+sfUrYNx0mj7Gggc36rFLVaJjmxKnSVNQwXFCcXvr9hi
YIPkeljl3wkJnJrqxizUpjsoRuVEZD64MBx7TA5bFSF7IkpgbgTjlNovmPDNZPWs8FtGcb9EqZ0R
L/0zUNIOphKeROxO+l0JXhQWgAZ9izsiaph3gAWeBp97f/NNqXR5vD/3upy1J1XBnLtBkyAiinAP
oaKab04w/ZE4+cMp8urrsd4Kvojq5Ifh1zh9cbM5Y5ripnhWfaIvHji+/ne7/ePnWEMagCdk7WQ4
TLAzIHf0/1KURJazaGcEzOYLzMofhgYIh9qcLTpq9s9aG01nj0t87cJtlgyoz3b4lIgyv/uYoMul
wTSwL8W8qw3xPcpL8EnUPBGGOXukTtVXuj8k/FNXt3la/XxntEvvTmSW+nhNqMe0xysP9ryhYDtx
atTfNiSGzKqGNysZzNNf27cNnu7zzk1fN1QlYWnouK5+l7mPMT3IbDYu7kag6hdOxhce91GHKZpF
3f5NCOSzyKiiriRvbHECx+jCOL3vELIG2BAjznixLOuPO5I95qtZjQd9AIBU3RSJCltovXCIHYvB
InWspCPdPvhFwdKNb28Xe64ATkbI4G42TZ0MFRB+gBWLhjTVWat78WwxZjwDj7X0gU3qKD0pNYg3
78V7MAYkIse4W4kdEHVBUYkCRdUO8whrTWx6pj78wm9vI5cUnpKoUnBOAXpro6QzYsej1ksh1mZg
nDJ2pcs39nJmSKatQmr/oNGKNpvX5SxLoRWVcUbKtRPtoIP2DN/3m/1AagxrFgzvukmS1DQQGdLZ
6EqwZ2u8AbAkkVu7GSNLGKLXFOrTYEJh6PmDKDwg4ezTlXQTrloKqTdTSceQ4gUq8gMazJowOK0n
ycfEHR22PxSLw3BHmn7HmuOxv9/oHkv4j0TEI696WrJIk3aguPwa+AuOwdxMCmnKBhej9ySoVLza
P1o6WHh7wLHi/eph0QEmlNGwWnvWwiZ0BYOD8w/oAcqPL5moT2Q6Qps10JRzuULcDNPU9JjIdlvk
qzsxpHC4mdYp/GkiqfswMoYnVDs26ZHFUTpYotqRD0jD/3n0hiwmx6Jb5Ij9yzna7NFLLyRvYrOs
u6H2Lq2Il+izRvLaCAAy7E+3ShrKyHumpfptWUCFPHrBNYKTm19UTvFFOgyKoM/9Hl3M9Iua9hKk
tHQT20eciWIX4EZbUZc4gqSU0m9advMZsYN2wMoL30Je4H3Si6SU/TO2ZyLmFTOo3sTE60kQXe4x
RKV1ue6Z5t03jsdBXs0Iar9GcWr9JxA3QO1QT71ItDfFqrpCdqDNQW/xUNud6hN5a1WnpcZGZdzw
d+pte5c+e2MaP1cV+SqdXGMg+tU0zOxOnk9LYuF+yPQYEvSHVAAPDbwZ6OhUsvzE36JC8kEqbR0u
R+U53jtb8d+Xz1NYUx9r5IzXI6LRwd9VWjRvTac27iS87nG9QKHqV7IUogKnyGRG0c1znQvRUHLe
sR25e/o5EUXCG3xp0xRqGnK58xnDLYlJRo+t0CZQ+Loyq6oIYRyA/PoFkLw3BTHE24GeJIaDLFIJ
bG+WjBDYstl70VeHQBoMpqqQ55ezUmPM8nUbXqxcimpoAjYF3t7ug89pvEmBK7ZRdLiALzPb1zA+
42YDttZ7rT/vFfdOICOWIc58PsnK9FsstXjRO4WlHuG3Db+s75nPXkA63neFDFjbEZ9/ZXXPGcv/
sfABiTgqB5t+I/mpZFpxc/MLLXYPwSxX7B1HSqH3EN9Bn0k2FE/jGNuT/yfB57gQVBcP8sNhNjv3
bAtzgU0tGZ3brzAwvvgIPMvwiQNlWuOtUXU96bG5oIMOLvXC7u2E4wSiolP5sL0r8fZ7N0Qkir++
FSuCreuX52rEiW7egryJg3V9Fv97DEkpQ6fTMFsSQ4jQWGTX/NzVQ/ZCRQsFo/NmACBOegqTIMX/
e0POQcg0S/dSGG8QdnJTpWQcsvNGK/6dnJO3IXirqHzO4N+6HaID2rXkpfRJu7neGnYLUt4RG1t7
jp2FrsJS5I1wOLPtP8FyV+zJUxHHpfGTz+rolHPUnYZV/gliTuu89deiNoLQ8kw9oNR6vi1qnwIB
LlE948NaqsoRSlu5b1c4jFfMBH9IWRQMqswl5xYYXNtxyrL/d77hfxXk0jlH9KaXG9HWRCHViYm3
w9UIeyeknnbwzETFlVBN4qUt53owVH72F0+CtE4xPxQ8WKhKE7Qit+601hVW8S/yssm+A8euMmq5
q2l9PoaGPEF1owfQMw7oOCfHEVv/C6olTQqDtGdQL2/Bb1l74RiCtl0tl/pGRfpixTN2RYWJtmXA
HYCmkLHet9WKZvs10AX52PoK8Z9ZgW2ZmwXlB33ClOfXtFfuZDOb7OkMZoXmTwjVwqrVjGd6l2+W
/gEL/UkcKsXnPtskVxRyOo1I472qkO2PavaaiAcW52/MXRZ4G9CrlgH9dUfDRgKZQDUxNhRyPbgn
pakniBOqGcobLteQNb6KhqswqNTTXup9ro2YrlYFIhfDYerCjxBZ3eig0UvPQGgWU8CJYhnCUziY
oMce24jbY0KYSMHgZK0Wt90SQ6pFffYmf3BWH9T6PQsM+2ezXenpXtiLoIWaiCZE2rg1gGSR2bf+
9oOxQErLhGe2lkJr48XDrp3sxcKrVigJjfvbCf/CN1kQHCS2ll8sI+nI5WEZIlSKevnSCvUfmq1m
AWsdQQnpAZN431nZm03wX4Fy/aCSdT16zvDxUZWEBofIA+nzH4KUeNJ5kxDM2B07lVVolCPp2SP1
qSmT/+YGb//NAZkjd7sxQ04OvQyjCCCd1Q8iTXW+zZOsjbSNlpGhG39wqKBjPybqlq94cIfFEKas
Ow001OJJxkdWHyW7pozMoCNkVfnq9q5cldcWFe/dpXv/LXCtSszX2AzGsqTomR//MAE5Y7OuhE8t
CqMJfhXpVOd08WbNgyIXtS3z4aurFgScbt2fUDs5DZvC9kaTwD5NG+8oM+uu+j1lwSuYo7U5szha
Psbhj1K/7kAFodoxz3nvtYn7+BDtYiwHef6QLcumCDKco3yPaM9TTuY73YWoHKxkEkf0eDOA+eQd
6RYoJlWtef3Vv7tNIvFeJ4W/5EvjUNzCOKjsWk/S34F/UCEmnvp3JT7osJ1zSNhuAzirr4xlljYo
qjAdOo/Em5Iu/asI9PEll3MT6ImqFOCgE2Id3J8qQcgvN+5uo29e3f4lvFJ0WYHScBboRmNr+/nA
eBecQWPEXO5CzPS/Kt7CzWXfpg1r1Kjk7KH33XuXApqwZOFiHq/SL8YfbizAXRNevupK+YEFbVM6
etGIB4Jiu+pEQ49WvvXJR4x82vnjwLNg3uT+tmd2zYa99wu3sI4PYZXAsf2FcQTODQGt795ZxxoL
ND/HXGObBS9VilpJKeUxdwXR3wQnxeFXmaMbGSYbt49W9h9lt1SQKQ1rxoT7A3FdsOp3mYU0u3yK
Qhdx+5boz2Iqf9ABGIR6aD3oeF6C9LC2Y0VwH6GgrAq/hUx+sckezCtu2+jvukgko8C4gQDOdMhu
Rgcpj+ygX8zzdMeTIsogf2W5gkEXCVnt5ry/wuPURXmb8/X3jp1JOEX2BAYY9aUEAVXxFj3c9qL3
2/x4rvnEaM6uZCQUC0Glj1kHerOWqR10HuTWmjpx4cS7JUjbj+ZsAa1dL5mYAxt7FNauH8Nk1bdj
w+us1T7E6jn3PrWD4Vq3vzQyTzMyNpKl4U9SPIHUs31/0qxAnbe2NKAHtI/WSt55yaSOBDK/YZV0
HQ6heE+SRI9S4EG3NnNskKnIsMWbVfy2RgG1ffoeJUkN0i5rhtGyIWlrsFYlXt56s7pr5BsYSzvp
5HW+yXv3WeAsq06DK7FWwyihX40jSo2XZAMblm160IYa9oM7XifwGbnGG+1sRhk+o1o9lD5icEdu
IblzOL5nnbeBcmCLkTbb6xW2xrs0C4vtnap449Iqnm18nzyR6Dyt7mYdGafHlzly/raw1o3tePSC
53EwOJhGNcoT4b5y004AdsoBFf0mb5dbSWI1VHsPNdx6KdX9SuAGtwLrErqXg/N4hWMf24S9aEzZ
PoKOz0qzP2VY88IdV0gQgiCeqcomkpdi/WIsmYKOZ/DlpCnbKcvJUfFG6OlmACpz3Kw1pHLiuIer
epfVAGvDNfbLilqvRQmlZ5E1yGTo28jLVU82jcN1x4/ANhFtn9CbpNFfmWIcys1UjhTq5bNX0IEx
iyZ3RciYNqsl5V8rWHXTnilfi2HS0ust1XAlDBga7bc1gJCbqPZXpdBQCjZANO8kVZ4joVHEhSeB
sYzZFSC739Nt/QmIan4RWRYhy4w5BnSxIC5c4wzhIcrEJOCitOIbw7g2ZLIRalf7ubAV7PYxZd4t
DkJrrFub3GONp1frUMVfrKSFGny3d6gBj86z42ktlN2QUef3MuQiR1nta6wwzGcxQ/GABrJOwew7
G1uOQOA/qKLXTvq4Qu5ILtpmXmVE/C9nDIXaiVJmzYnAD+idZBxKDpuBB0XiOVtZAlrV5GHVzBca
y740btLy4wXnXI0NkFirHrcGVzOPcgtk8GhDzMS7kWYAAZtEbIDaGakuorFexWns8bcw5QpBltIW
GIYXet3emCzQsfFx12pmnpsVm68X4G3G5fiwYv/nS+tcO9QC0QMVdMCSZHIkjGQ9KrE/jePWUcTx
s8zmWs3Uv0DaeSjfKFpw+SHuTsEtMkaBx44R0MI+6zt7xf9KdyAuG8tUyP2HFVqlRln07P/23tlw
Ze9XnKic69KBjgoBNKH4rmxlJG1CEbA/3veLHuXOOD79IwsNO2cseR8ls+cj5d2Tqg9aeJsrjYWz
8W3VnNphtATTKlBp+7chj3FQ5JjE+W4Ok7O+KZBL6/ZX8105ni+kho+7kcSOMQ3SADHq7l66Qe2Q
BMorxnFqmYanY4+c8SqcajCQI/NmaFhv8zubdTGpUlDhFP8icafYI4ub+w0hLICtNRdt7v0ro/+A
mIdGFCO7t1GsCR3q2iY8iy3vVuv5M8cktesXy6HPuKxRNkMEl9AfQF7rvHkCPTgs5u5y8eXWjfqG
d5ssIaSMDkLLGj/GWJLUW6ajIKJgPrO29BbIGgZ1bDDttpJpiDnrBwn45lJbii3pLhHCJVgUDKbv
TxGwiw5OF/8KapjRh2H5R0Sp2081/mQNquHLz7QS2tUqMPG9WziOgu+xiY0acFExKfru9HVWVqus
HNBKXab5QLiP/ND0J5nnD5FxYi0P5nlBouRB66+DfeSFuRHqc/Ef/0GdQboKQbFLlUBeGfK6j2mt
WLAGsSIkIJYQeWCLBG0/tPUEKaBOodyt3QWS61LPJQyLSNU7hIDspmzaL0bxlDi/HYU0IoHJ9yIQ
Qh7UBWqgVgY4Rq+cQabzQS/LQl+mXY8QZf47OW12SIIyWVk+dMaBE3APr2tst68cjuVpf0Uk+Kg7
jo8Hb1CMCkerro+Zu7EhNYLAj6OU//iadPRjHveg1RX/D5i0IyGXvD1pQFzyHt7qQ5LrjZnXprI3
wjD00rRHg1HBH2axm55KezM9XxCkhZI4v/4sbethxroGmRtD+Yi+icvgSf9p5kw65rdvufwneXZQ
cyt+xM1G185U2PzwyXM9UxgEd+vvqjMX1jYaFuKtGjpd024OGvhXcAczH3O61ujef4zUjGUstOj2
+fNrMg+A1KYQgkqMsLoO1aUGBxR+DB07aVtzJn/KU6UME3VGtSbmplyjdyxxHk/5tXswvhAJds2J
rqWsYZKAU5uNx0qxdOWNFiVoZh3yzBYorrCbVCql9XIFSyH/ywnl2P1sYRtL6+k8YOQjhOu9jmLY
Plqxf39W1H5u06sHY8AT4Pq2Erc+MsE5WeEGh5sQKAXimF1i8SX7VpbwMcRAKOWPwionGgDDoWlp
Iznvxv332u5odoCaVaXWIQzCstz2sM/OIA8LgHjg1OegosG8ci83Gp3X25MHFv1b2IrQOWbBpgnb
NEIBRfSbSiRS6mU/+u1I0AOFaG1RqCHtSmypXu5kvKtS+1WECzbpF4lvuv6R5zcq+HhsSjnSBztt
Z0iAeA6AF9WmqCn1v9kdwzjt6byfxr/oZRQBpwM/SqtL7ghguiPaVHOz1cpicq12zqnB8Mfari2t
DwaxbumXu2OEf7ztl067iaznnkEgp9vOrwtrw/rU2yTTNri0s4Lddm+yHryHymU1lBJw52jSDz/K
C9QauSiWE8/qVgxFpkjzp6/4cZK56W65VzcC/3+DHQp1nZ2RP5GyxJnLeWcA1xN4L/fJhgP4M5t7
1A+njlNKPk8cegEHOH6p5+Uo37GPSaeyrdlgnrZ3UKJVD2gN2ErjqNhXfh931k9vS+F0A1qoL5p1
jFvOnD8XOtOxm0s48gVaFhOu19M96j2N8ebM11zVb5qZ/RZeV06IcUrpDOFK5qp8UQKbI+ERJNue
auGtWTAbEXlIW+XGk1kHTx8jKHffa1ocJDV1XnYOGRokK+fKqQJvBdwWxQ8Tv8Z4IuW6ibthuDEk
aQwKveluW7XLw82tuNKcHLDkGBOcAhm+2Ypv8FXx+qzVffZxb/fMgntiIpQ86tQNo+KmcsAscUqQ
e1EE3DP6OFAl+zuwv51zGid2rjWAkyUDNh9+1C2OiqQkufwLbpsG9h2hoxFo4m9VBmstTct28EGo
K7MM/2nsJ5VVNZrzsDOWevs593HF/5rqEH3cHlgTDJjp3UwqpAFio98Q7I/Lrg8wNEJosRTUByAV
+jM0RJj2Mk/bfE9u+ENJyE9RmBV5Pn5jg8pd3qtgi//2XaQLff4POaEhhRNHCuTNa8QRHuD9hgly
Z6aDLeBXacQfosXHF7CSHdi7Dtk02/C1TTz6u/9XwDwLdR6F5CMu44sAbdSnFcF2xVwaYkxvH6ZH
92I9zNlcHHtNoJpHZnNhS13DjT/2QPXwpHUIKwOlrVgJGiXNEd9STHAaDcmX0aHG5jwUickX0ogs
h4uKsMhhsVgbxXjt45K3YwRb4ZdcGG5DqPf9KdxbyhwR5oX+pa2oQLhWBzR7xJ+nITgnAdNu11CX
d2u7Por3DWFNHOYZvTIYNnt1b6GOz0itsbHLu8TniAe6vqXAlBNAkxyGLXb5wouKtp1gDFgbyzWq
6M37t7rGhf6K9syrpS90/Ywe/lRtaSZ0Mxo/nKQd8Xjb35kKbneCnLVVQwJTvR6cQzrNCr4X7I6X
J/p/sFBRn47F2nIr3XjnUSK+RSPflLyJzuqqypMYXxO0ig5Xr6L1J0DWiKZ3QggISIM2E7mvWJkr
SYeRbNJuQhYZSMm/Kfb596d9bcRLeFiXQ/1gKS0QR58DW7axDgq311o7sFkpO9k79cbc9UYOBMAa
GMptREZ8cCPqU6QO6lNVPJcn2s2xOkU4CBYqE3sWvQJ9iscqGnAvobX/etPK12A2g3yC399+BJjc
TobGDttzJtWFoyj3ta8f9JwlS5Nu2zFgJtYVHb+UAvqacWD3MFTh7Zg9Z3rsOR/1eaNvuCXqOohG
Q5CkKFSRUpHroRFHafNokDWjcO8aLAtDWZCssI3olC+K/p6IcrbDL2NizpMybQNM4+VrtUorWhxg
8XyTGqmSA+2AO82d8zfw/cBAoaMIqavNegLCZ4WajM4JtyFyS0PY2yUHBMcydMmjpUn3RShbQnyj
MXZ6ni7x+/ez/8MBKXAsa9V+13HNQDVPlBNETtAb7rLhIP4ourRHceHgi9VeoONbjuaoBXGfHd6+
L7uMBirqq95d1XVPiLul/9GRu9LMhd8ocf95B5pToFhVTLdNdxo5SsrYTGnjToVj55e5iJX0DUv0
Od+cZbygbi+5HPfkgASUjd3l5Oee4rxHgjNFN7mtuHNsXv1Xvss/B1Yrc50RAJuaCXX+ajC7Opmk
b0OiQ0dpPnTDhjWmql44ED54U6okPJHV8gkiZc2qJP3jSSGAXku3JaSmaG+ATlnmX9R2IlasLkyQ
fkjyf17f3ierroBNOOj6+OKcPSMpH24aHw4eSnWjvMypqk8M7kZaCE5UL50gY9h/kCAFZGO6QL2i
ge9hhC+G967hEhKvYaISHGiskJFeASDgYCpmMcehk0T6j6Z6WcvXtlSlLMYMa0pKkSeO9mO8TAKh
mmYep7ur0M3HMygV5oAesI3+8+V0ND8CUeKbUs4xGUz7P9QFRm5Po2GkHgud/knC5fSbAr/XmWZI
Oc9E8pgmOQ/FnB2qnXCa+r9QJCsof/5xlKUMmC2EVIV+GvBhPLyw4tVu1Vw7UQmxZIzhTs5lMD5x
RJbNVXwkHVZ7LY+Wo7cH0d0L/RJOqAuFkrCWdhNldEyvDx8tIydQ87HmokoGFRSURcFt06aBulAy
qFvR9a5eWqElwejGrhcLK5Vocn6DzdmtuZux6M627F9iQ8o2U0QEWFJAuHNtYSGbbvcWc+FCGNUd
0wK6eWaD0pFk0Pn/O/AQ09McvKoZfWTw+Kh72DPtHYzT877L27it9V6MK0gLGzM/sM1Ebnll5lI4
MXcIRzfZxvBklkerylIdPgT8kkXCyXeeR1SwKKBCUdsChgnnE0Nyzvs536no/7bCkW1jSGVavg/m
JkdJaDd0eKFavYsGTQ/wpN69jG+eCOrAxlnY3+jPyRypmJetSFZBm9zP0+kVH7smjn0d4mqbqD8d
lgO3p9rrrWt9ohMraLZZbhvn3kSULk8PrJi1/T/LzWoVFGEYpY4M4LPZPrrqklhnSwJM8nqKdU1q
Z7TeT6GRK4ad/3EM4YzDddTnTwMVkcHdMTwLON/0QBVayvD28b3ULBAzoRrMlKQJvgHDkQ+W+FDJ
0sdLKv9MRZmP7ffQP+EnLZwSfMDiFHUSpBTpU1cdys92/HCxCMXb8JYe9EWiIHePG1QoC0XO0UzN
hQrCxgV4I8E7Bsm20JMrRcOXFLGgk74+szC8Em6TRwfAD33KCqmamLowGDkMBvk3X79ntZ50Bewz
QQBpAtr34xQTVA4yF5tMuoqUdMcSIqhPixCtnWnXIyCy1gtSihy+jqa9XPFbcRBMYaJYAT7Z7+sT
yGhXL5Cg+Jfy4uvFR9W4kj++2Ea2oYIy/EVcJ4NY+hJF07wCch9mPqVPkManzrjMj7qErPBHsoM2
ctPG+Hr7XD54mCpuAMvv8OYqGNqanC7ULAv+kYuMoQpbrttliMD8i8YMEIJUmFLosfrcMRROs8NE
q0/vb3xteN87RwzqU5qhlvG5QIcosTIhJSzNT7c2IhrLFKhuwuOxl387Xg4rhtiHXTqvEQQ3zV1J
djlgUCdwFhnItI7ht0ORE0/81vCDIcfA76VczCyFuLLc8BuAS+MRYWB5+QoT+FameLGOHtR06rc7
+l19QLn0Ew5vkqq1HsMBC0yy8Ow/KXcfSWg/941MnhezfasJwOq/QMtCbOHdWK2tV6oBILLC8pLo
F8BaArYEIIsuwliZgB7uXAcOr5Q03gZbgiHs9sHK/I42Nk1YJTT9T7rS3PJqbf6BIGGGc9ahdukI
kNCpGokiiTIqY56+VE88G1KkhAc2GpFUHuEqHPfV0vXiPjmV2OqBWaRZ1xmzucLozb2bxkR+wAXk
570q2gmDjbfGYcm1HC4lGDUGvbE0O8TshATs5P0EakuDIbFvfTLfA8F3pRLfzIuvMOK3VFbxF3Fb
1x8La0Fow9ajs5yJOY0wkdYVrD84KkHO53VpIkGeTUNMeHupiCaxfKGY+6nu2E+flNZKT1mph1sg
NcQrLjbV7cm4ABctUxyQMVtUPcyKRgX/mn8Mw3gqCzRQbnlDAMn57gJ1LIvKeefHVehkprh6uWAb
jlyKPChdgNsxAo8+fR3bCfvFZUUk3L6fcPGOYqwIyDl3RpcyDaTao0rGNmhMGGBojhLAtzkf6fo8
8Jt6WNGDo1qOIADAZwXCSHrKOr/z/SoEbP2BbTOVWv4GnFqvq6wQBoyWKJ6h8YfonNa8hX35xWgK
b67prbfbDMwSgVnYDWRiVehtwhRC5iEsxZSbZ7c3yconHbAta0XNBxV+HfUIJm0Cf3PrXetCJE2g
v2XDqMcJz5jQil2iGwaipxWJjNIXUjYz4aibh0C4KYR9ymzpONyklBFiJg1iQ4j2eiAduqf0uBGn
b6XcO+fQ+k6n2ttb31hanz4vaQrkEQQYxXgmr/TS3j4ctYIlH7kAGiN7rsQL5AmR4CwpvdNaJT7e
477tbK4LSZ28jNxtj0pR5RkHz9BFDn4aGA8uY+vTFCjvIbwkPq9ZKSwrckUkT0Exeibk1UGwWXkY
iN9aDbE6vZ9PxN+CIj3NO1/18vKxdVc/9rE9Qtwsq+j1p+iIj0S2wVITr6YmfzbVSbv9fP7KC/6a
n11iBakRo+XaQfS2lio2+LIjow1qfCjCK3Ybs+wOQxzqBDfWee3xtPZucMSbaxqKwWimWlK9fr8V
uGvYLvwCprXiyVWnfnCIMokhDzpnwBNIGM6Wv1G4NvnFJd1YJna+WBg1/MCH5iahhSTEyK/NU27g
3B5DxoWQp2jWxPA6A3ewjP6wcLo2WKxcSe4HE4LUKcbmxQYiGOfLiwaDkBxk5RXdv0qv93IYlQqa
xV7Jn9MDA+m7MNi8DmqwJrh4RKDcg7Jlm+eRJlTn99ptBJf0kIHp4ohh2irFCdEF+y2kG3F48jH2
zfuFqB1lGkFtTCEZ50ihPLBT+OLXzUYJVFVre4PjHj5P6CFCmK7catk6wmRbX0vjDdX0MkQM2P5d
9HZCuSGmWzsjNfw5YrAE954hTAFFkyMV/KLfnIzu1I0+jxHeKqUUbxRF29AI1nBCaKOSkreuDmEK
sqYCbp0hg9gbSaxXpnAbLMK5J1fh9enhy0yxYxXeGnEbOUNlOJQysSfOmuG0v07pa7i4fakah58m
AlF4zs3tk4Yfu/kfwQgOVTkkWQTkjAU6rJQFIT7R6mBThVtaF5FTWnUoo7JhCAh5v92TNIYs6y93
1XJma9TPDhodGGtb9FeLv+VV7d+FQQMpyosYM58S5CbeFtYxTg5iYA2nvBKiInj3wBoS5IPMmSgu
HAl6EO+pKhWg0W0rRWJMfmKXlKoDfw5ysocUEM0bKq2V2w0BNY7guBfb6w6dRWW7yc5o67A/88QP
1KaRu+C6VzEGHS5ehzPJ5DirieRfNChtjdTUDwWc/vjMLuFRgtiUZEvSHbADu3GfsOXUwLfcHQGn
eFlHyHPXopxCMwIreE5goRLN/nkj/V3KTg0L63g/xAwTLOHAj+usG8XesC+MtCk/tr3j39bw+EiQ
2KTYYGtkRO+unAo6rC6EZdQhy0s42KY95KrD3zQUmHelpBY1hwmbKzfQPqzQs82PuXXFu+HTzIhb
DBWGFNsMwPVT4H6onG4l94bEBzsJOW602KK6QnZK6Y8Saw1PMrDP0gFCJ1kxkbz2ajMf3ci2uQx2
/qERYxL36pTm5Hl140LANq3NRfPYAZlsxxvAxhPeN60IoyRsEwMmYJ1ti9/9kHuALQkVnRIU9t09
73AJBL2/Qy78VidSXa1Pagt7g6k4CqMFwS7j38bZr1WHR7s7sOzduZrI5CQPeT6dRMsleTLuArSQ
pT4iQkVUvoZw4fBHFjlWkri6yDhgRJ385g5D9wJXifItDngSp4Vh/pxJMbXlnMsW4lVgxi8CH0R7
pmKqaoTUL9nlayOlN+nBmxeuBZSMrfQJ4hhq98TJ2HI4fsBiGzwXayOaR6n0oq7F7i57cURUC+6o
EYok7jAsLN183AJ5lw1EQ/sfy2mbPvQgarrI5/omUcFDpCaO+5Mr+IcU+YuVYQtV5/VukKtzJ+iy
b4VJu5mG+ycKp/Qs9COpDk4IbzZ+ETiEauEBP20x62OL1kM+LOstYYD8T8apw5iH18ssjdJ1Wx3H
4B9KkDL478JlbzxfasKxwe41BaVCs6nY9pvxA2ItP6zAWj5dSvUbPbJS/AqW3WSxj6p/wcr5wJC9
DbTAJHFAHYntcTXTLu3bVjSDOUQK+lgGbpqIIa23K43jXmWpfCgomHHylBq1QShWyejHRnpG2lw2
I1fbqVseYPZ3Z/rchwGApqyA15sbZdK+8F1OjbLZh58MziKNaa3e7cHVMEFugZN/JYQgEvRF9kpu
SszSzMsdX0LYQQGWvm8NLDDzTkcy7MmYPK0PY1ZRRsbfIGYlkrNNrF5Nk5CpHpB0AjCN9+wUpYiY
CQHpD3KxutOw3/poZs172b7ExKCw64k2S9q1ShPoX9L/UUZGO6e36ruCY7H+3/A96sChp12alOB7
RdkzlOLPka6a8EhDIHs6vE06rDpCRK+DTCMJ+7xq4DJTD1ciTanKScVYrfF++VKP85j2lIzNs6uH
1PNWmNBGgKJSTesIwB86TYmEjJ4X+73Q8ndPyHD85iKz5wtudUI4BTyWJp6jOeIAblmA8CrC76PO
e8hwKMnSsDX96G3ZnQpkVb9NyTbMsNyVhlSdDR4+EmZ5pv4O5Yk96FF4STehO5uXDYhgLCcWZ5ze
SmtNXqoT0xIqulodNwqg2/073vLEG9OOBXPNVABQifx6HOhJXl9963htH5ObQlQtZirbvngwbegt
DiS3yi+ALLZryfE/u0e+znStdYdwmUpMu4CPQaSN6EYKG3XFclRD2QECtOEMVRcyr3XyAKLiE6kL
bPjcthuy8iQc3Eav2gC8R0OfS6kLO0JtkJHqQE9E30xBs8pQZpza9l8om+MyfANngaBuke4Vtc9O
rW+Bu0U/lB6xNigzLQ1Yu9/AK6pgZ08VlFp4B3FLSJRtLFje3vyMYA/ThbAI62rNXTq3P2t6oU3D
ruzCvAISWcF7tjV3IWe0dWg4w0ZWSW3rKiv2Nc3KqTrgzRzZkJ5/X43ayKJfEVQaePnvtyTjnRs2
eQgWIXylaL5tZwGbCkD1VtiWL7rrHH6YdOg0OXAP475tJfYMqWWSIIwHjYIM6N98XvtLwxH+b0kG
/bxq73VGsxEzmIdE9dTAkz9BGFnrEVyg+m4y/WykSOGsFnoFobRazX9EofMxrOp/E3T85KsDzyxb
u5x9WL/uY4KyE2sKPrvMCvwl62Q/tu/hiIXVQnbenwlWhtt6eZU1phYV5iW/bEnQeLrDx2y38/Zs
/iITfOgyfdo2rqQey/7y0BKBgE2N/OVU+iArXnv67qV7tZZ4mTrtCS+VnjKE/6n4TEBrNV5/piwz
RdYXcCoIRlvTKFDLLCYLPxePm8GxHhPf5ltVPHvlFzG0yY5bLtCuD16vCL9HadL7t6hHdvO6WTOf
iKTZG5fpb9m7AUjKDkRmfBGZAhuj/63Jd80nodDkpMHP/X6yNW8BcYQgYbuBQCLLcbaorJd4p4z7
gfi2US9FVGCAPHLeFA9s02acn8rPS2tLtt2VKfq8b2pg7lwNdp/o+FOM0iO4Y0B88r79oWGOo8HL
SGCV8jttQ8agF0xjbacCZgB9tGbeHF0Oacn5AaLLO1hwfdyCpv63xDSOb6gd7LIUyb0NL5KHN8jG
Cw0Myqxy6Vr3r7J58SEpHVkiJEfRD37HyNhlljXuqqsj20L0lwjcT2cEXyFzHSuOuEnuETeqIyb4
DE749zy4vkp+moySGQ+BEy/V2d5CghuzZzjF5qOAG9N5tZMvT52A593rLkjAw2OScxg9fssrQKOa
psQXfWC2L7DLapgohVJae3/pNqYLOo2rFtrncJ3QubF1DznOAIlFtzlDP3n4AtCHJlxAMR1OrElW
oRixdNan/m4NKcNDeVsM/Z6omCPbTkP1RQznEp80pta6xgSV4OpLr6xLY56UF/I/lsvdQTix9TDA
ubANxkMOmpZwBluxxh6QG3P5wQNCffbDA7XW5NSNPtEfLELznDZ/DBnxeBQNeKEuaSv9Td1Mx/Af
aPGGuUmt0yaOTAELQNmeaoTDG3h9xSdniXpgLvbqXxD6I5rkNfGK3dxgOWcOBcZT3fgGTi62ocPE
11XoTzQcPrpDH6+GcFKEvYMGbEkqHVNWSArV9kSE9drSobaoMI3y2GoYGyrvtjIhddT8hDeT5dxL
+FvLGTB2pf0HJNRRjNBmI+w6bA3hCFFqthBhcLnTA4OBF6YyHAFCfvHEv5SP04GuoumY4QWQc5jE
5xKgFJxasEHTA02+pDAp+kzbHZkA1jToqFVyvpxLgrmHFmA9uvg5429b7aPsQCvHzQ4p9Wea1g2H
YpOqV++5dLeA5DTZMLTjpoCOhayFqxhxBkAV3Jpq0XGuT1A7eg6KOczDW/1990idVi1NiaeYGWjR
ASG7CRt1qa0A8S58fyny1MF9f7dlufchlIbcjN1vVIMxVQQ1685qUxFkCRHfRgg4Nw8EpvI2o9iu
ebnzuyy+Gtkj9hFg66hA3+CMjRtkIovl7uYROiqHOEQPrkQtdacvZTH1Wh7h93y9bKk3bo/H3hzO
iY/75jG2K459hh407TGgSJx6YY4m/qjU30wIeSekQglEvHBX/L5y9hxfPbH/mGXvpqF7CpPYnN8Z
AAWH7SLX6D3ZcIGiBGwnWaNQhbjlyjgVDehllTDtiUzqlYx5Det1tXwm82n90oaPQ22UBXC0BlJZ
x0lhVdalwSOF481tiVpztNQk2AXz00R3QYooZbTVh3/Sxv4IS0SgqrPpfTzbH7WI9C06gSDTTSlk
VOeuHDKxVWm6JsA1dLtZRlOlj7dLQxPnZdz1ZRWRwO8SX7SJqHBzVZMxKqANtCYh1jpZpc/3YI1Q
jLpEggpy8RJ2CKna16PnVPsUmVdOCP3ndrYvDGOmHugP2e1wjWS02mlmtbubTfqsnFE7clY0pHQH
6mdH8Th6rd5gwbwpddmHquzpGoXh6ITQlzcdt73l7IUhYQwg6QB1Ape74IuxviC2iClPR/cCEi2s
cLFp20cfDW1+QbZ4s3JZnjWMIyncMf/u2qnSa1N5cZnvE6iigaterqfb8IGRGKyjUT2GvSpcH8Sj
+w/dcuAR5zOgO627ue4JVxflthQNOGH30I41jQLZ09+Go5Af+mDZ5GdfrPhLnuP7lHU34BksBcEj
AlHQAFzppnh2Uce3luN18IJDtZxHSn1r50wlSLS9PrXvrw/pIGsAhWosndnH/t4rXQ5dB4FSUNtN
r52TfCEXPjDLi85UfOkBx6poh1jmZdGnJVe0+hAO6weHGKQkI8cvC+haSn+kGAig0tABlkbHQSTZ
DwFt8vuG0GobzO/cyPRBFxkjSdTnEeY2WXgKeMmoZTSEMLbLT5byAbj87rHa3BSufNuMmhSynxXL
Sw9sQM/RrX3k7J0IGumrxNOiClHHs6Jr4KRi2pnsPJqKG8UgDbXNymexyeB71FTVrWG78IHmuV3Q
NVfczca8SWSJ1KBKF27dV/tU7HcM/0Fo4BjE1YREZ4O1lk2oZXCmxkY7PDlV5m/zg5ET1lnmB6b0
24ky5JkbRv+2zMBVFujeLEs0Cfwz8HE02/pysSFEMgmO6oJh/GxBKD65yK0TSKEiiiV0ibBSmakf
2OSWj6SiTlj5xrZZ8p/ANEv8zd43tyoFkbsNf2cKP3Xu8r70ynW1WWRcBwDpV0wKkoL3h0u7FZK3
PXoGS6BriFyguzoji8AX+MbKkDnnMaV9rlSBpwtx3zvn0zO/8i+A5PyPc9UKrESwyjvTqBTEaXXl
aqK6jXYhHBzihBrCdKNX3ucezIZ2+PnbfrbakJgyJ0lEpNPj1x6+Xtg5eTc3vdfA0mhdQ3uNX1V2
Mjm4/zDbsaFsN/E/TAWwaVaJYoWeF8930DS69hwIyv1emm7JIYTzxd+2n9nHLxB8EQVioOiq70nU
sKBiG+U4YKHfhL9OdZoIxYJQUTHGlpKqybukdiBfLUS18+vqjGeWDcg6PkfY20mlVAbD9fm2GJOB
cATl7rm/F9chK3QTR6gIiXoOy8+Sd6e6PRiTyibKknppMy+8BNM6dwGea/IbUHc3X87nkk6Horjo
Uei6ayzF4BNDuXM8W8t+xPdPhk5t7VQyWSCdf++BaazKmnoDlGAMqaNm/FnIio3+NGNMpyDe7xRX
b6l0/yo5yi7dRa58euWo4IJSH0NkynbZDzxvGr4nUtuEQg65stLWn34J4PfjIZd9/w1PVhzSuPhb
UUsoEvE5bhSs1HHPpEZuWaAygTHSDDIK17274xaRzPdop5g8m0suYXqxgO1TZcB8E1GKm8E67hlN
iJcki3uaSUhff1H7XGBJmD7PUo4Q3XjuSOURkRs1Cl3xifSycVM3XsPzhUqApYwo7DOPyfu+NiaD
iB8YN8/XdGpjv8xtRTixm16VYSF7YO22iZFw7OfZRkIcUhqBtwwiDDsUts5C7Pv8nHZ3ljJph02e
gFFJ9K9OF/fvj4ionHYGcIJ2i9wTFD1by9MMk9JUeT6ADS2iljjPm/ralQViTnmNSqS5DlwDi/gZ
j9NV7DiicOOlIhHuSY70E8W8wMLi5r4EdckoFlTi4HLCdTGTSUnPrMLmVnbXcFp9IesKaj7Jbxeb
1mpAFvpjt0kL1kzEwtLp5liafZV/pFnVISpchPU9P6JsL5isohg6JQaiZO+kqkp41iWYOW5iCVe9
eYKT3xP3QenNbrqFK9o5xj4+fAj5BcTReNfT2xP6nQE0Ib5/f0mBUqXu+JNFQMMK6nfCaqCZQqk5
UIwv0QRugyoDi5eHw2VLXi9kjdu0E5ELLKUjk6gqyNKbj85LcEfYQlQXP3jkNoGmYyEn2izu8Egc
o2de9t+8Btd7NivFd97SkNyEUF4EQcIWOVuQqnI3Pni6dGjfSXRX3Cazavm9pQoCXd/QH4TdQoc/
/KsAXeUM8izcl+kD/Fbj2BYcCNy5A+1xhLaFMn/ng3cVtEhxtliWNzp4tJ3YHj9GVxs8hOUfoK+l
CpYK0+U060G+KSqgLVFdo26ArMoepSnJRHmZsq22pU4QNDPmWA6mf3uhmKIljH7INtM+/E6Ywqew
IJl1PslwZJNw/4UjW9jS02vDfcfgkshYFZ6MRUGAU8o6xX/CmR0Kb1mX0KZB0o0OwBGUfsZelOQu
YswGgMKy3gD2RDWuahu2MzfStgzt/+OqTaHlg8ZWrDmbxugs6BiLaMoxWqk9IOISvYXCb+FJaqFQ
0/MNJEEJ/QZVIFRuSqhCmaTFd+cdehaHNwQP7m58CMYDGPai/D2VdvvsEJfP9tiXSZG3a+8t5jWL
V1Rle0WMdHS9DEqu12iprfGY9NVKd7E2gTCNTM21qK/5ZQaecSPC685Hnov9ibiuvK9Fy6/6lzkc
I+HOrplC+hZFBxyKQrNJUzQpEhv6j78Pk6eNMCiWANwTBncEHkslA/Va10bZywzc021D6bSUAESp
WLqpn0S5GU2BZDriiAH1/D8YMLGDvPYGw9NtHlmI2Agj0UO6MaDij38ySksnxf4mCjjEfFyy8fGZ
/rAh6Hrz41Yrg93GPWtiKdZ5+nwx2ap82clYLRoA4TGxl8kNJT9NP9QSs6zixca4IdlDqDpQXCQD
OWeOZmKVIr8rV8EmaDKYzlnioW99RMlfc4DpUC3rUw8n0nGfbodoYs5xJLKAVCtAN4TSpaHxOqvT
YKCIU2/guKyA8euxcoEq/Rm43Kpc2ZxFDq33zSqQjr6Yva0rK4I1uCnGIW/ZYxCdRsPvamE7EBVR
OLOdj5YDHBp6+PKc0iAszxavSnA7slHsxr+2H+BvAqdQeFzvamblYWrgW/0AiNv4Psu0TAnW9otI
WBceLRptqSrm2qFaC+6gNeO++IQN96QjqdR74XkEEG6lXtUvS/ZEJgeWOSMueOx0z+YuYsrKi4WJ
r4Wi60ltsYjPq1WUH/hZaP3HcOSrIcInIMtaNuujvV+sPrjeZXOrkGDFZXMiZNZjM2NbjutBM+UJ
w4bjuFM4hgamlPdWnkYXsZt5lkgHfFb70rszNS2EmtY/9ImTXnK9yVXTk+SRQcheAfe96blIdrGJ
nS9Mm+sQQWlbVBevsz6Hrf/2BaY+JAKxUkl0BmQbMQjX75XifVPWF94r+cgORMpQV+044rZHUiNB
gETCEvXnXS3EJMWPwxdSTTnc7XdfzMWRQ/UobpLg3gPxldCSmJOpv0cevCsmhOwVZuBpXAJA6Ekj
PubaT5Gny8bjFXyWJj20yojqu5U1M1U2VxqtyQ0y7ORm4aMrdNPA4lqRAxyT8/HmETC3VClvZ+Iv
DVGdozLBSCuULSa36bbJXpdGZyLHeYTiM72QRVxo47J0hgqibVkZz4VS2AdD6OR9pJbxTERpfyjs
wHXEESnGa6BSRdGKs747G9a4oG9ex80/urY8M58SDQyvQkuNnrQdtrrzJDh541q3/hfkUZWLa2sd
2yhhuZNcxSfiUVN/vXWsSD7fWcPv8rCRc6H3TCTuaRdogBGUHkHkvDbKpsNdFxzGyrOwRd4YVQsp
nJifCahudtX8sZlRQyDrdLmWj1BQ/SjbBRYfjnVEzqiqVp/lGd7sUXQQpjLmfeSoYce2YSyAbuRL
LdNP/rD5sXXAXB2fqBPRHKEFyAtwIsGSKx4JvZXHiKtsW3YQFc5gJek8E9YqU7ccmfH8l6pWO7aE
kRKkDlTzpdQfeQyGckFTwP/hDFJiOb6MK+h090HJ78Pkx+3g++URjm8tkTseqzCKr0hYSBfTM6qC
sGkTzxU/fouBdrF3tE6kqwvSxynG9pE793R6iJQx+fwLJEeVpK2mjIHjP0WkHLxh+Cx2dhhbReDu
Twb5YScJHcrnHpBA+3fJ08SlVdR00XW+qUvZ/1hHzIPcSCu4cidZuPC8hvBORgP5Estn3B2Pz/64
TOnd0QzDLaPHadqQzh3jggLG4DCySxBDzjnG41/PCiJhCVQeNB0zu7I814ptvS8+tLTAec/A3YDP
ac4I9C31q0K1XZR3LRtjq1LD4FXC1hHIgB4lTF1tgV36q+4gvUKTbvLhFiHuCr6VLG6yAcwcIYF8
rcV/poZB6dFARMyjkHiOLI6N2n1Txag+7ugd1NOyRLjnhpuiY6wOIvXwKTDn/1iXCiTvd6XMzVkO
c7M1qxsFFOw0F7vIGuomPdQnf615Glxygkk7A4jjvBYuB0I8hlmdcvUixIc93mRw+QWZWHpAh0AR
S2qRlwPLpPCtzz81Aio3EHD6I5AWodPc6U9GbunLerTDi442bB0Jws6vkaQT+jnQ7gJDnUGShFtH
fCHExDUE0j/FYkSfY5qTevYYYSWHIkIn4e7gYGSxYNON29s35/UxMz+1QC6+xabxuYDT1IZRtxIR
KPCND2XaQJMOCaXZDVqfQvMMx2yTaUkNAkStn+ouCUBzeY/1DCycGQxexKsCqIKWvn8x9F2fyDO2
l1WLWyD36WpzT7aoFyME9vEZXd/YQTIpw6AzJf9UcUS5gh/nb6b0BdGRw/RPjA9cZab+dmGLKNOK
+ltcV+qTfolqD5mpbDxRtTdxZj+EX85WbJMXMDnfvdRIW7/Lrc7zRjoA9Hotii+rRED21HKa49mq
rpx7l3Yl/Ps2nGPJcukCxEVz1/OCq0jpFDhUmMYbvA5Mh0AAhR3EL/YeZOj0/2H7So7+yKW685XL
wDhwMA6esB4RoOrYkwicLN6HXGJvGy1vRjsUmxJH6F1qqxfR/gpukPHmHnW5fj6lf1sP9hqVBNVB
c+8lfb8Q0ZvCcaTlm4GIZy1dGpgmBpwYhTjmHoNd1fYINdVv3dsYN6Y3fS1CiykkskC7UtfwMSHP
3XjVWMMU+v1MU+7wU0tGL9oQGngu3VbbbcIHd3nWahJrKLJHE5c7yDnqQEHEthgBBOEkI6ptHdk/
LbYfY4VFbYujrCQwrkg1fm5K0nWa9KtIdlKEiw4D3gnabTMX6qP+5KcvsxyrKQtOWOKyXijxinuz
0tYd+CeO56cQEcWuy/IcawQgDoh5nrqHCCmSiCoLFqDt8kof9S9znSkwjWRSLh2+6YW7bEWhPEQ8
gEczbp6im4HES9z5UT3Qrkoy1iffPh0Yy4CraOFo+pR1rai5UlHb8HtvndkZpw4U6g1QIlx8TMd1
7904+Vl+EFjeKlGcB4Yr4bpPKOjUcUpv5BRgJxQbRyzELmLEqxv2QOlom2veJFXJ7R2V8NBfDOZp
zWDeoVHqNy89WyCKP0k2SK+HPUO0ldUsj+SDYkhnWIv9lLiph8svL/jH34P01QwkcWRcNYVSpJW7
IpRwkzhF+DfJWRCcHO64vCw+J5qTGDpWyMvca3Zz1oRqRoHoPQ3pewIpZ3t0/iTb6PNgQnsjRcXq
wCGixZnOfUPLYDloCfbEYKNixmFExZxtsPkuv/szAoOFi4jV5vtX78NqBlHIZtypYpkr38xb/fPK
4ZMdTJStZYK3UFdE/3lk7k57fmOxGyTJmd+odeQq15TazQ9P4PUNT2eMrbkdyC6EZMIK6Yn0plep
iTMWHCtxQos3YLMhi8HUj4275pCTPNvw9pp1TYlSN42fA7DaHllXzMtpQukEJNfDtcuofEcIKfBC
fRqsKCE2kjnhPSnOb6zkRg5P5XiZKZK9oMFqath+sLU2mH6ylpQaL3ydXS75n8UrJsvPLm1iEO94
Yi2jcanTiejSNPuiVZ1lS2rDY6ShXV7YHudOxl6zioVwSl5QKPSh+qF+Dk9/XyFauLfORooZbEZZ
OeRRyYN1zW+/TKAfJvY73HEQOpTztCX4lTwawtgodmwkSSQYZp3yDxpc4FhKfIYU0RmT/xZYNNqC
QnF+6T7mY28O3gmW+VIze9DUhxUnWuHEy+8BxC3DnNjdVcK2Ae2ZS341R/gdNGqhBuLh3WVomlua
0HbevsBbtkWdinlQu0hJuUBDUnvZhfYShzVDNJb6+W8fO50mO+CrW8/CJRooHYrgQoPYIJiHBkwo
xmtBE5/KvkifGHRSgEmHobHPzOjhq2kKA4FJnbVUEG2LSNP8im3SK98NnzoGPJJXTiAeViyamWGU
hERHuIbGYqAY6c/C4Fd6Gg+RAF8SGxC1awxvc7wYSW0wKnimzGCaQKSnoS/slC+OLP5g435lyDH0
7d8mPprcXm0PQcdHLRmmF5R/kmoAslSERRVNMpVt7/d5gg48Hw07pOf/Qvdx746NPA6V/VTK94gb
xHhyQHVb7JQZq/IIuPfVtQxW8+7LBdsA9fXKvqXGLT/6ckh6ZYqthXrWsuydfJgdbiagG5EA+xIm
ZsZivlhyu1n18Aq7J7TMVy6ZdiWP+coBO1IywU3nSTR4BUEaBCADMoanC5vFO9WyEN6MwaOmciy3
flt6JPv5TgJR5VJu4U+sL9UVKYh93hqey4/tEbwsWLDWyw6IGMSozGJmW1qUlAojpqCKXBn8P6eV
e1qUP7AOEdenDtuquwYzgVHj9mfSPA8VB0P+JREl3sg4zZZ2FCnh06VjXM57dOEgXjkfS628FuoC
DMWb/oBCc7S7mpk9lRy33RpETN/TBIQy157bFO3k8uzK1rZI93oPnyxoeIPkAN+oFX9Sy318uEPh
Y6XKIB+ht9CN4Q6mnW+EfNzQBNz4vMuq7PlWrcBbxIpzJX4td8/JqWcdHPN92+QUFopjvWrxfHmS
uhg/VYBPINNmqqj+lSIqMMCbXIF9I4nkv40dl6yyH6X4mTc+6B9EYadrp/0IzjuxJWv82LXnlyuf
fLGzfzI/3FJ6Tfd1v4FNPj8oouAnfGPeRYKizgZqsrU6kRejf+jwFQpvD7VmaQROJCUr59q1Jgyq
WxEX4doEO2A10H52DODWGz3Xf7rqxyzr/EfNrY3RzndcMKlgqfvpiRjtHAZEVgO3b+jEU8hkIzGZ
3BvVbG1P16rNBUmMkRkujRfy3HYeXkk9r4tSK9Irj5Vit5rAmSG3EqO2vUSHRyfRzBvM+dZecyIY
rGpN963OetO5GqnDp0FRIhPuoH1VKZXthe1OvM8rek5e0xBC0ic1QT+cJznVI9I9vNegCwtaeJ/R
UHEPZ7/fTvD/okl/1uuDSE33sH/NEoebhwktdA2D92CI9s8+mCxuyJY32LZAX1+ffOBnpu/sCasp
qTmiL4b0CZyo2pTCZyWohvpilwAZDsoxcLKfv0UOXfLLAKkq/JrzxttW1x1o2QBpFo37iFwwxolR
NNkt4nrhsWSQBLfCt2eF+gZAnFHZpPbv/jbHpFE2KV/Egp0JnScrWenYXDANGV/ldvS9OSC2ULkt
fJw+4kqss9nUZKyXH6ygKAYsFBHJfFoQhnIKYNNk4ygRofbM3bYqs26uP5O+C1Bt0RtcCCY2zaoT
778IwLhZyLXveQ/Ni5w39zntoTND6GjMVal1OGsPjPkzxzB0Oyq8Wp7F3NZRGSjlHuYtCyJHrjFo
Ad26puu8NpdiemmKgYYmGeR2GFpNtBVVHX23MUEJwdVw6X7YPJBbPWF5VYC9WDzDxHdhfN9JRQ9A
FUbLVlEXHAKfubGH7A439FQgVeiCFNYUZjrD9vQTPSpXRaZ7r+hnJw3ZYWWwjD2R+VlGYP8LUlO3
HfmYUneRVP/jNrCC3YINxzt5PmERR2c2KaxFjVGNNMTOrTu9iPa9ih8+dNupMypOTvZT9WUUSbUq
HFve93sNkQM/eA1oKmsXR4f9kqbtk6qM/C2rbN4t3oB7YrAY6LqR8E7Yxxfc1e9lRLNoX3T4sRol
Hy7Zcaaww8ZHSOyGXyESowyDkCIVGOC3jsx1D+EggP7s7LvPMumJXkw6TR9aTK0yYuB8megA4N97
2Ksga/mN2BdIaSqLTpKkrZ7IAi02XeBX3N+yumbcvliIZ2bEa2BBmfHGl6DzuScCNoMdx6Dq06Ch
8TOG9YlGahbS2PvjB91j9xQczzqxF7gCvSh0pP67cDO8hGNd7jbzf0Qtz4K0GDpmGNwzhxHzqIkT
9HK2z9IM2yjNL6YX2YSuBXgHnyXnCExrYCwykE2qD+ezdhuOMfKvfqQHDsIs3PByfQXgXhPmiVh3
vPfbc9U6pXNQvVqArCYvqpT/iFrd8gznd1ggvVlKGvdeT9SYPv/fr/1JkV/VN7P9ytj17pD90jRI
nlE9R1+ArwUwo1mZptROmkCh4xMNIVTSaElhdYqNzRlIX1GH/hFf83PRf2tN5GIVOIytSaWs2Vpf
eMt9/AFY7lE02i3bfgiPSbXvP4fjBUPvI4WYnDYfyejFg+tuvabfAJVPdPpjqXvsmU3A6hLMgUan
Tm5Yhjvre2qBw5DxhDnWxTwCvUWiSFNDTi7iTwxtk3rBHbbcENYimr7nTzJfGd/waJVTkzGwS4JT
9D7SM1e/pQDOwxc2QUAHuuyzo5JSBGyPHOwh3ikJqBehyi76pvDJ6RJvggKmuUlBOE39wewsW8Fq
I4y8a9A8q5uCIwMO5O3YEpTQvHVB88xDdxAHBrYHrUy5laPAungcxulG+FcaviTvxtvfqKA9ATsn
up/h92kkUuRNkb4GYpXESspcKh+snnVXZR0+neNgyID047P9mqGbsRnaTre+8cOeFoZtoHHHsckl
TSbYjBQMHPSUTgaipAy5kZpHzoUA7Or0geqKdrHCMuOePwZkkR1DlL9vHSf7+PeFtB/9Hpo+isrz
FB+yPeLVO3MvdbLvV05HvqL5vFt/Vj+lJL50lzNMGTnZ1NweeEco4d4MeGaaPJCa06M1UHfv9eWm
IzO+YoHlhJcC5OlSkmHKqIKq/VPVOlKIZ9Vn0gipJaBP14mcGSCPFU2RfsNvprvWHxko4hYY6sE5
k+nUYFWGFyiFiTrdDMNtuAhVHdkJevFbOlvplwo9Z2pH8t3qQu7dJ0T1v5nOz5zHjmCYVJhs3G5Q
vVn2Hq7uDo6ZubSeKuVgtzx2HxxyjIyh+tzrKCq0ydn6bc9oA0kdPF5sAzZeITyhoPPRw66twTEb
EmMWbtguQbt9HP6NxRQeEObiIoMg0boPSLJEiO3xfn3YtMKFgX1TDmqImvk8nXy5kr9zCW3X/t5t
mAyxlGDhAlQ+6R2feZjtV8XJgkPXCD3RUGcGeCRzV1x80zwuLh+jrkVMCKTwpgmTYYJqefgoPZ8u
mIcpHBR0Raq8WuT2IEWsiJ4xX+WLLrDUgUVUHmAM7oWboPnGoNRVcblTrChKX8YMMPfLZDXzBL81
uWdm8D8kQW+oKTItv3JG2WZ5j1zrfXt1C2AMhTwuU+rNFhFeoo0kFolq6lD8X92FfVBvjJdnObDe
8UYRPnSGlHetmSYkmUv0BMzJytMkiAgBto3V7mlCK0V638X1Eknn3N8VR02yEkJXCJDHyHJM/wMl
pw00JTGXMsfUrSMJGUpJXZp4VmnOhX0JftHel8AQFIVWgYp8PsPLuTDTSs0luigYzxGNZN29uLSm
KIq4AJ0COs/BHWO26gv3L0hqw4pH4qq7ye6IkVRdrBrRkNMfgNj74BlYT87cJQ7ya7OY06ZfN0tJ
zroyyHYR7YMnLXaqgIyUaxwhs5gXyeyhwDug6ie9bvpT7wxMjaCBgAmyG+nAxT9enIsAsX/NsYFt
WfMXD8r26C7J9jvvtiQX80/in8qRCi1S+WZNoRPs+v2MsMHekgJXV9/dxYeg5om6LGmaxKTP4W+/
HxkYPoBMFSmZdjFSkiyHSYzOrcV2yPL7A1/E7GOlSfr8P0fAZhcphaxl1rXhDitJCNinxoY1Jm0D
PUJsLAT56e0p9PBFLZT/kffPa6mOcThDgaefms2bYmgd45e/LDwOGholgrv/uAHZoP+c3FMR55Oh
yFwnMmaQPyOlWYeAJNFzvM/E6egRytYdnZnO7+GhBJiWekKNMrl9JJj8gUzGuOyhoFx3+cAsimJ+
yAR61plJaJY1Dk7BVodPZYS/Hb/esAXBkCBjzI5VdPEuMGTW3+EtSOydqFK1/V6gFH1INXNV27Xf
bLAKM6NVi9zwIwQinHFzj8VY9j/rZDSXS/9tWoGSqHFg56nOi5+dzZ3sJuHok/dOz6IHMepvHXsT
AkSmFbQwq1dzGD3eWXmGsLFj4aM4gr6ovKrqLCm2k0WWRZYs1Xg/H74P016Fm0mF0gNvw9CJLWyv
U84FqMMUujE8gPrt/huus5imjgc90krIiQF7v4z/ntXtmyWiV4KY73q4FZHh6DBtNIBxQQg7ydaw
Pd66+8CYi4mn3AoPoppRQifMkDgaxZx6NCPUBG0AuFWuFizOERMy2gdSNBZ5xEnzaCz31NbagFzi
tBP8Q3sbqAV/qZ9nRw3gAMUIU9KCmv2E21hSgDXHQNEpbuJfoalXBDb+kf127MeXXuWHfwA5Rei4
U4Zwk5g7j9RtGQxChzfffWXdvm9CufCUaQZ+wkVfld60TtUsru00soqgptEYv+GCdQk8tpMPBzRT
2wbk3OJAYtVhmSyDbYl1SGNV9sxI1NQuJTA6SloUY09vaaI0O7QEGnv9ObLFwrybwH9lszG8xsyh
LLfmMft3IQeOJe5tAl1RUn4vfKgP3HSYmUvOLExG7FwlAWHYPGcWDboUChWzZwLy/RElzCs/xQj0
EhGfF0geMSwdaGiB1XExJCMKw3xCrjkDCSKZwQHXHaW+nJNGoIG6EGQeqiKXJwVTNkEIAWURU31K
0H4qpSSXtWy8AVjMlIdoiTaxGQeYDyOrBKorTHleczpHViPLMxp0ynsOoawHt2k7RqcJCibaW22S
QmOmf7GvcTvmCUkk21HIaAjKpIG7IhQBvHfoGocjg2PISP1EGmiR8juW3WnuJyUq5xYHexHfliyD
ecWCggC2GxtkTS/8ZxC8rEEq9i0rgq/Ku3Iu8hCGBAckMiIADqtN1kx6q/p1mxlKEdn0h2u0k9Dl
ZfJ98NF8H4ljntfKk1NfsSY5lOoCFiJMxpQddC9d5un761RwEZcGmiKIKhCKZOBZqkQSa1F+yR4e
GJoRGXSzIGxQBgRyM2FK46HEdZQ+4ZAPRdyWqwWx8k3cpMcMEMTvjPOEfRz5hl9/9ZOrau9nCPXF
Llq/0UQcnvQF25slq/QwqfL2IyWjoCIEs8opcIta6RLeLLgrQonQ5uwbWQRSndQVgyx3D6xvuTwX
G0rWlDf9uM8XTcOsD/gYjRw7ZfEy0zKmrQIteOY9lPejibSjSMRMYK98OyFUmB450IcY8S1RFbpL
5PYP0i0pv8nltrcGjW8p6RWbnq4sNIUny2IIpA7pXsfWEor4k31a5ojPXsqWz8BVaAzJdDW/jnSZ
2WM98WhQP+uS5/UlcfIusgQj1OVBt53RGDwT3fU1yIRKtcZ6g/Op46Ac0RYZFRigXnRMIyYUEsb4
QoJO8AMGYk4uDJGbUja0jCLM9sVdIaan4GD4nHZdM3F+okmmiwW4U10ZoYDK+WbNhEMU/5T43vcs
Y9YYhGi3V7Jimt7O5sTJ3bLp4qsX2/kAi+xvOc8XiDCcD/mhjilUPAC/8OxPxKNIEvuSE/eCQhiL
010ecw32F6fz/p2Fk0+ZjM7SX1X9e5ILwx2k18x3YfS86GJjU8ywoSWhiNfsK0+SpKzNjBFTvTeB
BofSpxRY3Hs2bqsJFo3UPXnvr3JRj1Y8S37o2huNTtR3gRyTPpfzJGIODalznVkbp1OEgDWvvxQs
YQTsAhdr8mLUwR95i3O3seR4xgAJePelqsiaQOFK9QSFMaYxrJw/cmPWFmIo5zuZo7DdSSiGZjAV
PHL0ubj6Mi/1pBctfZ+Wa1oqvJJraWj2l4U+HkzFLVOsmh1dT8BT8xaiCsdVPCRqze9cNLKHK8ia
npWlxFoVBXUMhmO9D/jZCwuK4ZAmQeCvb2HGDVNbcY0eqbt25GcFTCIcJNVlUUNcrCCAsZZ4hH50
R8wMQxCWUobYNNIPEKcZkYclh3nn/lemAAgbyIUR3lo1RFI0an1DiD+AGzbVGB5HyORLsA+5zysC
2pwgCKSUskYPW5dnMWBd5QbaYRtlf0kUrI5zFM5Xj9V3CKHpKk/MsJLyouWSL8I97Fq+yKg/IZUY
smojhgEDmPJ7O6gJJdXCZHHFvXYD1YYURlguCs9bN8/newZ9LHeo4IWJ92ezbVGTiIf9ssfZSL+t
tGeCY8RrLBpQl8y8Y55fOHHyIEjJG3lmYRIDggJ7VzDy+3wb265yEUsoyFOvQPX1IDXzSlxyn7oa
nR1XLxJBQ2t5gAOTm8+A3bTJIVR/97LiSosjLmaqP2dcHOXUpiDuGkkBjVuhTCcuVerfB0VVLe8p
SOyhng8PAadhFq2GTyNTKi9p6uQ1Hsj58Sszi/O229JrVdms4xBn08qSVr5+3PdU03PWEl+w3ksa
i3bgx5agH4rptz0zos69eCKmTgWj4929ONCixG8ThCHYljHz+vPDT76LkoSmKvrp2GFMJD6JpUOr
B/s7+yF1vnIyFnqSZ0WZG8oaiS3rqQi2EWA8CiaL/7KESv6+lcSMsM44LOu7c6cZ8NyY+D9lACTx
zQP+9AG4/ZACFPU6Oqqb3bGuA9N2OFZxYJZnj0XIdrP1TR5zhFgW7swrYVYJLMWvadX2aWM+gTER
2w3dO0oToPtpMkWwpYSgFNW1x8LQqINiv6t/V09BRo5tNH4Ipr28D0bZ81YpFYJogBe5N9uvix61
SpcPH6yom6/lLxXt1ngcjzCNvHhUA3krnU0U8UU8HZxaxCeQKocHJBhmpSulS4YD9je0GS975eV6
qcFm9WdASldhGg8PAtqDqI/2H04TZeN6sE9ar5IFmUgMm/UoFjs3/Vz8XC7w+K4oHJA93aUpYQwt
UDUjH6r6MoNFfB0yI51u32CZjbeVlVk7mba4BVO0MEVG4r60TaRDI+ti8hjTcLQBdJsnjv9veNn6
WbUVkBnIyjHuia08VE1tIBGsgR46O9Nvly+79DDo8vIUnvWOeRN0HwJz0w06VHs9XhxvQNDtZ3My
x0/vF/ZHqkShSnxYxRMm221+lz0Kf5t9Gv60/Zx8LwYCTqF/B8KmlXHUIAHuKtjktkhhA7VZlfEf
NF+lF2quxLg+Q2s7OBq4W0yZ6vB3t+Rbh4FwMu83xNoVxAi28VXbR/GQrO5XjLkLIv7iCdn0gfRu
jRSKthG5pYYAXQv3CN09PPYqYwQFG/bscj3ExqS9n7ZWG08Q14RHFQVBAQAdmiPoOHWcWIeDkNvL
1MHiso/kDH2hw5eWQsTgmyX2pEPtnu+sjQ1w6Q6fm6rmFIV52tHFGflma8dwU1R8gJbHIsFe46N3
MrUHpkrgwDImPYj8/Nx9h7ryCT1nUKXEK5MJCM+wgfvLFtzJeuiUOZgkLI5pkYUIVDZz420BM7HG
sXpqmX1fkMsTn+0RYSVVX5a0+4R/pnB/NtQD9epHsY0bQComhBbETLNNxV9fotIK74jBukCeqw9N
OwkznTXomdULa4fJBxMtVaqMj0TN5/2knm3JqOXnpWVKfMQJ2bY1H7RssyzFo0KOtTDx8waR8Dls
jGUfBctUvodip9xKvQ1ejTvrlm8SgmatxM88B5xPibX0vwnIe+AR16aW75xO/0BXQAqPf54qj061
DEepjZ6Sey0wUHoBwvc4t4BA8pRFw+lVHpFH2H9oEAitxUatMaxa35UXcTK7VFYpSLZ2NUrncqvO
jCzXG0qTi3XKsSj885eVuRD+cq4oSfGV8e5ba7+KBb7MQgmiKBfgMULJEMr7JetET+4myUqzzINF
icbxvWQXN8ilUuyFDlTbH+FwaGKvUaUE70fWLQmkIedhKcRVokBgLRCokjmxBFiOYUI5AY0ND4UN
6nUCoWLT0ote5LrDrH5Wr8OpooxKI4nzQcyDutDmCX85ajVy+96jdM7Eeq/2pKIMKGcqSjrAxrcw
46QmOY4MkS7h1unvqpG6AtisGMvRqKJQeolvUU9/fHG5O0PjnCNg23Sx03SzHarAyF+LE1+YwK69
RQTDoGPdk+SzPOVOWJkrc6O87K7pCIukpjSP21i9oR1bLCO30BoRUpTK1np+3FkuUKRkrf0RNt02
7uZELTHCvrlcIPTFEKBNn30vW1Q4l7o2Roh9rNmeNjBLlrJwc8+RHTDgq8dbhn5Z6E180J9VXh+I
uxeAaPldv11WzEO4rbZeOyPZg0bA/VWL42G6q1dVVe9HF3uy8oK0SX0GrhtKe1hgfGWBsOXy50BR
Hg6YkwZhPYPqZvEuFVbc9aaq6H0KlMYm5cB76qqlJPr2Z7RR600eyipeJJNJdrvhWiFvtwtJ4Df/
yJCjxVlG+hWfrA3t9G5X7LsDUpUMg+dU3vu1bRW7jkpw4VnxPErx8MDCCs+CjEAzcwXOS3Ycod77
qSl6ueWH40l8IrS+pt/oLwgx50tTnCPc2mOK2EpX7MMYegU8978IhDzphz/DjaFiRTZpilr9E4J2
FCMOOTwK+ZOTjQLpY8LSxDMxj/19O8JpoHtTmZbxJw9gMySXn+gt4ZTxz9NKsh6DzjnAAn3PuVR1
O28fKhzLCXSozkz4bXj3Usurs4e1qqRUBVrZ3lNCgAqh6e7PWUvN+9fTTVhdJcCueHHeiuBd9T7c
IkrOZsTKumQyp/j0//wI/vz2TNrGjhOeKTkY1fcn1lHdUEmCP0DGWvXRwEsHskFY3wrlGr2phw0W
nA1M1qA3+Ygof83kQGqzwbbvkHjp/Q2XwCnx4ggin9Lj4s1LWlP5pPwK97geoymFxve3xxaCXUDi
3mtLayPP9wKWi8Ms4DYA2/7nIb8vUxPKApHZEAk3dC35jENuclplcILP0Z8/9gqH8AxxfYk2kIYX
lwEFy74FS2elCUzp1I7cJ4RFlmaRbW0r+GwgkloFetixGEhDoUXKfQObATO8eSSzT+iJsqTphqQY
0j8Amouh51SxFzXn2oqZY7RNtK2/MPk7c8daW5pih+jEmKFDp5iAf2Pz7DpmXF7VToYKuCjBMyVA
UklLtjPYf/4EYqkB1RUHMpVNRwCJa0S1Ocw12FGHb4JPtCWBUc0ozEY1fOTvjsObM7DWuZPrLaRI
cXvMdRkuYLI/0yjPTcQ/xcdriCtyoTfPlJVjELblYxLRYPAW4dCn3/14Fv4iT4xTOFG4C3yOg/gT
UB/yyNRs8Bt0Mcdx9y/AmUO00k2U8pTD/BP1Ba/+dsHlXvbKAv9SBi5Qx327JZXAOnC324gzImdT
DxA0NH3KHLyjmydGZ1u0tgh3/xhStn3dzeGZAvcrpe1E/sXwb7O8d5XSMgMNlA7W8lWURnYvx+mZ
aSyT9HojOJZVZp+phClOzcPv6lfj81xIAnTe8Xp845lh3uUddP1GgazfP/c+9OfXknKisb7cp9jL
7JhmUTJjXEdBwV2I+1pccrVgSaJGkCp1oJixYAv94x1bnAbklC45S6QfnAgaYlkY50yo01RInZFE
2zPm3Ku6/wB9GdPZHj9idEtwaU34ALKorC9u59fKr4nDAvo9ZAfUnW9I148vZhvekHd1UPxjaIVN
l5GIbnyCFrOZGRCURre4UriDDKrNyw3613gCT7cvQ4BlfaELgvbO953zpMihYslB0hXkipDR1lIQ
nKYMFsET9z0683Si5kPMcqgTugKMpmbAfF/3fuw2SONcGDvS48Ml06aAx77wManP7GLgrgl2kxmb
7kDfZCCgsXCfPn0/6uNCg6gvYSsDr34dXJWpenDgenZ5xHydgraWGfnBkdsoSJWaw4bFuGyhjrvN
O2hUA1fON1bIKUWFUb2wvpk1DJIQhxgXRHtVbIPJDTaEh6KuNJ3TLDFY0ha/VXdOr7WoLuZJ2hgB
Vzal00uasVlLX937UCwEB71EqVtcnr3b3T+jBkwsxtyB6fpXUmxVaLpxZSRJSyPMwwN8Rmdnd7ov
t3QpgkxuAZCL9LvY6wHDtYonnXGCN2TtNk6ZLTLWuRHacMAgn4nXFFQb1njZiXI+xOtLqTierQuI
5n9tmG7ph/u9qAwFZE9je0vE26D+Mh5/sws+aK/W6b5G+olFZBkDumusDKjLd5bMs1GhE+TumaxS
4wUoYWlJ4NlERQbi1Py0jw7NPk1Owd/Hy/zEFCigS03VOhCxlfQjtwQe0rKu2BT+hiMcx27C2dL8
w5x2FGeFfLNk2dY90uRzCDVzGEGu0mQ/01csn83/PVuqIlGnpo2RlHtRibDbiDBHF8F6Dykg1gp+
4N6ZXOGjDYXRdPBKCOm77/zSf83MyogFoS104SOI16aviRM53SaobQAP/mF4LYeHT0vigp6PzLvb
Q9gbjLGcIDE8JsZds1oJIdyzAsh3H3eXVF+CSEMfCQfR5r8SoGdWF9MNkYZEBlBC8PBVHqA3TVsE
432x3w0szB7wJ1ChPtAb48z6W/kcqXV/Pa90F3fHThiFUAqNGWcjolRiL5z2L66QT1lb1pTRXoRc
+4Ez0FetlxVCFJ7qBhPp+aOEtT8mMju2YXZMSBJYMAC+rJabLnsp5Ig0c13a8u7a38dgkA1x7quV
L8cSn0NoX1ZKdOtAKF1UnQG/NLgmrcigr/Ut0d3ius3LfzRFiklk+eWRaQtzWxgBrAkt6rhOX+PY
6hB2Z4oM5jM81hVivL3N3i7Xc5jfqeKfqWfg8FvHlFO7+FyWDxf9vU+rAIyArghvVNjwBQomQTdu
Xy8kzNiN7t5CCo+r3Lcyp1kkSMFDhADeQmRwUNV/wIriGFO+XjObuLTOci2dEoy3nHP8SbNgXl0q
QnhKsV/9mAXEMp+UIWKCAYW1MjePsXYTGXe0icSq7yJI7l26S0fJicDTxEvakAjvZ0xXvVXE15H1
wuJM3u8HqRBqmmVB69bMIlZV4CF+xKJ/ZZNeosoPzisser/3KAEFMbteBW0iVD8fcSRjQVXG8JpV
0/diuMyUFqXbsNA+W34aRLkpG/lLpxoUJkrlMSvb2o4BT0ph9WcL8nxXfvtK7W0vV+a1WUTXSQcF
cea2qXgm9spxSbKsq1bXRuAd6ksNuLdeq3SiFcgQT5+xlsLh+2/uNmtOoE21LTPdBJqSoeNUlDjY
dcQX8hM+QTDeWvBJuQIXuCYQMw4GIMBNw8Mr+JKihefyte7uJl1F/xB5t6n5vxOn7zLnDosUdy7B
S/eYG8Jeb1hARsfakk3S/aaR97EaJIQcSG0JJJEvCL5VaT3GXCscm+9MgLortblzZzUre9xJ6syi
sCiUbdEm23jF0gn1tDDedOcui4o81nQEWAjaRNnhZ+lYziq+ppzpSFMSQjHGAE5d33oL05rPq9XR
4sQRGgBHBVu9I6sb3uzWk2P0GKE32AewE2wL0TFW9WyesnpBT78bapr9gjnSujqY0yG6mgQCWY+M
duFzUdLEMuJAui6g8P4CDT6ZAF0DJIReaWDZZS6QF+1uvLklyWR8VD8LHDIrZbYo1HZrxnr5MHKB
r4J9uS1N0wQMtnTDvg3x71tu62vobciUrVTj60OQ7clF1g4yOuWQiLJffa5AudA7RtierJAVM8Bi
7Y6NvoH30weK0IMrkIvwsNlt/p17JcBmBJBOaubS2xP17q8spfHOzqnBjD+xP4L+dO6lAbqDG85i
oimD7xO8Rqib3pwxmO5AT5whlhLVfIN999EduhxYaMOMMgnvGJyNRgGNejAA7WDbu7MrU+k7a/68
nuIuHbWlm2I+WN8j2659dPwAh5kD3c+0+Ezj/e/bKXMSD+vbk2balAoSeVHqemXfQOtCCetJDltn
tJ3vO9jVRcUe5BC9XxiOp4SBmXJ984PYZt8nUROH0uOhaGkF9quWKJO2VzDfyeQqm0fmOjS8MJIX
xH297svG/JMmpJPrIy5XbJTZjWrdwKxB2s7oyrYQuOjFD1gvsaLoZwwVe510B/iDQnU+yw5GDpLQ
eb8b+QSI/1vsyJ3j0N01PtAKjhZ4Yl2UFqufgfDMFQUxZI8VXsFoopiZwFFrvggPNcBJtGYdXPW/
gXD27tofb7DgzHPTa2ztObar23MUX44cQowG3DjrRuOnfq+IweeHHN0oSACcdTtQLg/mraSIh+zO
D8husd0ZjGiBIL51I/lfvTkJw1zq9fwCpD6pcO4TFeGVyq/T0071/lvGTa1zm2+Dly8F78uJav+t
lwLSorUXUHM/ON1W8Khwj6WBxsONqL3Wj/j9HginpSz3KnDRwk2UA58xDHqdexhBBsclcOItIHpx
V8dDH6kw02q4qek4DlqMMTNeZ5jcR1zt0i2aC1oY7g72Cl3m10vIJgNSPsM4vahCx3KYFAhrkY6+
CKcmuO5u9iireRKC/xHQKC4tGG4kNoGqsWbtTvuC8fCvQYsnVKgot9UpQh/Eqzo1ck2gub5rEoXk
3HScYYETypK1Cs3JHC3hrsg7rhDjuTz9kT0OrYBuFMFW8Pr+C90QoGKQJb6ip53mIs6EvEzZ5N2R
60AVlrVyN7KFn665Wnptgjnkh7mR0uNfenEjgvskd+QW2FqcJzXbmA/syMy3NNGXnmG1YTby59LW
RtsptjFrRRcO8CHX1uWpPFvyaFGlhT1M9oKVNvewRWeiCHELv6EzSOLRYgJCeJh3XqaPTv4CRI6O
eVikmczTpHRnkcd8li0xFBvcUV15zt+iZc2IyJye3V1+citwN9OFe/km7XjVe7p0gttau6mDRnkk
B0V/XKNpoBIoncDeG1BJfOCFzux8BI4SgQnsxudIVFVLqtF2s3z07PKBQZCbqMoLbfASGxVi83J6
Jijritq/sJjsGZs79vA5lZohfNlWaPL1AxfjBsR9fuWQjFaZqT8FveTM2GkdR1VIcl710+DvRktY
onnmZ5KxCGN2SioUXIePxPZRRTHs/Vo5LRMxjOSrrYjRuNsN38rtYI5NRE+Hxc1ASfyrkFu90XnP
hN86YU0OZNkcJBrueJLvVROfp6TYVya9zHpVPZL8Wvf8Wz3MUXfHjsGoNnWdDvO6SWf32pJTqJCJ
pQdhdm6XEN819q/mnI5EUEVwPjbUm0lSuBQcFY8KjdJRRaGDufXcGUcwhS5YUpzeKh/Lw3nlBePD
yj5LBchbtP41YU/n30Y8PBpp1pYMukKF01f+dOq4heuIFSAjZn4ObbqX+P4NJ6foSnSC4ZmqEs5Q
y2YNqrZRB5CjwrNN1qnE/ZTLysnL2oLcPO+p+SYvHxRtaVnzyoTnorePl94vRmNC9WeokFAexxU3
0OSpYRHIOD0EQFYYEb6RCA+LKXMW/qwnVfNW+Jgt00FQlx5PLyAJCoUumjfL1L+1OUa4aXQhLFJP
lyZiMZ8nwDmWNSawHxejDZh3PWgOUEogFjedBshdv9/bd4Ys81e8PCbuukFxJYtAx3dx6+8V8YFq
D29LuB6dOuDRQ+Z6sRYNbsQ/p8CHtG7CDYRqXz9pr5X/Rr8Du6e35RshXKlDBkAKmgha+KlcFuZL
c5QVq2yTDUss5IJireVddDbjA4EKk1y17+A2ltPq8zq64t/YGpHbUlFpaIfX2b1jFdDKZAZh+twA
+E3ID/i9ng2wj0gfOPOBn3Y+P/DcLKqYTx8dRpe/lprnx7fa+Fa5uLYrg2AgMYDV7PNT5Y+SptOI
nZ67jVgAwhZ725fFCdaka4HH+69Qcm6sWbh3Rk5E7U08syXUb00ON0u9qHlDalRwYo9FVbMUH01O
KP+7dlIgbYmf5SH2Z7VI3KEUlgEpzXzxfqtdyyajjdDpM6i428afqIoSGRqKMeyWdJ3+dpbqRedN
SNELGk+xbpnOxvNKi7SUZmG+1jUv3L6Pvnse2wdwXfdd7bfDs/VIL+waLr5Yo85ZC+PCTj942d2J
XEoqcNhFOJs1URM02biSz7MSoCkKmfRG9rvzix2+2/FwxtMvTyvTFz+Q73a9Rja6KxjPS+LE0egq
8FiDOj6hq4bEuKOhYxJglWsnIgmE/gx+m88nG0lMIAm3mAKal0SLLNK7DfFCBAYwdN14pC0VeezV
y5cUj/wQuwDzQ2hW6zyvZhnoL1DwPcSYJkih8XetR5291G8+Uyd4nkwYHUlRyzL4Bx0ib+XLLssc
OcQ2G2yi3/mXkgTBrdqBGmtB6wH1KDWQimJvWVzessd7eYfgOPXpNWKBA55BBnScLbd4ShO5fHe+
U2WcPkxjw8cFDDz4PZVQl7e5qOp/o8hJ8VyPz1mBsYf8k77nYETIBPGcG2RrRycRXyDPAh1PMGQS
VuxivjKduSvTY0uT3cgVhTxdiSFJk5m6cdHxOG7I76th+ByWpoo9+2KxUvIC39vPmj2W9FAMwVHY
NQAY0eQVJnzpBjv9LGYdqtYJv6uWAzx99yvlz7ohSaeVHoDodOj7du5Bu6dp+syZs802UNH194Yg
bF5SYUB2aGLws2nWK5387lAnOkQmlxZ1C+8i7tdmuDFGcHa2tHcFQBzSZIfcwqgle2t2SsmMtn7P
M7a2kCe8D12NS8V9zO/wQVMD+atmQ3Hw5y/c/25hMP5GhbH42c6nSKRyiSpgWd7eL91dyKycHlJh
pfsFYfsexl1/8etkWTkRiFoLD5MoP0lbwOJyvyT//1Al/YAQmMQaoUaXwu9wlscWXoPXKKrlKRWy
aSrIkBe9FVvvN5MYyApbKcUMQcA7fDDtSsn5KxoOtsdYwSoa/nKgxWsjvDthY9+GE0hmjO0CBAzH
dVqXvjMkChF2ZHi49FdiPkh/IIsfANAW6rbEQI6Gues3iiJGdFAmSH5aJCm1SGzz8PiRltd9hPcC
LZFiofzKCYu4hVZfIf1m/ws85k9L0iIXhXi0rqvMO3eZ3PXhOxzmlHdactiO9GXYlEX7Sd8UjQok
wCxKUHh/hXCFAtZJDPTK1UqFrK6X7+uccqSWtIPJWIhFNpjmuGCdKjNhufs/mFzi38RNCvoCCGEV
aDiTfEYX1Aj6cRridZY3pLM7/0VLYcvsSY/rYOilZx+XCb1jsrIWC1VawXFnm3MyK7lxpO/2iXTL
LJXEjKGIAUV+UXE0lUcq7sWazpB0TXYzJPaYWhi4pief4JnyLl/k6aTlXqKo2U87A7ZunyqWwTJe
je2Y5m3VZHYM7RxzGZuUJPi6PTxg/j4uubkgCWakSrwVOShgzIr1xQ5ujnbMsFhhdaYl34ZE3UJT
CqKgbfzhNuG+quhwdmUph6n9DOL8NJkd4XIJtqYGVkTa5sw8SwoSggjeXX4d29zHsyVjlMhHUM6C
TiM6ccacnOYANbfqSdua7i4VoKHNiiL5AvMLlI2MIYfyfBNHKBZWqlrmp/TgHBq7vOrI79CcK99J
o9OoU0ZmwtMf6WkJLTwsRaQyR2iuW2GD9wj+TrdnktK4GynY7ZHK1TNPVkfSomD38BLbljgdvOoj
LTwMZ+pnj9wT9xMMs27XSb+9Yny8qY8vgvYmCzKjjMTRkmrnA/XJgNqoYkHnTUh9+kPocROszeX2
6ZTGEH7Qgec9CShtg+fgeKGHKTu/eVE+bePCz3YSiRD3vGaOhS1YDN7/Ty19v9LBlL08N9WqhfGH
3LVAkRd4nu3vClk4oyVPNceYvGFSYosw/a7w5fPqB+DVLjpmuQcCVtKmPVyFupICXgdZz794Ify4
iK0zl5ydmCcjZSQoyJ6U9KuRSm9/9h3p5UbB10eI/oL5jaQlXd/ZidWWkbgdtV0Na90SK++osqZy
2Ne9qnk9nZkRXuXWoaawNYhEJhBFCP2MGh4Fq/F7d5PPprMZfDhDKPfAyNeYanqYMnQZDb3mpauY
MWsKKKRhOvymwXHYeKeB6j0MexS7loleyKNdyhQr3kq1DE0Y5BHOdbq4EO314OfA4vNB796q//cY
KF+7TyyGm5E4LXq15RwhxP9xS6NisUVvV5J8vMd+20w2ospESkEnCyig7REY+6HJSENHV+67d383
hyvjOg7P2YaEKsOTDH9FGIDD+VZLjkPyUHA6+U9GV4JceeJREUYZDqpBNhit8bSiwcpHVlfNh5SH
ZvwuP/PsIsv+oMR5cbYFvNNFtsPdH/CZhBVZ2H9JDu3AF7PcqqoLv080uKIbHOyq4gcGTI5HThgx
OukyqJw02Fcoa+vQAgDODw20i2QkiNbZRNzzWt1FXF8Z9ieQ1DyQJrtyU3jMFpRCgkgX/l7qxCjR
BMpd1Eyu4fCOBUA1nt8Pdck2DEKR63Q6CUxa/h6REPucyBU+WYQhOLgtCiHNqsrmBdFI/epANH59
x5CSRxrmj39s8vY/UizGgPdlRt3YV1lOx+sbVy7EZQZKncQXkahHNbkEl5qpcfvZHZNqIrIK4SaF
Gwadbu0jy5OL1iTsLb+5mPAC9/rQey8XaY8kvjV5OWSU8rxzbfEB54G9mwGNLGioYRxyLlqdBbU+
usNxms21acw3UwYhEZulqdvBmNsWwsIaHqJyWBGKXT1MKUg5C9f80rNF+8sXSgqRyODtNFQ73jAy
dRDSj+BH3cJrMG9MIZrsKpbL1Nmeoue4DUuRggdV2f61XGHNMtq4WESOVv9my7X3fhKO9nVm3p3K
12Y18Mu652cVLbVffJoNPoVjN7mHX+KhK8TfidkjKetHKnyHg1hbLK57p46a0y3bCp6yq/YhVzT7
BWAp2DEX1cQCiSI3OOLH0BhNJw4m6gP1Rv2/hRnXI4ps+82QzZwBT8WbN8OS1vL9i/HcglyJy/wJ
+/oFy1uN6IVjT1zblETALmzLtKnrKGq9Gt+Z3WAWP/eNIbSvId2sKG49dHEnlEJ/1dn6GTRkbk8i
95e0QW+n+1cM6G/qeSrJNHp9DVo9GRuB2SQP75OyKB0uUA1/CCMqaL0XxoSOusn8BQpGW80HBWSd
z00zK+KpnJEtQHtleFa3RYZYCZ5cSpi7TccL3Z4mzCaqrUHS32lPeVTL6jgNGvdx1ooOsWqgA7NP
p5n3ntkLjSxG6W+dWk+4pzKjcObDAOjas++0KL92b54fHQ/BzWD1Qe4CANNsCXrMGt0wqwJdaeWm
s2K3WBd5CSbumsZ2C9fmV6g++gvT6YElfgci3CFFZ1MWd/RQtK45xOtfEmowEJ2mbQlcXa4W7ZTg
83tFTuyEw0xCarjaf/sNjRYBdPRntk183e6mP4R7k5ODR3BLfE6g3wBFivIxYeSxEL0AxrQIzfhD
n7Sx+f4JVXWMTQ1+rzMoTfsneYf+x8zXGNeDB16QfITcpUi8ew4uO4NnoyqqRWkq4iQ7PbiK5j+K
xDWUYnlZiRly+z7d5Lg7486McYkfaQazfwktLqJva3WRWLcocM10tVFNn3HjmAkGhbz9i2uTCQ6L
qbvDj9LEJnOVOMfBY3wTGSecLPNDejoLg5WATJFbsnDIcKV9O9XMa+N7MOkX6CQ0TF20E74ryouB
3+MOQK8k8x2zkSt0fhJgEfd0v5aBO4pk18UsCke3C9s0vKFU/SZLG3tUgCrdsbxP2xPDlVLUamTi
9WhvgxyhtSGog9tYNNvx3aRhE26tWoiXMQLrLEXqG9kJQFLhCqjhllu6Wh3wkLLxPTsmWdqMJZaT
KRelB779G2s9tmCPfOfrygDH1Ths5/D81M2yedlCa8g5NDJNE1+VT8L3USH+Pe2Fh8FV7ixN3/5H
mYUQEj+BMyZ5n+49c46rqtvr04nTFs3xTXxSuup1+fKikozSJTxzrQBE0G3rlKHyRIoVY0vCe81u
z+ebyH01ramJr2ClXbb2mCws5XK4BfffxvGSIMUA2OCMx/c5Da/cILgtlsyjjJh75+PHx+68Yhg6
h1tecUmq84Mfp0gnxBXHr18ZFgdrAeFl6Yf80EusUej7i71fee2YJToUtJg94y67bgYRFTmeCKKN
a8PcENup+vw/JlLBHHsP7w0V/LCU0l+yUDOm0KF2JmXUDFIYERdQNqxp9CH86fyimbMtT6a0ycCy
LC9WbEcUVaKT7NcfGYsd7hc+vosGXc5Qa+PUXhb0q08JGc3FyYf4PDcVzLAS8f/C9Zb15p1qt5kx
ri9CX1qzoo5+W6Z1r7mdgdZOvGEI5T1brw53X324VSmkD158R4EuWozGzNZOFMlpK8EtcIMqm8sI
2yWaFaJAOswzmP4wN42/0ATlVZhdYtAG02SAwB46OkU/cKmJzq3FH6jOUg0QjqAKsEa3awv6LbMG
tUy5CSDCbcWUdTzTUuDzCjsWbLXkj7EB4krK9Pac1DRx0EXH1SFYAIKmu/j18FgIqu7/OujcQ/oO
h/JFtP5qs5kc8dQlszfzioaJsbz75TRwXLc5n5Ruy3WNxlrmFaPCzzkNNYwC24e1Qu30Z19FHahT
+EfRYRebwplUl8NjdfBBgdJymLalh3HuzxXNCxfrhXoJ4jXVx/lH5BAnM2F1hTAE+NKupWDKDEBs
VHqkT4qoKiivyJlsBP/XTFS+woKPSUjAo/0Gaozyt1CtOSt5hybj+XKvhuQxXck2Ky15Tku9zHJf
UPPtl9DTlSsGUegUvH6P/pkFaA+dBKXNor0p03BcVskNKm1zQafMbCM8X9vqzeGm06Y2UmGGUYp0
lcmvNqx0W/FHPlCb961TjZJXlNSMuII+lvCmYBSZnd7JuMghA4wefqC+oQP3DxBfn1w7X64mfcuT
JWaip1/MydZk1SpH6WnqtFFUJjUDMtySvtPonbreco0ddAM9hnZuOFYsolRYcYDdPxPomGQOo3x0
DmYS1b6qM357XfOv21MNnPWVV68qEixRekGv4pjLFEfKCU/xBKKMicn01RTQ0Osjm05bA6SGTxVw
+qExRyTRRX0s3bv+Fyo51ZSzWiVQQOx4HIKsjTIkNL4PRwcLnrN2qtZeouB/2LMo+D43FTBFiG2O
2ew/y9SFp5l7cATrZHUvu+EDHz+rYIQqawNBLQerBlsFrxn3clZkkyThfFUDR8N6AXSV1jbsmITJ
0AJrUf4xGS7lrYx5EUmKDTDDLmXcA6dz1fs7dF4HFuKeGwaeopJj5cqIxJUGdapaIZI1dcJfd12s
rQNPB1rrZFkPSamIn5PLvp3EbupWI0k7SFIYeGYm5Os5vaKWAJEoVDENSEb+RRGSM37gENqsUgiE
bOdNCrY0Zywy+ixx5PaMC65lf3rwADA+dX8plf9o1077lvyOgDhFxosFpNVDV8h6rbrb7FL/gmf9
5TH3xPup9boHxldeowy0xNDC43c+CvBr1G5cy7+U/rPlQcZXyoe7rf0sd5e3Fl+MahsQnl22Cmnb
ACciiPEbl/KtOU/+yo3je/1Oo0ZaOeMyRUIS1jAlPgaFiBkNtM+tU/ZTDe2SKzWmgtXPyOS7Pmxc
TlgXKSw/HZZ+30lfTDpVgPCYZpn2zEaBbZIvvL2Qdg5EWz9GPcfBD/OKB3uGYBdNuFR5I3YDxsZE
+Xj9uN12EpTIgzvHK0hH7FTHrgiBhr2vQ/NihqY8CwLlp5eUoqKvkdzPNlv/uVEqmozyFThKAORn
haiydRcFS+RUYBW2mOcqUWlttu1VG4t1Y9x4zQDE+gp5JAz4o/AXQ/D38Sb6WrvHBP1SA6D1S8pY
BvSQJF0NM08R9hSZqEMLjLAc3J6CsV+r/GLaMZfL87i7EPsl0CDmpNlt+hLojNZEJDU3A6rxeTcv
7pTkC6pTqduBMlTl2eZO8gAg8PQA95XNEXcJc+XLlvpDEY0MD+pQ9EkpPJzvoO+QgpH+KwzjLN0J
+ZI81ZLsXtHYnk7P9CauzH3k1HU9aATSrwzIiGB8rw7KsYZlRzYC2/VGDjdSw25XFTOUu48uutxu
BbyANKEf3xtkdWYiyV1JzTNMA7Zo7zcSdAVtk4BgeroueduM5UPk4VHaKn6i5P42aC8ISXQU0lDp
whe14htSBq6r28TNPgzhkSbZluylxiyZJXaRHPxddvt5mRZzqE9pIqGkyFn9T8DCc+WD271E0u7D
RSeUkSbcjKYyknXJ9XeHu2iVkDKj7/71KRBwV/CD57dEQRDrVMuheBmTih4EcSDIbbzR0E2s5lCF
BGvYqDBAxJYjVbyrbZKFKXNKlTyFAKPGEF32+m96ospSpbALF9JtQmTcUO62oBMi+PaY2wjMlm2R
lTocRwTvR4T+Y+B0Yzh2z383QHctjj/DUTPPxEoPBO6uKmKQdYoBeT3lc1weoZYFps/YWPoSYOQA
LDem6b5iIf+v3C3HD3XK7l//KZnCGHJGHdo22koFjD11NjrPFnIlLbFDZDrA3lJ45VCspNzuu39i
TagD/btKldahgqs7W4UF/jAJZY5S7xmjQW7lIFP2RakvTmXE5opOAE3UzO5cgFeSAM3+xGx6vnU6
f3sQ+iHCbl8ZWWMkjYipuR4qRAS9QrK85OKDxDXm8Ykx44VQKnDN5Aw5abu+ZJ3HRcpLsZ/S5tKs
bF9ss3H8ZzYxUW6Xo0x1rs31Q41S/93Wn2ax6R9HMZgvmoVhqVERAOYQCdLZr+0M+rzhjEtrCkuy
GDryHOe+sajNh81b5aThSCV1vC/97IWLgEUAmi2vJvlLibnAt4ai/0Rujh0hH4UoR5VBPUXhPKSd
6HNeTqgP9zRu6VCsyScsC/pcOa1/aq+i01buxSEMyK6SZfOyI7VcJHLfhgqjrMIml5WQ9brGFeoP
DKi3rmgWb1u3RjhYqujWCgiPDUgzDqaty53mDzeD40Kjk45FPXsnX4na2rKjKvIgcyk/wMQoUIjl
+m012FBgv1Q25gFwzNW2uuVR2ugN98IYvPIMax5gSy74yqwnE2AjvM0FO2ibSG3/nfFVOaV+8MPs
54v2dymXf3QhLs/NGGPUuhxz7uilIXD2/oSgspBr6ZD6p+wu+2qk1qW0/u+ZHVMdIuf1/mgy5or5
D+//aAFd+R7ySEydexxmprMoYxcOxMTL37x/m30IpjQFTbuCIYqze7PA9Z1pNcm+mekAB3tV8Txu
Dm9L9Su3zqAZF7JhXx73FRPAM29yX/KdqiUAHZmAGvpVsKKXI5pQL5wupL+KahSMofZ1U3lnl7mV
szhys5FQk9a4npf8FKlPPLql3Ib4bX6aR5ILcW+ZWnImSx8KZKfyFm/j3Xax9sLRAF5kMKwUSWhR
xm6QRFkNwVZCIPx9mKJajdhHQeM0KpMQB5xMJCGLKBiWswbrBm0wxQoXfHTKqEVDR1ApaLjYmkMd
sgfhZLs2aSgMvbs+Ij5doQTElDbNGofjFy0928lxFrDX4EPADsH9yx8befIu3Ac98xCFkHYb7682
O8FyJFqcKeSBBQZEjqltwb0hZ5teQJK5FlA1krEzcMvZKcnFKdYyKnQPb9XIl/DfAabY8s429HvS
K8+tZaKAx+VS5RRUzuUY5THKFVD5AyxVxYtSKGyRKMN2yb87JoWeyT9xNGIRpyIL10LcJUFYwLqS
750Bz/uhyFgFVniHIz0odGJPMYtE8vZ/8LvE2DqkSSdFyuQxUM4LTa3qpXqqTDSqXT5QVZWx41l/
anJojsDTIVOnuiAp1wI/qXvhmoPciifaH6LtxPzgjBgxvciKFArdZ1BeouNbCqMuauTNXkGkkbgf
eq6opAMQvO/jXwIPgw6wtoI4XKq+AnlGYiy7N2GxouJk3Ev0PfJ51Ike5jaCmd3mPAn6hzSME7Fv
Ne4/WN8icXrH69iQcKZVTvUpwgjT4MlSHt9MzlM3K8fPpNn51lKr75Csy/HYepJzZtDWuDlviGT6
IMqqqeBe8KsLczaBNYYQewoZb4QCgeTGeVjAqX+iRKR/Ti/clLddZHgjnpz7wtCAIHinPYMNpwPM
GXcMeaAOkZmQcbcr6xVgqll/jXMqZ1LJWGGLWDMpoqqjHrOOb/fTopG23KZEru1OhQiOLbkmvJwz
rsyOC9GaRjnlg4gE/Vg3+KN8lN19gmjAqN1I+D1sBlwAXfb2yHkDo+uBRFx33rBmOfE2PyYdUPDR
06Ul9wob9ag8vrZekIta3TahE5sMUugvf6Viy+A+MEw8A439Tb/rNECvW7Z4cWAO65qiCFurngSw
fKpsU183skSgfDlnJapU/5Oz00fjJ+Y4HkD3J27YRacgm1BYfPBEa0mIifKtn8nYIUDXt6WM4CDI
Ec8J+UqUhIPjp42IO9qtaFPLubCY+lyDVOcBiViVYqU2lbTgmo+E6no8ouPVIch8s2ZevG3BYLvX
3Vk6vPO3BZNZcTPp8DyXsc8eXrbpk/vBOv5u+RCZfw83lS/SkT7O4Zpr5KdAW1JFOjNxuhfEHXfU
M2mC/OnJnoP8sXSJ/bgrqj21T0HfjijRzwML0klN/rt+7XZkkkm2gZsQTPYkDT57NsqPKp8e+th8
VYQhlKpzZbVS7CzWvrINC8hUSSpBAYKiglDhmvfouTsS8NZhpsj4mLD0LSrXMEZ0W0rFN9zL1RUH
kfv6XKxuxFYdIUasGkR/gPOTId4QHUW37S5w2mMiVQRyLeQvdCpIxpP3//YSy1AWg0M9LoqQAXX7
zMzjgfd0tZHqTH6NgnNEoKjQQ5okoIcjbv12VGRvKZ4M7i913LRrOLFpHcO4Wc0weTp2RHdy4wmG
uBTeRAHF0LjmW9FN48q3R6leJSz400WwzqRm5ALu4+ITjDKIx8hExHnikuWGMxHVSh+eh3vGKcjR
ulKBerGrxmHitbh6mbhSkwDT1SHJcZ5lW8wl2sRzS32HKNudYhOxsQOs9rZLXh/znBd1EVyrc+b+
Wse08biusDmv0+2pcHbOibYLMHsXUkWUt/m5V5CeDEu8MYHZAyv+PY9NwljCFgtAsZa37v66ljUx
6GjlS6/hd/r2IX6NIQE5LiWOJB+RVVpsyAOC5nJU2bGUabda8yPhKCVlVKrneLbQMJNdoj+rKvjs
MIjT0X84DUQ8hntiSHI9Wc5xEXMA8wiZvfmMxTxCFt0m3A/G3HyEzQlkroP5+MbZd2KXCXdNJFKE
jiR+H6woIgzhuyQpqWksH23kiUPPWxem3SiunHD+or9LpwXQ6weNxMheeUMYDflSqsruBKnNa0tH
tg9d+y1zM+nFQGYE3rA8mpTpoLd1QgaWeFNXI4LITsmUC1SdaD/IG0hjyRm9Svbk/tWnU7TnzgmT
Prd56B8T4VXJSlPvIbDoJ4HR9WS/dO7+X8NcBZlKY8PBKCz0V+AMAHavLxvRe2Dapnx0VuAeNmyn
ryzQTIMNTx+PfWhl7nK8HdY+Th3X31EsK5FWEhNxDcvJp0fiN31IMIQtCCD2o+bxo5rn+eXLOiRt
0p3VgfFG2/Lm/poalK6arOl5g10Y8M6Njae1BE8IM/yYnNPt4rSWH0gr0t16aKV73uBnvkA6uVn6
gEcj7mtu12kOeRAhPSAhMj+vbHgBFNM+v0Vs08QtOCH31zDwJa0hPfZeOmKG3dTC1d+Oy/JCH/M7
kpGrIwSZjcn8UL8K3xbwdL4M2aHqUZKiO1kCXGyFFrN1j9yB+/5Z6Y19PpF6J0oqeduMpuXriug1
DQn1iyQ++SF22vI7y90esC0j3c0bDVRLT1Y7uJaQYgHeDqd7WYzlUf7HbjRRU3WTlyHYBN97iM3O
/5qSKk9icX8IlPOzq+s33SN155ZI+JBp27EHRpOG/Pi+M5PBpKKc/6ukpEGWj77Cl/0ir0RNoFm5
MVeLGVpplALlwiXQvZKKdmlM/iY/UvUVXvg4E0/wpMyDX7Yzoy4M7RTYWkTPTkrUDFWEyGVQ6k3O
7u1kqHZxRc87JeaSxUiwHGCBnro/MF7v5xw18Svpyd5RtnkC52PRO3vI9Ex+j6mKslNBDuLx8n9J
/6xSAcSrUvW/gdWs+MoU6oSn1gsIgWW4/ZTpBaZYCioUgAdAUWxgvRwF4AfooYFSmWNZl6AsiEpt
kkG4E0ndQ+Dk9CycO0QIb0JIbQ7emQPBgVj6CEEbrDjrf6+n4dmZmTvFLu1iFmIgUVTACymoxSbA
vjit/bfgbdUEdKWnXwGtf5htcuINuSSiQR7lwrNC6yR8IvPbcdwKSqySeuFZj295OxVZJGwyjiJs
C9VTsDNMIcKo7qNmpq4ft3s1P34k8YOvthpnts5VI8pbwcwTNo9kDGG1TQvKWQ34oPV/nZa40s6g
oGpQtDm8w7tcIjqeOTw88LPvnHg1Y7nOMiWQPPTK9oRvPMCPsH9msl4Rn3lk042vr08neQjt6tsY
mLXolHY3r9wjUVB/wqhXWPHqcX1+FmR99OCoZWJ+Ywvh3B4i8YfFNkKaT3ebWKWC/fyNZhVzeYEy
RL+K5mT6AygBD7a5ecxbB5c1LxM48ozhLfTIwweLqJDSMn7mzWSKNAl2DqjRR87T93DiJkxhQrhG
C0nI3xPdWAuKkXqSI+IV4y+F+u2WO2JdnaBAkkTRZERos3WKxFrZXsSl2TwjFJz9oEmlI+YXbsWV
3ieqGH/P+0j6UrdSaKMZb8iJFXxAi+X8AQtMdhzQGXHRV7XFp3dO39IlSYsCAi2erjzBKIwbkHBy
bhbXD2e3MJkuCZjIhHuM6SehQbPQuuFOoL5gYaEg1MkLwo8YJ5Rv1uWbGEuFutfhCURtG9nsn2AI
cpDg9swF00vxHdL6iP3Iv9UN50qqv8F0768i6X9wfVqqYUDz73ShQFASfJAxi0K1K3Op7lf2wun1
e5c6CLfpyMPt9A7sG+kiRHVpEc+/IoQc/UyORb5nhOGFg6wHRBRK55gxV1hD1J1XzIPSRLzX9cXu
7H9lOX1c/md1QOUVVLdbLQtI0YnFZHYFPi3Xy78ghCMrplBaAA9WiFQGl5YHsW3LgsVLwxea8vHh
CNcgRsUmFe7k4rHQhQuKdYx8gA0MY7B+DNRu0AjDxjgh4WEYavI9blJpcMSVKfqRKAXfmCU25i9G
RUbQz9R7AcZBwix34Hyi+AYdDgDtsFDE8Gib54279X9PE9lfHcLTkTOb7/RLYL3hH8bREcfKxXIB
KqeEXFganY6WfpkJt+5fns3MU5ox5+wq5dw0Z0WI+rZbt5E7CsGL06/kVTlo7O2F/bHkb2fyXssC
Q9AgPnbcPDAfhQaO+TdivG14tA/E+XG3zQZsQ/41TOTQJvSDo8koLNM+zNQiCmQi4kRF421Mn9Bu
sx66pbIEpPIhTNXF5GUCivJpiXIEl4Bjg+PKaNLqMuTCfr1hEKWOfjgREZDLmfraNl71MRb4jhWf
47oXEgYPQXOEphri/l3n1iG6P/pvNXFjAvXOP7ZK4pt5tQFi29JuCqsDpZnoYF/4wMDzxmo5PeLX
TSZm1dxhU6P4cD6W65O+Xn3DVd7gQjw3rNSBkgC6o+5+2yQBzVQx/lwaxuOdx6NEsKiN/Tq/4WQI
jTAAp44U1NfwocxEL9pyXwqO0DwKUcCMdM8A9YsVQeurORdwLCzKBWiy7iYCGdycwM+aCClJtp8E
bBOXqyQuQkRGCmk0a9RmGoXFbvLZg9Ty7U8a81ier51nPBXctVOON/Uf/r24RtRKv7Ma5LQo+ebY
2q+iHR55esG7IqEYcOrH7aa+0qgoH+fYHOgzr2q2SnAKbdjjv8QI0W7XAK4VJCj2EId79QwvKy1v
1Bnl3/KblJ87n9ximglbCby476Qf/aPxkHc0nIndeVypHb7UTomYm3AvVre/m88c0IRdmp7Vxz8g
yVq614qJOkSb8oz/twFxsCfIV3SxmUA9vWPnq2EA3vCyHFfYaJZGj2kBugvR97JqOubHcQbwnb00
t1M6hz1JUT/UD7XZc8kxiwuLsctY/29G89xxD7EGyhQMK+CELukPxiQHI13WvzCycvP9GDpCrZx9
QIEmBfUEQWmFY+VOg9qIUcBD81tXZt0d9lEq7soBSGmWKs08agINL0WHvfLZi+ngCnSiQvHwk/YW
6HbGvN3qfJ02iF5+bY8rTqzur/lJvnJpGuCNdpueyemPWii7pgo/T8nh/wTHsfv2RqyP89B3FYjh
8JZOzwCLeqKRXZEXfUgEOREH6xOBWGgwA6D0AwIedYMIHRA5+YRzWx7iKmLXCiW4rT5LCds4hQgQ
cwdXB/OyGM+xi5UPmMB8FBBJagUPoTtUom2YCkx5KXjwJ2sE2JMBkCAKuFuJBXOdqdK5ZwZqEWb0
FlT/YfgJfMf1KNCzAxzJvZjyUxLoVBq23WGla+cTzrUIKqU3GosjyDcUaIgc7S4UWpd7kPbeM8pd
jdZxOizwR0QBLG18EI9EVxKbBUcN9YgJI46oOcZt34ini83GDKTcVOnsWvO5q0ufgh9lFb0kDQWK
cph3ukij04rQ7KELnVuFX96uRe8CXkpDkl8Mda1nYd9AmEFiOKrmjqjdwYO7BJUnnBZ1LLcLHjhv
RuKoQSqnQc23qemEr0nLcCDN+KMkqO7wZHEF3hny0lKm0pR+Z263/a4nVxOQYLaLvY7uF6Ue4j58
wh1YYKctSYoFAiqVXqXd/i39arQXG8DXEZr1NZD8Cp1VPCV87w77xjrND/r28H/ofzJLGhkCFFa7
yf6HDbd13oEeDyrQlK37TQ5H0yOKXxNRtvaTG87QdMEdb11HDs3qIzN3wUF8b0nRVaf0n3sdRLtp
Fm3+ipfx3/fpS+sWplxEE6pJAdl1CWIRiwLdMRnX4aoare99fihH5BeRh2ehNp+3lTpOCnDw/JIn
+4nUzGZ5x+mt+We/N3kj1FFFoSBYUX5QpWz1/rPS4OgI8khR8D4X84jz0i61d002DVZOGskct1x5
8SVEhys02Fk/v9zuC0Jgc4Mfl7tDrZNr+Il2lP/c/ePkE00MAMPhsQyhObtUlVwce1s7vH/RniDk
95i4x6FOmQvH2pyB1OzYNTpiewVjOFCwdTBq0HNGuBrTsGtWdCnKub3hqHrcjkcdZIR2FwyT9iWa
QjGK+NQBjZxm9Vrus1ufYknLSWr1sHt2Qe4nHt8mYnzejGp5zOJHxyE8JyJqiY+JEw0QHh87E1cB
z+1VUkTeb1S+kPi7sW1iQP/bPo6ONS5j3TZGYwdCs/0w739C3XT1F89vegP15uEaxbP/nzn1QkXI
0ekNcb+6kC4FlzzjNx9i+UBDK4pcuy8/jfY3jRpxApxhRWWg83XuILI69n5IjEaA4np4T3ANPyM6
o4XYPElvqBw8Wo56Gxa05PyoB6P2otVIvLG1oUMYYsd5buAPCS6dPFwKq2EVYNvNmX7lBcgD++GV
SljBVpe8/L+/owE1qF71Bk5XoF+qH2F/A5KQpwQszkncIF/+XUk+wDuO0blFQcC8KoFMwjGHMb/q
eI519MU1augmi153WExVmtS2ItjZpzPmDXK4I1D9z1fLvL2pis0yzvWbJvR2OrKLtdmMv8cAXsHQ
HlDSB/SFQdHMTKtsiAMBlAzlB4Ks3mosKw4KczWGgsDGFZyp+uMmWHvoF64435UEIS0PaJ2t4Yr5
mBDRdv83LMrBPyiN3Y9Qi+h+l6p9uhn6IFi71k6/A7MMYlplJhU+u3IkDW4EtG5F4pl60z2gOk/n
0QxcKwyvD2VoNWA09ejQrayPBYWsiFxKUgbJe14ixLj6sDcKkPuXjhFUeWPpnCgPJYS94jihaU9p
w7jS0SW56rrFdBsde7RKcAJ8CfA8p3zh8/Jvqe66tneAJSOw9xelF9PLuH/Tqm8oEzpKVqUEoIUs
lRG33cUlzuY3GCSuMyxMniDHGz/PR1++UEsTr1wEI2MI7R6FA2vmLsZV2pjrtknQ2tPrjuhfn1YM
YsVmOYPcG2fO5wa4OH0m1eF0zb2rhGvqMh5tu7dA+4n1/3+72dL5Ws/QfooErpgZmU+nav5ykxhK
a/CoGbDkXn79nLjnTNRG9ctvgL6fvM0StmZnihSbtxI/+Zwq/yVYrswq5NIwXG6T5jkJ+WCW54Gq
f2KzAQhhabpFaiIDrmC1MKnmlThg5ZcsvTCr2t0EqQJtJtWv/2BzjJoOuYdKyqVMEEX4IosXrfOO
7oY2TSauy6RsBTWdyH7a279gok3fYyBDUoQbV/sURsEBzezk9Of4J1HjA7VtfzF9jyIoULKQvat5
rl06fbcZaaHOA4XARcXrCQD7VzXuNiA38OpP/KOLUyUu7x9iuvaxTvD54ih1XijkwGGbbdRVqbrk
3KCuC8A+D0t+C6kMwuIerHtgf+X5kyCmc6ZGzpXKrmXLH7xdz+t0P3/uI4rEHarH+3frJo4KrSCg
aqxhLa5efff7QaaWeWdmRC1LULIeX3X0nSWa1zc13A/8i7P8RMeJ904Aafk3DrIrrFkUP1X/Hkjc
83AnruXaLpmE0nWxmeUNRM2PjudoAh5ezIYq2VRr5tmsagBGPoPkJpoUQOLOefQLbQyW82QZpByz
fHYqrUey37MEzTwDaIxMtSeuBXg/WwC17SIKsDK21LeWa6qiPfWtgxek7LSCHkLC4hLVJfucWJpl
jCIv38CvQ7IGCumIZYk7FApW29e1dtpmeoSDwxAwc/zxyxCdxIr1Cc7Y/yf5/sfSmJVeStWcdjfF
Y5FkH5KOXJbrSwozDqMixFv+GCnkfJnBtcPS5UaepQZXPZJDhBpEb9HusIL2rxrdwjiMiRmbnBtu
/m/qpNxqywOCL+KlMQyJvmw2RGBwyGOJAqvZx9jDpqx5MZkTdzVRSpBUz8er1EWEILCFCKwp1kq+
p58xeJMTP5s59HCK1oCGq8Sw2k9DDxlnI6SlU1eyhwd8fr2EXhST9iIFKZoe4G+z59rdFb+r06BS
yg5OFZGknZKx6X4ZlzCI//z4U8i4PCEjzqugZBX4/nOYRga8XLmdBPsPiq9VCg1PaM9gnQQQwade
9gfGdC7DR+VaWRxnZuc7tIdpKmgX+UC+8Y93CaP1k2uoN46hMzwcWLRbqQ7Rz5GrVTqqtxtYVt8J
Pm7c5TaKHkMNeBrXJ4DpQoFHpkLpiQTesmrt4qrK59BrcZlQ4HdfUReovt5D0sdytlj6P3Fl7fpm
Z3oIWfGPHqYJvDyOf0T5k4gbIFDXZWUKM1TN99WIBEMD7MENSEKbtGGEsbjsMYAuuEJcpL9MFjUY
Ol10sb7iUQDmdq3bF76TxiNGBZjcttYceOAIftGzVbv5AjPlqKsdhoUyVkpcDQvmuzGgb4UnGi0A
f8tVCwyAJpjllHhxbrMlOGM8v+EsDo0YYodL2zbCDo8sVpujnrASSKqT0uOZNH1EgB7CUMCIc4GK
OkOf7qNDcpGJ1SSG76KNRfluUZRaMJs6fm044/ouas93MdLLev1WWR1W4I/ol51sqrx+cOaLqmH/
d3X48plLtZW4XoGe+ecXYnu+BAEselDR6xcsXNKJDkrVVHA3HOBkC4cEfU1F3GzkXLmK6yPUB4qc
V991LAra7X4lF1a/PrfE6ZzL6kdNxxQbpnyNGP1mf5NpJz0xjM/9RjSwdIoZX+wckRymr0fZiUYq
wXnHLC53BdF9U7LB8Eo/MJmgXVm1MIdqZoWcFHQVopUUWJd+9E4Q2Je3zwz0vzPwi9Ve7+zfjYEn
hGuGzdbhpckFuyNB67QL48i+TsrGI+FHT5wJZft1MmV3Ea2l9i0F1mAL6m1Wx2IotuhOOTxGnJCF
zIRKi97Gi9dsmsL3udLqNIBTTjpB3qu6Nw48To2C2RhpYdCgDXj3OoKTHZSgtkpGAcs3uayV/tbQ
7YQDu7LTtQZnmKabOQWvHK1zXa11Pe0jEYnSlpHVApeZ+L8mMkwKS9Hua1lvOYFEFvyLo5ypCo/X
TeI7aRa3edZcV60Z+xqK68tAFlO6D/ZlXfJxN5g5fXCDpMs63SEqnbHi9wlySVMztMLjPp1O86PX
lX7YJSVE6f+VCdf6sHThlQ8Wigd6SgZTU+TeHqa8nGauRjenMU0K5Of2+71c90Y3/+hkOc8vkDko
98GP7Ym5lX3NgoGGH40U23itb/VPo0U/sdh+oyqJwJjeNgCdSTAscySoavnaJupwgNJ41GdmXHVD
tVMm6bX1FR50Mjj6LTedUCyCi1VXQyoRPka8AaOOILNWO0C4ougSqNMSIcnv8VxmuvmjSPjV4APA
haRbpmw303MJWw0exwjTZaYVjxPOyuniKYtUKpcj7+d3/v8/Pu5TSVQ/hLfujU6bKju/dx05vAP1
Q0+UiECdXJxDG+BDudMe+2hjjY/ZmVcU8+yyOOXH2NQpkXCBRiHr15RXhxhfzh0IORIh64m03uoG
esRWuATE1cxvhNdzX2ShFLSCOnF/WOM9lPXSnpnMeX0JByjhNWggbKr75hzaubuA9m0OMrqutxDD
pscfTE/fWY5lkRFcqEhfvYsmhyLbeuw4dA/yghpzQ6OZjmbPmYHpYcRlXyZvMIPya4+ZbHj1VaxB
WmTWMCcHcDWNLbP4ziKSFixfY7bma0y3yyVwaxkEj3YpX6RiOBceTydcAdaxm9jCcetMnqZhPDuS
OCqIkmCmIWymRuPI3+TG3q9fyFukrkmCELor6AqAF9dI3gb/0alOuLFtQz8ESkFNs50TH4D0ddY/
KF1IP0YEthRXY5Jw1zI3MjfvtwQj3FonKHGhTcWDMx6NJdMHS20//KBo88NGHZazEYG3irOb+JPs
CVWPFkzipncoH/SqJnA5JgtMjq5O0RUMiKYB7rxua3YL7bnNK3hssMbgRXgBg5arTpuV9o3AABc3
Du2kZu56cZETZALya5QJ1NGrlIZkdAfRnnWs984VZQzj0Gl3PHOwohb3KKiowoSlZ9SoMLt6IHOe
HXkhBBeAGF0JftLAlI4IvFAe3r2bMJLM70BqRIk3W08X6yWFkTXA4NR+R+ll6yDNq0ZwIfm/94zL
KmvgXX+qITztWf4QyQENffIs4zyGt20NkJvOIStQAfaJ18UjWe/xfgXZwLwwMse72kjtlatGyi0U
WDQD8/+LkG/uVowhUj24D8GQJ9GVP0w2WOJ+FXdp7rgnSizYqWZe6a97YkVjzd7cX3CYrBe2Klh/
i0CdUznUeuHzZpE476baPLTY2rO6wvGxZhyaT9ODrauzGLCMXlnqU1zR68syq/EqkoFSf3Pmcg7E
5zVVwlCoikWEqcoM72jRRukGOBhe8MLzhyHnfhqFIiVFRu5r7oi33u6mhN4LjShaJdSvq+eRTftz
fPwk0LtMO1MZteHfo3l4uBcuPr7OqclHtpB7EfJR4in1brLhyWy0QPYmfdz94ZqVt7SrpKw49tTF
uC/QWg1myduQrklXgQXY0YZ9P0P0stCRGO0OnpgV7KZhDpZyTsM4my+ud899DTMG216ebGN3TILB
UT6QMwtrFNU1zZQk5ofvxIWmjKnNIdq2dTQpDwP7w5DP14pE3sgoZ69JSHY5AJPubUDRk8/qgLLz
/kiITzP6Ln3DVwRv58UThUMkKKO1qnVesZoBRafshYGLqqCOnmi3zrR1srlIIV5InGZdigmlWF7+
tpa6cI5sk8Ytn9N+Baef5srR5NqPtMxc65HS6lAZBQvsJMXZ4HMwIw8L/cTPFToh95e1h/+54hI/
TRtVw/hDV5aRPcRxsM4FhfRdCwPigbjZszKr/g+BhrFr3AOtlweGPPzIlgKI8tiBUCojiruC3bD/
srMGKnszDSggWzdynG4Z/nlL5kpG1y7o7acaVWx5bA/JU5Z3vrLSTAF5w98USDiF7THA7r6M/UfO
03YOX5/d/qkIPf2FnTa1sUh4/2pInSCaJ8Q3Dci32slHjIrremqxGmUOeE+gUr5tDT+tYsJsauoU
4T9ML3rcTUsoLWVEchou1FM9Y9sPCmSZl4OkaGIlaq2gb4t4MNKpvV0yUe1YPeLgT1Hkt0kyl4Hk
dfA/WyOoappRSKb0p0qvwGQF+eVcIDoP2nD7uu/C6eBF/ezp61uGdZt6Omf7GHE/dScGox4/9vNV
VU6659zAUM9p+0n2W7NdYui1KguWKasjMxNJQTMUpZI3uvEtCXLLRh5PbHInHG/0r2l85zgt2oE2
zqJesy/K4IiSdHYpfCVW9AXUeDl9AS/DAdMEB8VasodRFmfp7/SEMciVAAh0WLWfCcWT9LuoqnTK
FjQZ01tdTpqHaThN7kY3R43rXzbv3EaMFjB34cOY9L/nHxHrAIc4j6G8Cb/cbCo9O6kOEOFnPLoT
9KEIEF+mtu7V7evoc8j5NBsQPIPOe87QJD1SgW0IPmgPkTfsQ/Kov1SyDdEDq7rW9gSJbH8ORM2d
1ewsp8dZrOuQKP4lFAw0DRP+xP2vQVxWNhWC9/BeSQ/Rf6UMBvYp+tBSORZQDYZxo0h7R8VtiyOA
s5qkBtqjw8UO1Q1TfD+R8EjafGHZGT5/Uk7HBDlwFp9cRjpom3eadY4P62+W+KrPgF0bT7WfCMoe
jLfY/vl/RmYgoylOajGgPaxW67tprlfDy9skcx3dfH/j33Z9nM9QmnFwSSRH/hrtKPtP0wy5JaA8
FcFTkwhCSVJDDxCDw10Ut9OkTehiFDCi4ZLYO/NXxvOijjEKEF3gGUhK4MqRiHVr+dX20ql/c+tD
mvXosOFJmysKfNK+h+5vMtWRXc1EO5ugM+Iyp9DdQ+6ufmwAqekEpyuZKX8lKp/ZkoS3NiQ7Fa7f
1XGdf9sBKGKfiKlKSQ52VooUyVnGMbn1+oYBzusb2zt3dGO2AIche9Go+dfbz7F3ZyloxLJrhRzM
UGxAQIm4fBSMYJot4A77JDvPQT2QWosnGHw/g0ipjpuGNWU/6vwksnGZnufJOYM1GHBghKUcT8MY
CdPFFOmDiyaPQGGLC63MNHBtGgVtYaaql4x5lztNjXKs4brMoxbfR1xUOqCkw39BSnfCmgSd8o6/
bTcbIite1wpgKGP/rhtsJ5U36YXcvjCDwbYhFaFfG+WKPZNTqBiDYNMbUsTJMvRl1L9i6N1cLSm6
m21sMQajpx2Tp3vCfESDbP0mjMm9FtM4x9ZDxL7Y3VUK96tc18NkEVcdjckHuXE2fkWYxLEgzdtW
YQxk0bFSsoutcV9KTQjiggAQgwcJf6fSs5nb+EchuODVaAcHaRqE5CteF7m8B4OjvxhF3pEdw2My
ODHSTmY6lYEqkZh8MCpVaKoU2B132BjBrSSS5o7kotaxl8qzAIT0Qy4ZyQYdfJK3EnLJOWRtt8yn
LVWukoy54N55zt1gEzPLwwrZKXgpliiXid8II5HhTcInamTCdaWsv9PT7qCQ/jlDbtAPjegOqvaL
Hse6FQ0dwxInYM8G+C3DjWjqH/11E5dwslG7e43/uGlL2BigFDV7hOFVoj7Piihgdhv5iMCPpT45
r7PlvK0rkX8y03OarTGel2oXXNOy+wTt0pIiR3lzqLFMGb4FBgu7jI1eR/fxd1r57vQbtrtlA2hf
P/kleDKCv5yqvLMu/4pAbGTc3DLWvkS5YJiqLmtad39oz7q1myif7+5PdXawQPljF9X6kIYB0uRo
t3h9Fv2CZ/FzW+qWKHfAZpTPceMCqWpEGfg1AwS6GyGSXhAJjwvQEhgj68yCtTBYGyb0z9fW5eiD
UwTv0mAF5+FzJHpJEp3WWQT9LnEXIXv+LA3h91g4EcL/dJs9/5rX/mYv+kiJhmIPgwKG74DD70K7
nx5FtPfqbA8eJ4uYq4ceR2cqfjcjazQUpQgVHLLcT83VUI4unSvTgS9aoElBGeUorFOe3x97wJjY
jC5FlMUmlx3nHz9mKonEIVmxwd5KRv4bGKtcXb0FffIwNg4c+Hu2N01iZRA8vD27Ib1rfGIMamUm
myzafnOWT9IvTNIuVqHxJOPACpTysWnz3bbEiDr9vOU0mCryZCFjo6tyKw61wa63JMjaic9rFjdE
qbZnUwZXT/303mJNwf3HOitX65kxqDkSOs2bTovOIwVw5nLDxtMhfFpsYescj+54rahPTBb6GbBu
rRoTqUjVVQ7SC52up5LT4gjXELZXfsVvrDKkdWYDPidHFRwmcUQZfZFjpOjhRdSmsRmvyHcaTUO2
PKea1HOMnzFQeflfTTXgVnRm8SRuHMl0lA20MHCWD+FT+ILDygN9vKeK/V3pOu8ytAoR+lwPklxF
vFVhFjVSadH99BQK1SLM7rK5ikijl0RE8JlxkA6FSpUGHaH/ZiSR+M8D+tV8h3t0guL5j51Lh459
NriOHOW4iH34NCdFj4AD91zPBywQ8jfQWkA7wbPiCoTG/t6JgY0Vc5wI61qLsBos+84/KxdMQPx8
qI1WcnEZ+2NLwkkJhFYyadNVRPAMNudhhNZfQjmkSCZ450jqW1qLCP4DFVHi1zBalI+Nvdj/DnmQ
nN1PB144rPOScYAWu++Ua6oYipmxh/FoGRaW24Us3LPMbve3LSUz1A7WKMHkVy7LCVfCh7Jq3We9
vOJHIh3fYh0YQ0bet1RGOK6OtiFPMIU3ZjWOSv3jXc/d/SkKo//NpL3doNAA5avOAnzi79SQkG6k
r7f3pbU/tn3SWtma9ZZ5ucEqhhC6X49ZojerBpAW/g0SDJuVqEP88lpkKmNPRYmx0FJWEsd5pe0K
VG8wU98tGbxWHKuV1NPhP29PzzDRp/lIGUYNJld/prTOdGKagtD9RCs5etnYy+NlO3oy2cRn5Mmx
cQVBtrBdPeKGWHAnKrzqmyLsdEdlq86O77Celbfx+9p4iHqzUqC6Ud+NZxaBTeUJgbirDVOOPzFZ
mxzCzuo/KGpJZWM6h6UgGq4rbYVMJckuY2XdTLwRp7OxvpYzu3YTf3yqvC9FJMxbx7UTXenX9J7D
0lfrHRSE8Qe3R9wSSItqdQtFGLwjlQOTOdagxGwLBzN6hSOfD/fxTba1ve6PjLSJBlQ7APMBmxds
1oCu3h9FYvu5IxNbD3dmpn/x7xHtd3FE/CnmKO5FS9KdT9Ynxo2MfbG/Ud2cN8SHBFuFz7LKbOJB
BZR0Ia3uX3zJvA7zRpQsvLhnSOX3Jy6BD4lUnwb1iDnhyDm0IRMQHVFRBgFaxDC0PYKO3O/6okKK
JLzfaP25vBX9+P+KTJq3ibc6suxB4IIJIGI9xVEyZAAuaamSKy5PnINLcz8m9qNyh/3hjEBYZO8P
/7G3b12evv4l+k3Ok1RgfJF3LYQotIYfAd1zmoN7r/NFFmL3e2IYR1PIoEYCBmW9av7IjV2sZ/30
Ns0kQwj+Hr4aj5z/SqrkmHMEFOMiyo+hLBYh4rs/sBoPnb5WqURpXRRc+RmQE3sNuSR1+pWiVg+H
Hf8MUyFcv6wnmFR9hbiV4cjRJwhCrSkEhp4rkKC0JcxOsb+zM4+GAwkZDmFyauau2kTFkdLOgbuN
uK9ALImbuqhPsX2cKwI9oYW8igSPD8nQVO+IARM3GQV+TvVhP8d30+Za++8iJuDaNlOBqDpwNmsm
rQC1pm8wjYPmjFVwB0oYkU5ZRfeHeU5zvIvGAnfGlLDZNYiqpB+McBzOBpj8ymLLYsQZad9jj92Y
hOuyTykA1pDNYrakPRx6CLzXwibBYlkxIliSjr4i4E4VGpIjKO3nLk69T4HDVM1sEHizBra57RT5
oUWfikb8LASBmfzVQBofUyyk6xNf/Y5gOuvU3Ll3QNIX7Xv1Bv9CUdDbHEyO4UlqRlAZBUqPuVHg
9L8uTfJ+LPjTyD/DYKFrRwF3oqASbeZkXM4znxiO3WyPl+AlAPBhKR+oxghz5Pq2ugre85hUS3/R
f7x9kjxqJPYMsx7yQnrdLY25WUalsD8SS6WcGc+FAPvLxjkDrC2VuCXkaWGZ6JzuQFpxPJAnhJrg
f39ThH/1HNpl0qcSQQse4Yz18v6ZrtAvXeF+KxRzyCbFfNIk05rFPXi7cddDcKRF5ls2DdKjpE4U
S1Ktf3LTPvP2D9jAd/C8Z/0ehed8yOXc81j+E6lpKZchN3JqSVQod4aObJ17+Bo5ljOdY2UW6xRC
3ayaxSYm2Saac22Aw8DPqT6wRjeGiTQAjpeGT6OOBKYAwujTww3cDkyYiDv01CU/X9U4wDeEOxQn
dvKA9w6GyH9KtqFR2NQuig+PGYknS41/v1xC+54Zlibe9T5Uwnoay6KGsl2HJMBTe6uexpisbiI2
QdfSvxgfIZwVcj3mhqdu6IgInavX95cUGOsyGHtEVykjOYXka5ZtnYYzo+kB+0EsPwZ6BIuFBeai
FYN6Ik1tuVW8xxLTvh/sxKMdjwqnmHnLaI/S045XD8lWuKC7cTNDSpYpAw5YYpqNT5SVFQyroI1O
U1qswD7PSqRBm0ju2agi5rYLvsY9y1XRhyjhaskCx67aAHrRExSS/q8N+C+qaUXv7WHmRep6o5+r
FdxGOMkbA61lxUjxJMvVrYgJ3dW6JwjCoRxY5MQVru7nh7OmE/NBVtEpsztmbWrkIogSLlarVndg
Szq4VSvXDpd0Dnz6nxYw1OAL4eoPUAU9s5gcDfhcmIeo8t9a2I3CluljL+4tUa93J1edHeazO52z
0M6N8XDS4VBfB2AgOZVMRMES55N/hwZHugS9+nlPMmhiRc5Nwcpf03EZSNJKzl9fUf6Z1LM6ubbC
wax4QetcSx3ZWVdxX+Ofnna3dMEycopL27TW3k1BJOdjv1a70E+pr5GmVwGj0rjQgdqMaBgZDz24
q0hLldlkS+enB4pIxZDDLwi6yl41cuzr/br15Lix8wRsq9l9RWyxCiBFxcKYDh8ChB/1X9XKaI7h
kPM9ZsdnUE/6mn9zhM29xuZtphy0iGMiZUcIPn3laP4qabxmSTwfEnwhsrPIbtbQ5rw6TuAqUcEd
kxkZ61DiHGnLYsOqzrEWvNYxCVB7BvjMXx5nYUnJCXBR4HVmQF2ImHo1TpGuOscNy00w1ABqdGJu
05EBqXvq5UYPaQw/J5Gpmjjft1c0qw1V9Vgi1yTQQK83Pw0kC0VcMi0wxxjQExM3K37Celon8czY
hyK0upFnr/7BSoSbhw6uXHpgMU9Jc2Vfb+sxoroQVdNL5cLuNANk/Pf45Q/rIQwPQ4tfor7oeOti
lG4Tci2jF7BV35/RR/UxTZv7P7PJUpJ2GBc1di9Z+pK/++JQuFk/2SjybttmWM8hzt0ooYw4Y5Gb
BpHSPnz0ZJeoJHvW9fsFaVAFn6CnXiDEzSPa+K8jjSmFTCt6j3FVQv/7nHb+A83itVM3ra/+Wehp
b/VsCm4QuSLO4VpUYdekHENZ0+AINECxJQnz30vAXcVsctD/RURtJMsi3DGk4qKKtQbPTfqBt79x
89DWqg6WFRnnkRkxWaQ65XdjBFXEW/ahzg2TdiB4vVztXkWuyLGnvHsKTZb6ehsjKzvbYkOXU6os
UpUcFPt3ZcR1XUK1jk9TgJfuQh7cfD2P3FqikSVTooP858u/dbo9U9hyMZHJ4urxP9APbudinFHr
DZD3d4ueBeT1r1FgPJtApH3tS1la59e/RXr5FTkXHAQq6N2wMV4WhiAEvhtX2Sp+u+AvZJO+ES/o
iT0+39w97qbFEYykqYM24PSBlQU3aEMkXZ8CkIiKORYCjzEUTbxCwHbaX7bGI6s9On0EaeWS/Dwy
J2cFvj0B4h8QXoD+3w2j7bllmBz0lksDG2+x6U1tTtm8W1FG/K+OaAou9ydJVa1veKY+RzzeaU8L
mGZajbEc6YOYb7qYtS1wL+B/RCO2s+B3MhvG98sVgvSdQ7RraEpeYb4Gn1OWAobQ5w1UfyEQPLYr
tWFg2meBFbumfPAAYUbmPZ0LNa3fajT/hRB/XJGF9sANtO3BETj7oY1m+Hv1zBgdqNXSX6avH208
iGycT2Uopyipz4sF5BMsnagsawOAfGtIfQO4BU02PtZvSDRE6nnGa0inWfumNDwZ4G5Sa3qRyrhd
aICB51Yg7XZJGQ1i7JbdhsBps/oORAbx3m1UsSZdyW1p5z3WlujclpMvvicyKvGFn9uV2AiqzY+W
D7dvEJnFPlfAFiK7QkDrw7Mu+Zw9cM16rweDYqViYQuU01rSmRY8hsez4TpLKqdDHT+c1CJt1OrI
Pq4mI7lujfuxq1rxZR2RDgMtYVf6k+KY/smY6YCLuQkvfwdqFTrQtxqC/frknL2z7YuAQEaIANZj
PwATt7HwqtWmcd9W+08qcN291ReaFWIdfTaMfvwSWSMc4K81qAlat0GksFCIz+FVh0Dcaj0rpxyY
D8QLanhX7oDpvhIho5aTZOg4Hcnrl6Exl3g9YNNxmN9RyUG9EKXAPOw6iJzpYTWN9b3OR9crQdZx
Ji0cTcNUXgy+uVlAm4gdXKKsT9jx5tYoLMwFwIRUMtB0OeEtEe/M1FfzLol/Lxby5mcuhlsnRq4B
xhbEDXuEiyjJo1piLhkCuRnN+u+4SVl4r7Rvsvyz8S0vZ543f0SBcN9iOd1Fo3XY1shD6AyXUAzL
aF+DqxVD5xlEBOuiCTZmZ0DS3nwJ+SS5ITNV2mnHeVs2E1SWl1dAy0oZTotebY4f2i/faZ+j2sS+
8kdsxgcnxroTTpNOYdPK5wuY58SqUIRuCK10GEh3I0uYfs2W6IY9s6X30TG5TS4zZ6iMDP3njFoM
6K+z9gFveMzUTuYUpbQh5vvH4QgeNCqfxdZidvbMgTARS/7nEcbQkHowUwo+l+GVWTQroWMRxi9H
HxgJ8wl4E1XD/m/nZnvpmRi8yQxPghaLnsQoBujGLXSbbS602GRlPnMTusUFBl6rm9NVBTINafnJ
1Jsb9VbWATRD1Yhxu6kheJLq4aShJ3l3tGdDJ3vnAkU4J2iA0647aL1SnEZyeLevuxiR3Nmf06Uo
1r7FC1SxPNDk3P2NcTO+9YYTqwHx46tDLuqtefn3tWRYOJoBA8CX53UvPu9iMvYyqoeDwCqIxwRt
BOc8rzkGk9FovrlxLyHRu98X5pqdqKa3HMhrmRx7o9vdF1+ScVLb2bS4n/jVy9wKkoTXq5RTREvv
03No/GkrSwxef7zd2z1UDp5dom+ici9LbNsg+A2Sj14GRewrhAxTVfm+kLANRZtOacvZZv9b5bQ0
gx7d+olz4Xh4Xr3xrJmUMqhn8bQVawvqnp+35b3JmEU/J6daHuwRTXXfwUXUwIKWEeiBS0D07kI0
hdUxw1ZE0nc80rPqgnC8FZKUqURkol7W8u4+DfSjBJrLlJYnxiRF8pIzY40ydKaWFKbW1ZX46BQo
24tTE9dtjgG2OlkKTv2YlkcYY0YC0B3y+47G3UrgIqQ1fcFg/5QUFL/bPj4plJp5t+CqfpuMNJ1b
2HeZpFK7LajuMrnZ2IjT1FwFwH7jfw4dj3KkxNQ+ESkaGSSivtaD5Ae7R5Pv14W3QLpaLIuJfSlE
3S8wQbFQJ8pkuy0g4/W+ALMIfvM1OwvayjkorW0hhMWY8pXSogPEpE14tFPPCdgpQN3L1rgY5d9d
lCK77guDjvhE4F/EOzNvI8WbDHZE3aTjeCb8bGFbjALkcsqf3ea3WbSj+kTwO+bwA44PkqJAOkXs
JnHs+4CXbO3rF+8MDLHz42wGfQevH76O1O25A8dUYg7f9LsVlQtHqK8MIu7JeiHBs6q4ExSix7Bc
6vyWdtCGCtl0lbPlVeUMw9X9QH1THOODQWyuLzaREL2geWMBq7ZLPzoGPdGNZYj2paVTHxvrtfIK
ZScXmnE5RzKqLsXOeI/ITKFXEsNZWwFBD27xvTuOnXWR1DzfAGP26/W+Xxd1la7I9Tc18vKfBBss
qnQmcgWqmcO5udg7qLtfVROit4jvhPA7Qnwq6E4XhTI3Ev9LkyT6a51802/ul2g6i5Fsc0J9logk
cdgWMzbw6OEQDT8IYqj0oNTdHm+shvcbRBjiyKqmUpWJ+/RKcno6rx1z97MD8fPhaHov3GI6dihl
KmXG9NkK6RjtjhIJM2Wlkr92hoMAEVQ1QhrLPooedxFOdBx3lEzN3dOVKOdrxGrkAKz6laUFW/7y
7WeKyGabgWnJIMU8hfJ3FaCm1za/BiSLaBi1KYaL6nGGUd8EY8Yq1tm07S1gVkr2y1wd9xLWDY87
2yUNnZlu41CDTnsnwiUpf8X76ZfmjmqVYmSuQP2rjuabufveAEZxF6sltqJiqhIdm8Wp+zX4P/ab
yJGDbL1O8YsglRU1mt0kXAi5MCxSdzEEA6thBwVrlvBUmUiaxOvda2XfTpliU6AnzElHZKACUdYM
ftbRMbIKgc4ojZ170xI+FB2rRxfDW2eHz16ApzHhdiraX+XSDGDgg3okm2epgJ1MWpfZ7IuMqxvZ
yWnMlKCZfnWymiav2+zEQkB9Ykc/IXizFhUNKL1ZsuOCus9mBgAxY4/rrt5UqTfWPIePTLC0DHL9
krWtVjVAHW09LqGcFy1H+wYLd+UHqpj+dhXQbOjTCKD9BJJgxRUSXrnj3NcO/0iAPOCgm20Y1cY5
PJvBFDhaUOqFg8jtgmVf7DnIX/YT/yEkNNBN19RIcZ9Ofia03i4tyt1C8PRIffLR9kb3/otBFiVh
erLBBpTg+w/88TWOQM+oRDlV8NaQNTqB5KTRTsEScgMhOMQ7lur1JswhwUtnOUZP4GYjWlqtJ1Kn
WiGxHhP2GcI/3qUrAhz/thBjKg9qb4qm81hX7culYQalWaWc3LIqeOvV1ZgrvZmvJD5wvMpuixC2
TMyLw0D2BQlt8q/CFRcmebIg7Y+auBnhvVUjDkTJxG+Ui1pPCy5q0ORZt6nGduH+e1bPmyOIAisc
S9PsKlCFPPwPJk2VXp7dsXGIr4KWV+9kEzQhv+1C0+B34ImMXedlz+5mYMfWa/b5wuKI+By1VxYx
yloEeear34TiBT0oIy7iB2GJKQlN9I0M1xhnfZW85AOf7gcinDSulEU4skzJ2TPU3t+93SKVyHTo
/Q2pQE46B0V2ko/wp9zjljJrRcoImenBQJZ1r0GciE7yrgNMnpheK9KzwfJvWFxb+donFnxK2sH6
DETveyP/wrIp52sr5LR7zg24x3mS0dQiiSNKTEUNAYSsNAzT+N34eDHkI1UNd7QpMJGpOX9KVR4X
skYMPBfyfqOlmB0qWk4ZyijPqB19bhhPL6Lt+AWIM4HjXRd0pQ4CHUSotYav7VfuR036IXfWu1+T
bWmVIj0SXlp5SPObxMQmBoP5xEIOobpL/dorW1PhDMpgQi9fSV/ZbCoI49hWvKqyQB2/Uaat4Otl
rKiELHhCxlWU6/khjvKDZmcRUvpRmWvBuDVHEWQPQYg1RQiG8yN6dG4YIkbVq2q2VonhqFxoGHLb
7iab6OQ3lr2ewiLAKVqfn0U/kTendvJdttBQb5WtMibLNmmM6cF6V9VamlGqEk7kFYlwIhO1rgca
TuUmVM/cDHapjDL0vk2NlKRqkHrBKsJ7kju+LFkui5pNr6T13YZd28eOtb7FXPVHTC9aYLT3iawa
qvLYONbpHi5PWeqd/8hL50UZypMjfyK8+EHEYgfPLsOBEnjgPfBAbBrvQ4w/k5JFrFA+socy5NBh
ewOpCsMdJte+sPuqjBo4piRICh8TzAJBwWhvktTW8kQ46BHB+0kaUcWneSpcN+H5fB+arSdN/Bi+
4KaRY2IsPhji+RfyZwapAoxoUOeiW3TO5VVNjYUyHHh5y3Nn/m//8lfVPPONPXMu9FBIX/jKaN0O
yqzIiwpBw1pv5qGw+/Iy5Ig4LuOcByuOkpZqcBjHJkC9PDUYGydDxmttaDWfGLykN0WK6rNm6VRh
ly03K4Qo5uOysf/xOOxH6ISbCXHTH/hbcsPudLrZ2rs7orn7/xlm04TrkpgqJ1yxi5MgW8WGwzUi
aQSN3qAwUXHE3DFsosd40OMgM94+QJOkHGNP0qUFWxC+x3SA9uOqbKiN2YbM+lsE5F/wwoYdtBcX
zhhQ/CvIahAVNblHx2uqppQ/X0x3Nb0GvnFnuY+Hh5Rk9Pl2Dn7bCttw2n+tXTKdJ5k85/BxK2nD
ylSgIsRvxGd4n2jHDYF9uXiUJOvNBwFoVZnciOTHdLiVNfsqQUaD3FEMHMIZUfuy72zeY4w1gRL+
GsdPoH2y+9buOzoidpKnqzWogoNnCLlEhDTAkx962yuxYapyBNDsJccIbZ46mhyG9f7Hn6sNtQrx
Pgtjy+6ICEA8A7/UE4xz/ArEaL/cbdg/F3SEEL2Jb9aYdypzuSB/jvaSNruCqA4cPUktig345qXl
VhsBAboPdOW6FChXv/q4kFAhBzhlC8Og6GM55CfRjW1h+XvhFioUq2n8Ts7otKCnDbZoInobLIZs
uLEwUwbqZqn5ieGgwr+oikiPTCkTIOgn04jdGGdhvsvrNUmysVSp4dh1KbT43jhcNPGcvm9AOlSn
G9NdaO/ckTl97WmevsQpOzb46z1+iEjrhYhimqydf/3WSOFMMZa0dLRwCa7/D0lJuIDxC1lrFhbR
9Wkh1oMk6t8PsqvAP+FgUolzUWyOjtrJsYsipaGmYXiFKl4hMZEwJUdevBU7HBomKrLhEDIUILjB
RjrfQAX2yZhpfitmH3rWjmWTk0T4PZtNxn9ai1PwfAsS9cuCYFftV6kVFDu0jM5xjeRU0Qq0Axt4
4dugEGh69BSBOAZceO7Bcylot8ZMvMAhBMoFM38DvgWSG/NTExqNKgsilzKIdx6wA3PM2rZoZJBH
GS2oyGHnhBlGpeAHDNQKGPMCz4pJSLqPi2eJtwkxgLVd+W65SAEf/hsvpUSVDwJaRFOB8y/GfcIz
jWZrd+u6NNyhh2N1XMljVD+iF+YB+2mt/I9y91zyQ/0OEf1+gqYK/vQPOo8xitcdBCDr3KnODQbc
ad7N8eHoI/6NWJcGtg0Z/u3V0pCENIgXsProWySOqX+Pg4o+sGGYlkyuqQ+WRUbou7ugzhHMLdRt
+UXsfiVNs+tmuPrK7L9vRsSa/WOxesij+EsiKojXvoQVyAY9u4F5wXmiXz3ZgqdvLcccB/pucTef
ygfpj3Cx3ozp2YRtuO5UxNj0v+m8fr2aHzQ1nNMchDyVpja0R8/XpQtYTxe/byT8VuPZIL0mGbI/
9MbfH+X8jIY2KKb+373usRqzlwXp6nexnDO8N4VELFLoHD6NHLCf0eDe08RsS3rahZA3YJdcOx1S
Wt+2K6SfI6TpI08KaUAtU84Eja0kTOwQXxWAYdU3A9h2ymlOEl2EqP9vf/LJ4DG1jSJdPy9LvXep
htwPMx1LJ28mJem4FHXI9f338Ejw2pxUk68XTmT5JTgSfynEsrvxpy3+66b8rQetcNPew2RvfN8z
JZhoWDh9+0OLBueAKC26nuAWvL9gp6XII2irwm494RkJmo2rY6ZV3k8W77VZ2h0EpJL+VIETG2Wm
L8okbXAhLf8YkREAvxMUFz7LIcqR1Zdo26veQMoDo5CQCCQnkOBKfvGOGxtuMW5PZ3Zy9cyyqXRX
aVYd4QPXvVGKTkNyNfMwdDOLjv26CMyAwIMnErrv3pG8QyILeu+pNmYT/RWeTsycsan5F9vSutrv
gjxWb9qHk+6yf5HRVQx+gndRresErEWt0TpOlWwBg2gHUodEJdJ2ykwuqKR67xtS7tITt63GgsHp
jqpIgIuA4oGAfKaXmiRHN7S3VdmZvstJwCrcgxY+VACtCpCRw4EW/NL508yNivtTVyi2oqwH9wNe
h4ekKHjxQ4wbRn5acDZ/j/mGArnQqi8J80NK9DJMG6s+3NAJMyCMu6gu7X3w55YsdbqU4RNLt+Ci
vQM03fXLMoaApDiNtCT8GeWv+AjuakUYujL1OIPVfKYXtN1XKVk60zdkVaFOI54Pn7HNHYD7cjWh
8sUnKgtw8K/C40wwZ6DnJNFjn4AkfL+5XYayV3bjaDN5viVPcLbSJzYq8WERuqfAe/D5FU8UbaCX
lvj7B872B3qe0YidMhbeG++ohxzVmMcyRfFwLtbriwf6ty5AofRzAPRZmQkfTNgI0lwyt8b8HYc2
MScFqk0Ewm+90dZn3+slyc6lAyX5q4vAHNbdTKqDlxQ+/4wSatfE2Ewqh+PN7LEodUPTykEPStHW
rcSE3rdbuXEEDW7Cg4RPfGwzC8wbHW0pkueYHHdmS4OcM+3nnz8iVO9OBk5sepoy8FvOQg0G3NiL
oAQt6234Ji7OfZfCwBIpdreqtiUNYUPRQHR5NbcV0sJv7Pe/eB9Biq/2BzMsh4yVmmazza3rDLnx
2TPyrxk2Iws2nOQQolx3ERW/pKc4Lf1t0xgtMEDrTGWzMYioJ/LGfF9M1t/lm2ocXtwZPgLXke99
T0yc3Dc2KnGyiOf16wVMcr6nPqynwG5OzcNpU9dz7XA6VKJppOXhA1ru9JIb909FWRc6An26MMhR
6uSEyMwbxUKXDwmPxSwOIMZT/z2X/I0tQGfOZ6peLhkvyBKuJOphaENd/fYni/oc4tL9lxWx7k8E
uGEFABuFvpvYNUhX90Do4JqrGGg/yONRMh467kxkqYy648Aq2Mty6NlwnSJ9PPPImA5+OTIk+Xcv
Kkma0PLboQEskUvmU584arZ2GprwvEsEo9IInMD6BN0Z44xF7PWcGtfdumtmcnvR9ZxCEM8Lzlt0
+BBqMy4Rk1zd12be4BDMX2cRDrFUvfHJod43l7o4gugXxPBvTpWzWcVpm8zI9yjxKKhpELl+Yuxo
JuzzPOr/B+if1dq8lv0If7A/Tx3cWlng/mnEb1119dZjqJLdJj0L4GlWVglXXRoj6ip9sQhLBniw
hqTcjKoHhe6g4xAkqnsFEOpm77fpYyb40Hrm033ODol5yhmq7u0VhLgM6H2huowka7pQN5x7DyFG
Zuhu4VHfHY3uLpQhVGimUvc3piQjLB79klxAYegphMPqHAbVgcRt//+6PikDSVFTi7PheXtAHlu+
2EATLEwNk+Rcu535Sg6i/Cf9fJ7ecBO/EsOQhnisZ+zAXbtxfEPTsih/wi5Ogk0HPBnoGIqpWV0V
agQgsZYtHc1MG3AXRxzQDkP5ioEqQnzvrWfnnYkU9/jc5Mm2Fa76JHV2fZogajDBHdyj37a8GdPw
BkBLd+XLC8jG1s9uVX9oqIh29xRQZWU3rXGi4LhyVXctBWLaPJh7dUsmcy3AURo83hgJWSvZByZY
UlZ5b6jRpv60/VatByhGzwXIcfA7zz/73Oq/VGWktpAqYgNzePb+C7MlI89UvhbUdO/89S4enAFG
yJ05/OLuLxN5PdWRP4mVs6Xjn5Um5OCHA/58UkAD/xWkWSaIZmMGJu8A2SXxX0nCWgWr710zn60R
eGZze9ZMpGdv9kAUX5Vo7Iw4PUmXJvqFiyvBe1POUWjU874TtdSYblkPU2UlnyezxY61t1b2gLP+
Hr4FPFSW/HOI3qzzV9KRhhHKhHXXJI2FzV2NFqoW08W3zWaevMJxa7YuPtTnB626dx7v3N5OQUyI
cCwFIU2mKEjHx/pVAwrKhuCAtdCtnLKe1ZxZk936S6e441kCyf1m98ZZJRaAg2czkEjHYePct/GK
wGpz0EIZXVbexh9ZlcpDG9v0Is3wgiFE1faFd1v9OPsoCLYbDQ2CDpdCBl0d/eD3e7HMRFOV0C6b
WHJxB1RIx9E+k9JmJ1YxhVTsx44z4x+l3inX6DPI32+D521U51erga/wPye0d6AHf67ATDMtHYQC
ubS4izE6TM4SihxPPfliJ6+2u/pkSvNqaixKviJZhvOVpQE5stX4q51ogHuXfSyX6BIBhWLlmCMj
ktGJPaHTMN2k94i9KGbE/eMzuq+VfTr6GA/UAIJHtsYP3gYdmgiIJ4ZIwvlJlivnaVfT8Q3fEwB6
FptjbBwDXFQ8awUr6FeqSIzpmNJW75OdqS5iIaE77zVS55V1pWhGs8H9QYTKmhoSW2zL97Kv8fNk
Ccpuc7PukqlGL6up+W42ekYnYwI2jtxfA9LD06VjKf89Rk+Kip4wKWxMCO0VghYPffUGBvIxYJ5p
W1lxQEnFjjcHWUlLMGHOCFcMdd3HRiF0LdYgt73nu30KSqE5icK4gw4QW4wSKBae9Lgee3W65tUV
fsyR66lViC8Bgo1XnyVBxt1hPxbiY5lO8Q5v1lRg30iVCw3MTC6IJO6k4af2xNV92YiU/+vunFwy
VuK614PT/2R30naGOl6D+5w0N8/0MzO6xSBFheTzRqnKDQqJPShBNXD1qcIAKS0rAuyBWt9ImbnB
4uHWQZG1rdrqfl15eTkIT11imfiZwffhYEP+v+TO0+wXGJbXDeAJMuGqr3OtucK8aMoE2IEPXxS8
uYEpHs2OAPlC/jIjExaz4f+OZ/UrdayzX4wpgdl0969PptVWDUyDsluHSNWRM1AltnDCL+mhYmZx
hNhyNmyo5tBLLkkEgQjMXEQDzzyZxjkiWJkXObi3RiQ+LSZnj6XfiFfn7c69XxXOvEGAKstn4ntG
easAse96bAERWm0FF6Rof1DwLTIoECDkcVTGY2oz2tAgeo2cbhEOR538r1QEQfZj+3zdMOMcQ3WN
eAiWtpPQ1rHkyntC5hpb/9WdA9+fQArojdmCp+5fVGIVrBLXPvhrQSI+ae26wGx2AYZ0XlE1MHjk
H01LA7+7WO+qz+orUIeg6apwVPwh0VdSfpXJy8clgRsr35Jh8OmcbTrMqmd2nHV3BOymF+HHoLns
AjMYHNnlLsWLr8Pr45l81GoPJQ/FU+RCIodMTewGyzl9SCK4EUUdQmzkFz9lvOMEQjdSKsvqgI2x
JBosAjEgglMcvYEBxbD0m5rUmk4pK+q50VNmgwPUqPpwQs/EKT4z/cwWXVUtauVis7Gdy0u6YOmY
n7ABER/9KtNHHqqjIj7n4l19exN7qyVoF63pzVf4tbWGB1ewXlS5uxNmYx8pyBwxC1kipMKknGU/
BjrVx3sBRBqIaoiECD1Voa0ZEeYR1XtF7ubGtIz6DMqC1ZsbhR/478hI250aVlW4eBaGDUeUzRXp
KzoHh03Ibuc5YcMxQUpiNJ+VRHv7T4iwRkieWEDifaF81q+X7qK+F0DGoXDWSJ8esI+4FFOL2twP
4HwnmWtj4xZV+Z09nDbCFkUHKOmlZGU8vFvKzldsr2zXxG5uWWlmwewS1PUVygxn4eki5CnAg6pq
pI2RkNX6ivVOTHOSq/fIgD4x7WADIGK7flw5WkQ2Nzs+Zcev55Ghlzfi50NrQ94X8b8i1Wm+7zrT
ILqVhDFMZwul18kGWeAJ/l1wVJbznjRWJsNFLOYIS1wn96ZSh5ynPEyoDea8AkDHLMOywpBEtDU/
yGR5cTQj6M3eHGQIXwWaGbm8vqxRjxsPssaw78Wcm16d7VVMdTrs4GpAkd7H3u5klpAYKSdOtCAG
hMbrINs6tNgqNqP3qegS5rWLXZmnzye8Zg8ncDRXW1vE0CM3O0rjiqVZ9IBfPIiVowZWX/SKAQDG
PdBX4EaLBsDjxuiGlLpPbeDCKQoPv+TsbjXtmGmMWhgKnPRRmBvVSosKT+rQ9UKMHITzlis1uUvw
K8NAaEgrGYGRxcoW6Csm0K3bW++Trm8luHNJVAQmti1pOl1dOWmWDyVFGchguI5ojMiy0QAemV42
tMv94LPOcmuhVIwj5o95643JYa4Avy4T0c+GRGI2+jyJ2mhS9aX0WKtC31eL/+CVBNM/4lT3yhFL
Rtd9G2k2F/K0rAz1ACPkp27B6XL/BANX+1BPoukgUhB8UalgmawXD3t1FUYe6RowXEV4J2SlE3Mw
Q/hDGsOPzIZcn2YyN4njZIYGXhou94sLhtcSf1YZ5rrEHAXrPKPzpugJiL42Tlho3ulYCaVB2M6I
TYJvgpQaDKhab0RLNjKwo1fxXwXqdfQs6zg3cm1a7Kr9JnmYw8rR6jDsZpFdXdWAmV2u99RFI+6A
ULW8DGRY68CxqJH7f/QpuRKwUoDWP/MSbS6PjNBqI7jtcJkKbpFUes2DIFyiyQkvjNSmVWVsQnX0
wzsksb9NS8Bdk+jpoLXPQz/hr8bKl3R2r9fE2AELEZAAVfD8wbiT/13P7tPpkjzZz+CM/E4yeE3m
+CaD+EhQHlbbU7gEuRjsEITNED7JoUGhUsIsEyHV/tzzCP0f/ahlrlF5t5VzJ2pk67w1zoZaK/bm
a/EjGS2Dppvg/DTHqgrHL5Agl/9vt/v+UfkyEyAF35Au45fCYD4+Qs+xbKkG4Nfuqj9gkJTqFkqf
SPk7p+hRW/8A4IpYV/IT9M6iL2s62CEPGFOlC888ZgWjkDNxPMe9KnXkx7amjwiXgLmMAgoGUGKh
rPK/jTdslDTaqm+EQm62K1bZL6ofUAcq2nATLzcixJdI5qB9FjxK/YAwjCVCJ2tyGG0cEvq9bohJ
aWtqP6vOuhomNkcx2AnrTfQHN4PjtLydaIQVUhV2TaABfxaVh3TqnK0Oh7CHFmP7dvPY60fBSNsh
9tek9Nunyh3dzFjW/qsbr22j7JzthNzixQH7Ai8zP9oY4+jZ5PjJjNdL1E1ZFrboQ2T8TXXXd2XN
ghEsV5A8Kj8SsOufHCOCcAIwEZmkPJLPTQHcK8sUv5DFrQTsJR2hJTg2NC7jHZqiN6h0ibL548BI
aW59OKu+zlNDEsHYkZFU3Ik2wYJssXtpKceYFWY1UyM3xwI9wSRniEt8edHWQ088CVLJ489Wff7n
HpTwdlmsD9iKsVSmjK/021RLF+9z7z3Mvfy7A1tTic05az+XDOtt5h+D7meC5a5op9nth3bPi/dq
L3V35zIqFnsBxIMn0O+/xdxDcwPcrQIts54BfHQP6mKS4c6+Em4SeDOLy0ZveRi/W28XKWoy/k1M
OIqbTJwDuHBCy7NQ2mpuBE0wSpsAByJCVqNcZz0xq5UbAbqK7MhmJewpqjGepYyzGe2obvOugnOU
5yPGyY40nS/qPWS2PU5VrrFqssRtRf0ltDpuzZen6iATA47YALkEej4Kfy7B6WKwS114N/XZyEkv
nBWhT8oJsrcdwH28jbxHtIsqupo6icbcwkt+wOJIIhfLAT48jtEC6NKSOZjG5XjhVfqVfpeU+Ylz
0eytDOWcblPW/Re0Gw4PkIxGDv69RBv5DnPKr3cyYJyiKS/VYw94y1y4rUBZukE1q/72ZegpqGay
30HQ+KGXGsWCCsimSMWrso644/v/98KISeZNPK4N8H7zrdU55kMIn6Le4szfPCrAvcn9NFhvdwp/
feBRV2WQeVq0GUUfW1LaXS9J/LCX6gDmZhjD+ILVjIb7qfLr2LqArDS+iUWx40MDvr/kEh+GkK5I
tM7lIKgnLa7JwJVRjPYHcOq6Qhce47Selw8hac7yrl0h+d4NUY+D/zzXtNBGOWytQGmLVzH2oGEe
t/Y//6A8uyGRkRXcWQYrjcWQFxaf4o0DkwheeXAVMTap7rZUgjExMdC1wHBnSiN3V1GAJdPEOG/2
hfMj56ZvmNZAM9RGB52+91rOE7Il3KPk/d4jheOCIXLy0QNwfbG9clq9R/39Abc0HtS8ELMlXEV+
XSj1ZvvClW1Vtm6zWrxncjxPiHL1cWEdoxovNATFs0UPBB1mLZ81F8z9z4/7xURzSUK8ZGJ7yZMV
xB9Xt2MHFFIF7IEv3BDUE23Vb8H6x0Z1BMtRHoJ09QDdQn8jBz1oHdrhjoJiKZDc4P4O7uozKGWn
Xx6GWaH31Agd8HGi6PDGTSr8fXzGsT95fKGgWja0xNzZGzuMyXCGv0J1oKu3Lt7HP9ch5KgPKFxt
sU67Vo2lMZUT5pH0Sg1doqrJThwW5SkU2HpfWW2r3bzvAYQHuXvKN8pJapHjQnG9HQEdyLfEeAXk
zl5M/NmDH0I7VhfPqVIsXz/7Y90zJinMBzhexqeOVscEMx+SIYMBFE+Abtb+p+xSb9p9bdgYHoNz
WeB/m/xNywqUksgLlNLBB9qQW0z1dILfOkyS6+aLbT0+aVx/35xCK4Ss0N6V/gxnFzSp5v5LiUIE
3JySJ021pOO7d9DySSisVKa6IWCQVDri1dO7qo8ulFfZX3MGjmFIQzIDNtEQCi80aFCv4FGAzuab
GCmTTRRFQmvdOvWTDbbG2EIibz2ngsb5acc/lbvKOQLg3f17XC5TjGEk1H4b0BBNAuQE7P7vQTiu
BpM52jf1Z4yPny5Abo44IF4IVhFvdo50PGUMij2pLGdujFVeQZGuJlul3ay55Ccxyntni3tOpMNz
Bdpb5z3E6SYgB5tMR/Ph2knfIIP/xNA35BkobzxHazEBx25BAqSH3PgPaQYZIpBwNjTfXsYHwiET
DCepmjHc98tHrwTOiaRNXJdFSVbwMqHPfvRJVhSxCoAVZiTKI4/pW8YhvanaOmkO+PFjEa7RQoOB
LdaGdrWka3u06R7dR5WLs9Coz7/YOHDqhqj5rGIPgKvLskCYfAdM6Ni9HjNf6V7625o288JxNUcA
i13l7SLkJU6nY9Z3pQHzAgd0YjrxPONniv/dYcckhclLrUw5lcYICKWAKEeKnTdhG3yradetyf5l
ruVRqQYBWmi+i9NjG7XVR4gN2SWKmyKr07VkvcTcKnjDyJqS4lPrHvW2qLTdt4vas3/LMcKTtWPd
XDXhk+Pha77XKYq8HGZVDyMM1sUeqbNeemxizMYZvTl6OraDrP6zpSQa1SWvucU5mp1ZxrDSrrVp
c7zQHEcUIz+Uf9WE0o+ki36quE7qN5u2KONWnzaqMH2LEP63Z/3sXEmbz/Oy5nP74ndBwU9gcT4s
Q9rBXn/fHlt3jup9UmLOd5EYKMUg94dH9ckmVHR6DyE4eUsv5uFY5xEmwWKkT7aVF+thywy4lrh/
9nwAGCu7aLsQyjeXfW8lo1PcoHttYPDmST+6Bzn7wPfWR4y62WjCM8RzvDeIxlxQ7WMDO0K2yht4
uFYJZfGkEVWLADt9zoTbIpAB04R/UL2wX4PeE2kUyrofh8LY3WO3sgxVsDfWHt6kmiRNZxW6WRAe
johkIusA4uyMhK73dhyb86A3suZWek7RX7GKkf2hgERt59ygiIh3Rcp89exVQRntrK8m0BIl/1vb
VkmsnHy57A5cDz776W9MwkRbVDQ85CaoYv4bnaOyT1kabjnyDf3Qd6joGXV/v4mkSQfz2pwdFgV7
ulKLRbpmawM9R0Ncrpa0522GBewm7/zQ0pjmvWzjlGf8b/9vnrTBUrQQbtANLZyvIesbr2nEg4Lt
pp3q9W0nnn4vrtHgk4nyCObz3zEebC/RViNP83lQUpl7e4MghmGwYz4ztpdZZKlDoswSe4OKjRz3
V3daXIJF0B3Ko02DunCkv9Pl4/D/jqMdQPVKB5LJjmlFGLgTjms6ELkhHhRI9WQ2ppYdR0HnGGEl
5m5UIKWRIZ6elxaW+k0W7fWZwarpQad3rdg3Kp+qkqrEQ8O95Gw9+FDPi1pbDa4cBRjMsbiOUS8u
0atBmON2XLu+42cvse4bQcTneRz1mnKVT+bsDLpv6hLbWvydy4/xOaGvHNIN3CmQlQqyCOvSH2Vr
aD21otfKs/LSOf50GLvRbC94y9SLUGEhozuECtg0ClHszGvf5fbS22pRCSxsYUcCLK1NJFeZcGiF
8thUXW5MqOgqOmnhSse6Iuna0yMkKQAw6VU11CmUHDFUTOFcYAHWG99bADXXSTgpCZ8gfE5VK7XB
48WvTJE1C4xpwHkEYlHV8oG4Hak7rvK1jpcILaqthl3foGfaaYcap6PWeyujshxzQhsUk2d0VaTP
qP2KzxjjloJXBMxOsrDxWlgSPXfA6mxfqu+A4+7kky9WghYBzP2QOraCZ6w+CPFaVR7W1HU+AwlS
4dV1onXJYpl6+e6hWUzenRTGQOejSGFcVnxhQEFRw92trFSHwwiKqUztzNSmTz521KZg/biDS1Gx
V+AMrNCb+fmRZFVooJ9Rel2VPX+2OwsthfTd+Hyb9b5NzMid+nHKUsfVPczQswD2sBjsq4QN9br9
YB3zDsx9q8HOtCScPyohcUiI74jwobg7zR3c/tZ1bHlL+nFPKlISD/G3UeaQ2BUIBUTPfBKF7Psd
iu/mSHiU0o8NGAv4cp/MJa2bgmQA7/sb0fOREXo+nKtW/V1wJhoA7B2VjXnU0Rt07Vw21t+7yRdC
GEKFzWI7q70x36LSJcLo6wioAOv6Zh7jaF6+AAIRDNdkDYhvTgE6U/1LSrDahJCTER6ypjkrJwze
fLx2LL5oPXemPWiJVNgSl/3xe097II6ouUl2hAQ7HWxuPJwTq9uh9IaXvjbIpnH/zD2kpPow23Ax
AFdkYjhlNzi1Ky5MgMzDr9SGNrWtmb1kuvjjoOmzo6OtTCjEgHG9NAdqPSPKUc1fJw3ePdx+Il4M
WcSy2dXuZ2Gjco1amwUgGiaF2tDw6jUs6K9580FeY8tDkUNB9H3X8iyclkK+fXEbJiU7x1PdWJGR
onrIZ+b8/6g9RtvoEwjdbbrICl+V2QTz4EK/0BEh2n8Kq0wuqXY0EAsytfTFVHTYRShRIb/tZoeV
ScfnXzRtAToTwSjFcGC6ZLJjK2HMRpoL4FYmD+8gDe06d3E93Rc8lkF5hhtNpNNjvWZlq9B+nwXP
GnQGto09OWUu4sNaGjIhHSxz4df0ZKm3mvl4sUw0K130gJJGKzpf+MBn/JstqOzLlmfoJlW+nJ43
2Oh/60iQi1QyfW5CKbaRe/e72SUfyZARSPJBOE1rwaXcLjzGpXwxqgKfgyoEHFegLhOdN2MLnYg4
fxFcaQ1ag0NntafHZ9ChDryvsy0xAhXjapeYjRB8LyQXXwcsrAirpXZEbEV7R2gtNcUQL+wCltkV
kbQZNYtVN0WB4teID+tcBIa1MDo2YCl9qBquoSgfRQJJQR8TWver6rsg96W9ZbUAOVw5B+YpZ5/q
3DmiKJqn/CAnA1tx4gKGFA+/1h0Wjryg4pqxadOo2oUCgQLJYPVf1bexQ/ER0NKTDKL4L79xYM13
6G3UDuBCo9jOnc/UdxGpSn8S0O8Uojl3N9dNtbUrEu6mHnoOhxCoADXpouN6U6Dpip1iBFtHu6sO
9dh1G+xtE8XgVXc6uq/DVecgwUM3XnJZ8MaqPZ9iVm7AOzMI2QiMBg1NGQkijnYS5fyvjh9vxT7w
sREpR5DnZJwi4ly+F8C5KWMVLwUfUrwDlk676FyPDpVqwQv1f2eCHtAkb/s5gYayZYMamLKecpIg
lCthHUzJwpnk/cc3RfszoWylRbVI6cCpb1+XpRopEh+LCjxf1sfPSYfOSxysWAj9hPF0+vvJW6Ml
+da5cOQHqv0rv1wnanDo04N/dxeYkvu7OBDl4R4M2Y/gWPdq5UtBeAvAsxv99RtF/snsd+21QlyO
Dt4WhtnshrvclGKAX8a2OJVXGFpAxSvTyUVXcmPW+VPOyG2z37e+dC3AATV9UWfeD4HCH1nngeqo
CD/mZ086fXD8NoC+u9H2nLiemFP/9DoF1rOucy3jsf8wfjwjyPPgZbQE3Q5r6+7/W3NcHJXn94KW
QJgBitmjF0FxaVP+ZJ07S0JUck98feFY2j6qPaBEQfFkTj0gDXdoK69P6l8lrL+ciU2Q/5tmIr7x
fxOJRSwN737oF1jCbiNnkg4nv2JCAYWUCL6LRGgrj7/6u3vYMTcibauHhNzWktTmm0nFtaH7UZun
Wn4juhOQcFNfyv3HTvRgdc+4FSYPLI/1doHbdyB8uDjYCeD3t/E68XJJCckMLucHQXxIIPPFirFI
icT3SlPhI283HguvUJSQxaFsPgNxM6Qe3m7MPfY+qmKsBpmI1Mdkf//9Tjeo7lstJXu8HY0E0/A9
a00cTu45+23thcuhx5c98npKZg59yQf6pjudYP42QKcdp9usa6xzeuQ7vRAdV/DrPXHifXk//W0h
nSVf+rFvAFSptwDXvvK+CQeA/QekHgl6kWfpuTWeGLXO0YchFLNv9I09bTkglmb0WR8Y04vCXgEb
dkvP3iUhkjfVEMhho3pbUZ0TMl39+3vgml3WRWal/e+JbQrDETbQ7wHqNbTPGKoftugAvJRBgWQ5
8Qgbha1jeDI96Mu5L+qVvhZ3zwczppl1i+2PdngPwiPPZ2aOt25iliOZfrYQLsMcRdLaHvCUnc2k
676xo8K7tDuq3G7G70I301YO9FbvqcIMCiWuePCOs74p4yp9dJN7+a4WY/aFReBFvcdr3kJWrKS/
IrxPLSHIJx6/3lhyOyUXcxSe6oBpt/QQJHAsVzHU68MNwxpReGY1rjYpIragdKeq3VEqY0F3kR7T
w8P/VNO0WQlpXpbfbDtVD9wZZLy6fE5VVOKaTDykZn6BmA31ynBEjHLrsRYvCa279B6Jj0Zkv2Qi
wBtGmcq3aRW+TB0hkdALn5jS6GO4Ql6grhz6+0QBdNkDeEoEHXy+bLIXvmd6E8bwuz0xloTf+Y0o
tEWyGcrVeGSNsamJjuFcBTNriMJRQS5WImHPBn/TsKyzXzUbhYd4YKia3/oKQEFDjsK4y1ediwnW
1aHAFIgP0vdpXZc0iY11dYUrFJZQ6fbHDCpxIbMizyMo3MYN/YCArAOA4PNLvv2Aok5qIPxnVW1K
knjwcbzYIuXHa6BY/N1MpK0ref4aWQbTY4fNTPU4CMCYSF6+8/+gPTSR6/86xW4onRvhh64dGus5
wBgiTUQ5lnIzpiIyMlJ2BWDztbeRuI4zPxIvVPR7jf1CYTISC0Gte4Zniym8TFkfCIOrPn53MZBk
zleGQb5k4+Udt2hRPjPS1yGLucbhxFQPEGjl+JYIH07kce2hoP9n/fA77OksqyMX+fJC3OLNBGax
p10sKKmIkAyQ8ZbxTZRT9gjvo6BU6VgBnJcueaD2a+vj/ayXYEdyAa1HSw1eRywO1xUfnD8G9UcU
HoEj+LGo0nmznyLNN7Wy1S2zdz/pAkexyHT10/9LpFM5rW4SbQEGavgVF/m/Vl+jXxD2gU3eeraP
DyTmuY3ANrnMhd5k/pCI4x3fjksZmTeSg3v+EQM+QesdsHqEMP5vwdG3ktW1w5m8XaU6kK76zFUD
Rk+WdmwzKAQSLhnV8gKR6PVFUtMwUcG5WxyVSdLV4UrRIYm1Ms7oV38UjsD/ibOGASbeC6F247r6
7THo36Ye9rQ063rz8nN4R7vXWGmM7DAzkTystXwaq6RJ4LXarYcuPq5MhlcgXE7foMds8yLjswnJ
zEMPVuQTCDfsSta3jJpsi+fxTjDJQh3lU7erEVI1X7jH3tZAmFDXRXB3/bZ+8pwuo82eDypssu0Q
qzohQ0doKjdfOOP2/7pl9DpnyuJLk4n9WIoLudvUK78A6nN7IjLVfiu2by5GVlbks9N/UqF5PfAX
RUE4fS9e5YM5SZBpILDWZdQ9TlRF7ba2VJSfnMU4ja6at9lTxpDCHz59nAWBMEgNKnGC+R0n7zBr
Qld6ZhTwaj+lusAu9fLVo6RY/PA1ti3r3BRalYtcFMQdQduNueM1RxjXbHraUwmP8vnta6t2HBQv
soJJySA5rFH2CEmVwzl5LvGfcV4egQVkRQkyaJ6DFNLPGypin4xQnR5gSiYyhQ3T/Ow1cQT/WPhL
Mci4hQToIINmve0sSer5IqEHrOMMqqs3CnxTUut1XdJo9GVBdAS6hialQrZEq7CQWiKJxJsDWi32
YZq83i4j7UwH+nmYTxJFM9pH5h5lMDSWUM3xh63wy0M6gFLAgs1UnYM/cmzNAMXX44l6+ddY0t04
aELUY9iNqczqa46LsCswutIXav/sSjpwDyU6MIc/4nz5aTXbIQSYhgTeBFQY29QuqE6jOUFQqEu5
3YjCadVAq9IWgrS40ZlI6BFaHbW9mdYTP/+snL646mQB+LEa6UBw+blFThpGzBr9f95SeRaodwGu
FstEJ56x0tbWdENJHPCu7fWv5aH4JsqrbyawMYdYDvot1f2Ahd1xIprKrvaTcVPfOZr07uDAtvFI
W3DfuuUjb1gd7fIZ5+ZUOMEUzL1/HQHOl7RA30b/xOiqTQpL36L2881npiL7O9GLZnFZbYig2yDH
BPBE/5T9BZgLNo3AikcGn/6ubC7b3yPsvpVVCOWzEhgTcmJAQh6NTDXIfcJJLLXofMugs9HT834G
yCir7cmdH+Xck2m61lLuEBxSDK1eBST6z+zuyamBTQshCz3q+IUKsWy1ab48VtVxX/IO/Ah0X4pu
v2Rn5sa6INs6gBptJzHH+R95WPjgPNS4+66taKE1+QzlT7V+B8u0+8sHBIt7axtNs94V2b6UmwXb
vFeEcL5DyXtjAs+5GvOMz4b/4vqL96DPs0hihxtOlmg3zEEhUfAVttmaiJdVvofG5Ds+1vQGB3Ns
/WD8xbRBAcxjfN5eBRmlBBblINt+zd7YikyvZwOpNvOmetew/c7cJy8PHX2RZG9aPTSAQ2md3D3l
fSw1RVeFKUqKH7qUT3XbBiNGqK4udFaXgpBa6Fj6ELZD2+bwP8xiKD/dCbk0L8Fv1xKTwerRl6+/
niYdTX1w+yRNuKz5XItp2G7cfqJBRddpPQMf7AljSNug4pIr2zBhMzGlkHiOimSovlS7XG3gmlzR
U3O7Uk6z4zGtvALkg45l3HbD9HyWOpBjLWTEjaGjyxmCoDQ/7IA02LkNwUfFN59dibxq6u/uynUw
9KnFodzrq+iEEezWILDaEqd0Vjgq0PROy1LekgB9JaaAKD7sgs5D2R6Hi06Ejo9SsepMC9/7Drm+
aZPhMC+FdwVAzpn+qPwScsRNG/zyq6jkZJP3CfELh3xtFGXQyhvs+CZXqrarXZOXBEa9oXHE8JVE
/7lZhTvNWY0KHdXLWgbdMXP28XGANEvMCVPSc6+EEguJN1hM0BVDt1IHU/EF+Kzv84THKE3wUnW4
DZOoLGPWs9W13s++nK26dYgYOOWJ4U5qJ2609gBtMPzbtt8vQM2uleKL+xO7WSyzHd0bExOqfBmM
W5X0yj7buAySEnuxBniSU4E/UhgOdzv04UvCO1OMzefXMMBCgjppNy4mVwdADJPCjMqewIHekQyH
NIPa4kN7llei3yTVrSWMr4pQ2R8jz68wnWQpk/e7dVAsbvG/JHSppK08JKYXIkwUoiOUwS7RZdf8
t/fiaHyfwa49Ou2KyPDNJQw/nbhVLxyMmFUi0le0NCcnW/YvtYIcLyc0wQ50gZVGgJLNdKbZCqvL
ucZshRSVkoiDwXRCQ+QbYvAY7gm9bQlpEhOMeVvYztEXBUrOuttwl3kQXjevGeKKiJ5xUn/dcT5v
WealdpRo8ST7BgI+U9aFFEECV9aOcfFGp0exacaTyNY7Uh6ZIuzKyYoQiYP4BNFXfkcSrBRODC7W
/YuoChU9WyGmSv1lloyMeHLF3VKtM9ubFrNGPlK4nYugTdtiFQTGZH0ZYW/bmwUPg9PS62jaJpJ8
0jBigInRgNW6LWsCHhj5u4xrfECMjZgHXxgmYMVjBwpMzxtxNI9e+rXyhQUgLePBo4aJVCarYp/R
0X7aUu+0B7knqz8SOse0HzTweMXl+s8fIOqCmFgxze5XhXNF6SbnORiMPBZCD4YNU21zrkO/1kVL
uHW6A3xvmtQD1cIN7Zp+PbejKTil6okDqsRtpDGc6G6zGBvPpHCTT0xwyipjIBo2HVZkPbY3KGPh
cxQCxCeYqtUHOyIGfVIjaNZ1Jv9xcvqZ+Zg86L9Pw2RLstHMK96jV5HsiQtjR7/GmNtsTXbP3rkz
NcKpDNoZOr2EbGj9N37+lKpuy8NGucPsegkZOlI3xiYPkkwb0mHQpUg3H6fpjSD3UvwchszUA4Lb
zIadHBrAIwl1H2rfMfTW3q/7lvfe//TqIAWSo1OLWeukbWC9ZdF2NFP9BKkam+BL2pApJqpjMbD1
/gCP+ctvtdZjq1aRKZ7OhA+ALm73HjTwYQSzNxGT6vfIi64NGpHmhfxNCveNils2dvDokNnOLMTa
W54vIAiazcRkr8lQFMVv2IGr98rUCijmQYOVfgmP8qi6fkDlkWiWNZYqUK9YHrb5TP84OeBQMVs7
37buSXcky1BgixacYiyp+8HY/lNdTWrGRUQdVZZZgTLOpFzzR3k+HuWb8XmutOr/wScSK1t299SC
1xrwe4DVgel654HN51sY0AbKcyDri68rTU7CqtYdoHvayMjHEILxAcdaU6x1SvQbPR+QUxksKc3C
xNeAsP3e3sUTKyk6zVfOUp9FwJHn03yW1dR7FN/rCXej2y+xvV2YfXo7tow7s4n9bZCOG8j9yWU4
wbY48edjORwKUBLV3yR74v+j2idPok+XFcr06qfNkPE+cr+Ii2h/yHawwOs5yP8N9p2m/bCGysZA
kvup9DUjhoqoGe9VrQH8L9myEcDFEA6p0nQeWHfGREax0ErlyI+To73q067qSjRTYfUl/blxvaPq
FzQ9k/kgq06La2enxjwMN55y7oSqi/H7jbHvSASjI/emh8TMy6YyzY2DmFjdYTIdxD9f23beHy0d
lfMovOPanUGO5ID3/OGv1SV2FrsbDhgAp/5eT0Ju6QGZlmNSe60FvFMAYHC9xVK08I5pIFOxNU7Q
rgPki1ZeKaFCkJfpzKDl8oGIZVmmLMqzXHv67tTNSLINqtH7cE61gqC+qx3Nrfqyo5rCjszlcoC4
S4mtaEu0JyJ7rR4v8KAUXP3ZrcChGOk0LakHAqKSQuEYtfzOuwR5oyVgFkEc8bRJlbeu9UOxeYQB
jRUABmHDrs8vxqWYPLj7WAdtwTKpBrB4BMaAEf9jSPPCiG0ksJS22eLLUCe5KppMsAcmIdHqSxM4
x76HbB8YRVvyMB8ZRUcm15dOTDwOsYEZR/gOaRrXZGndcxEkfaFkKdDNjrVRudgXU7OxB4gLDhkO
m2alaHoTogh1QhZRvrsoeSylFnPtBAc8jMq395+j4ZhHV948p+Na4ifHw6kvNJTU5TNNCpmUhX5m
CzSQfR6+3w5h/VAqszwDJms1yxP9OVxuMvFLCLI76xwrlRo/fKZAsP7FTadI+yAsWQhZmjH7f+V7
PggVLyQUuNA6doOWnc6V8AU6AKDUoHEp2iMYgqWGtbqCF1J+ebweNEvTVQWgKLegVM9jc+Jc+TON
QVHVZxRIwHh4FLjE+bNArF5DaH5J79AQgx8DrW6WdzViG8JIo4DHNLfUY1tmaccKsCJRDQM5ZFW9
7GUE4ztlh5ecPXzP5xovs/yeMMuMnKWJ8vyYqaEZAuxTKGGgzZR9mLhJ1Gdu1DFz0BUTXQigA323
INR0URizc/rEtzzorhkgNYEFNSvQjROIwMsuRcFIlJqV9ecaCL7yyxFiF83jIMItSa4KecIKI4Fa
AD5dgH5x+dVpUy72fWqgtkybmd/8YOHbYMETI5bycUcnjXjbKHtor7aHy1cgEwAxwoxLJiI6M+UT
8W2rko08K26ZEBVyoZzImsfZbyc7odrIuGzeAv21hEXTgJyXWYUuCu3AySINwxwGmi1pyEqTy5do
1n8bxnS4n/lvhyzDa5bnoJXEMSU5MsUb50YFUEck7xLfeuE8Rpk4jOXazxPW8z8fmo2VO22hb9ss
J7biUHOAC2Wd4E5C3vxD4Ra061CrTug+Rkei2vTtYoZ2f4d0ADVG2uEckuLNUBP/9JaXtZyA+dnY
faRVinO4WfvscUvLCeJnYemOyB5soIszpSMCz+kOOVnu/jAG3cO2X2l6lbHEqt8Yo+XxwOuTZ73R
wyNumfwlWhkOmyqSznwjyquNxgzuz/qJLroFSoals1nYn4aJLZQNOMf+oyiiGaU11dfuIWMQ48rA
jLLuxsUrRB4ZazPMoeD3KOJmeQSNs3suyl2azHvLzlbew27vqiHcjwbl2CFY4jvfFgTryBJuVhDd
c2jXi5FoNBzeILP46KPpUYTdQGqQCwugDpxW9H2DIDTOnVLrauJ2AcXmTBlDx6fHelH3o5uomGkc
RSN9H02wCxhq0LTgiuLqwe1C9mLRslwvC+6od9Yqm0p9O2YnvXzi2HXfgY64WvCJsCH7C6sCVEek
uUW3cKJzRiUQ/E3wIOi0Wl4AxKFRGiqpBSXwYad135PGL5WPoQtDOggxKe6KBGu/m9QFz9ShGcCP
O4uhC5pHzX5ODpqEGjCmI3o88ZeN/KV7RdbTkqO79CIzHXUyeGkXzFK4aRC82jGKSSrO5HHl5NAl
brgr6rOBe3Vlsit18lgnKbK3wStkSDBFFtxhb1a3S2AFb21szDaawjgjYtGB1xiBJA76NzDFzMYh
jHPjKGkztPNr9d/4Fjx9X1n3VU5plG7SK/n5bXtcKcxkQJubxO7Mal7ttw9/6cZQCmLzXpNfv265
l7XHKc/fDEsJnpm24rFv2NC/eWQdppZfBaNauYerp+gmKYhiF0gx0j9AxYHRWAiVdOOSip9IjVcF
+dQijO/bEwPoAsjIwHreaaRCBhpEcZ09Nq0WbfmKyp4FBcIGfZ0RH2IluWj1/gpL8SgN1Na1mYLk
p9cl2eKKJjW623cKGkFBChObseMi7ua/CvS9GQ0W28WASFXyo0PpkiBuJqNLMBwVw89AKXZ8K4Hn
9aO1Ufltbz/ivEJkPKTtEIN2XDk66iKeAWEBOa/wHJLreKgChORMD/N93N3LS0z0rDA+nZ+v+pRd
TJs8dlgsWEYffHzdAH7kDSEKsq4FcGRuB/xoNnpVbD4uloW40HEqY1woPVbnISfcJ6JggOfGl92H
Qa81mTugCK6zYTZeqHuDkK4arXsZkwKfGAUq9HOIU1iLUb5N5qjodHHK15wyKdPx9URyiTaSJoud
KwpdXjMeJ4ApR/2XErOgbXpiJEVKll2zjBor1xkkEnZ8Y5RDIHyKGTklmNhUZ7V7Ero/nlXmQX8R
Ouf06lDXbFdz5n/MMyvct8UWxdLQKvpug7is1+FfCtFpHcZl/Vo/blF9o+uTFPKTVeqLOp1uD6xC
p8TzXGo6CveRs2zyYc3v5cbDcOhPNXtbbBlI/kRiIObAyu21bhAMAEjLCUP+Bu5TNdmrkqdw78Xz
1y8ZWEpIK+ZOneLD3Xxrh/fD1F5TwziDpZaLGFhhIDaN2Vng5xMNAo5Qso7XApBfN6D3EhF2rwvf
SwAw0cu4rJ22FfgCB0TjrDlLWXJrnfgA18htUqoEtbqc2dZ5+Eu71nNCeeMEmMK+RMwG4rd1CMu6
H0PYrbeQOVX/K5WQl0TDrap2WuFfqfy69kxdE2/qUUlN8IsDEECd0+DI3/ordeuCkK1RtJiYLmsw
ewX46fu49wGpQ+inKr84rvDLeUdMu0fq501wXcbhdtNLY5Va1MxjUBSM5szVGeN8Vz2V+fEZzvy7
THQ9j2sjwtg5HQyW+8nLOtQ0Gq4Lnmgx09beTcHPDDnA+PT3RhH8vzot87Fiepplx6QuxIrsAsAH
1pIEev3bZUzhOx+SHEUZLiniWU16tEROOg/oR3H6nwY7V7B7AjrMf1zzrsJ9UYuIY397b1/RHDrA
e7qIPBGHVN1vrFS4A6pSxWF1w7Gb9isAwvrM82+dTMBNgGj/2vHud82VSp6ANdZMLkBrZLD6ekIe
5yS9k/Z8NYKkIKV7U2iy4OZplWyMRkhJWW/nWREoIyw6psskhRoDpPEAfCDaT1NX7vOn9DQmiZLy
+MJWL2xvNhouGCOcvweKQLHHaKsPVKvgfjjVFiK+55ILj7jQjKbV7S9r7EOzYdLlwtrEi8pIHLp7
2e6zEyv4gkUmYARPQqe5ZPLd0Nkl4WiQHTrafe0UDjTV9lNG8eIsoSxdVdbB7MsizbnNJATedjmB
+usSXudWoeEsBhnsQocWOMdLz1HmjHfw8K8kpKou9QKa+SlmzeXR/0jlznb0z6tn5pHZL7jH5/AK
yApD00tZZh0GaB1zUv6T5vU79WHysRITwS2Ckmvs10iCcPLu1Ht0zBFSOxDFoOrXa3QOL9HLBPR/
fpPOdDxlhq7dOcm4+Ia0lBar6fEmAs65r1kFBTA08L++lZuycz8+ymiUU1N4xZQA7vQDA5ei/hYN
QZi+n7k3xhcecbeX5pocSBFlDCU+czTyVCJNIPDRm28jMGF4NkzFhvMerIcNnC3wJJZjZHPdZ7ru
Y0CyDsu4fmYMrn03n7HHiPncnvNqeUuQmMg4WSRwQyUOTemGtUO8lOJhMf+81O89ZS4YSJx6qnuV
na59rryU0/+EWiz24Zgwe+NoiUg3qBIvmNtN5u9o0unEH8o/o1FnqExE5zN/69TbS2maI2eg0Fwz
qtGBrJ3NRUkikP2WY+OS7gvnIY2jIq/4m+gemdDmWqa79eYh4eo8fmb3LuyrnyBfmrbseo4OzzeW
y9ly+d4Gm/lfOoxI2PAmE0KBUm/Dxy+qmBLBMUQQ9X5jBUYoiYXMVDLVAgWEi4evWvR13gbItA1s
UdvpO8ZndZ2cm/1IMpkGXsJ/Cin+HIpDM3lLMVU8tAsM4GdirTRahORn08A2ldQ9whdu1wi/AiW8
Ol2yyT4Tsty1jVJSUZ2dOCJiITnypi9lMvuTbCxBvyh2cSvs6TPypU4/nlgfOXtbx8xGtzEQo3Q8
7sQoRqs5GVBWn/7PUpxlNwYhZsVVEvPod4FG9Naq6vyjn2dLBiLKx/2PBYPY/s3aQZxTn2JhzqiY
nlFIZOfjbctCQsPVeAwCsxSqER26vu5QgN+d4TlNDJn9WP1izeu2BQpCTUXSM6l0lVPxCf/QtD5z
z/5MApvOXsBliaP/bdNoo5rvP3vuambGcm4wUYZ0EegQPaR549dlokt7sFwqg8OvG02UACHfCTAv
/+lhYfKpH0xJSuv0EBAwt2hRwIt6u3QkT+Ht7ZUwGfn6otBC7iGku5fZ2bSXOubSJfdf0R8jiOSL
jv3uTntD4kCuSONCXFfGMr/NAJXtPhUrcR910cNQkYUzh8iplp1PLBOi+UZmg6rxq1AiWrWg7qLQ
uX3+PBz00/uPmnzZzZWZsn3j9/pFMdz+KuI7SdNseR07pcWyVBXbZoDOyl3u0gPf5+Hb0/LTpSqT
aPAo1Y/+Koe4kvOiXjJ3St5NsbTzvhAaEj4Ial0TxcbkM7vJmlVo/ecdYa/kLUzDxA7lOhGVrbeq
+7kO5JHJFOHEna+zzfgrA1774I/KnqjnReg6SV/o03KN6O3K5YOR9dklq7tcQdPgeTe5TnnbOux+
udWGkfl8cTNR1yb0tX+zQSWSLT6CLy1C1pif6SrjtUT4ydn5TGjv4IiYiy2sNXqvJsOg8X4wzTN4
6XXWNQAQTXMKEFoVhifhJYdY6+s8njomT4VVM7JjOloWK5y4sns8bLE4HuBba1Xa1tfx2IOjoIz6
HgcTOqxHIBajxzok/R8jjmRVjeKY3vq6QPJ40FpnQgN2ryuhrieWeo11zoNMRY9XQkIrjanD4EGq
p8ZMyBQVA0XEInZ6fWk60ULZtSXgiQGfEoTf7SzcSdkdnQew8tRd5BVQkQl9RzRr0cH7yBVz6SA7
Z3JDPkkpVl1UxZDo5jSzZ/mXlpbK+MLEDc5rgwYgGA4Nb5IeZT2dhYEaZ3wO86Rn38q3Sib0tL+n
Arf8XTz3pwG8j+ipY+MAWYQ3u2Y1sjY+jSpNPauFfU74sV38aQ83U76JWOTvWeDADXVdzZmRLjJT
6QQ3VQGQGvLd5Xits2VizvKmsaEP9xH+/zMlot7LoW5/qDK1vtlSCfWaryIiauy19NCDoys8nBEM
/Fmz5OfcUZ3yoTERCXT/7WLXEFesD8CdtA8IHHHBB1iW+zlnI28/8lQKiBFrXXBSbzDmBfyy0wLX
3FJThBx9L0QjsOrxBb1FptVO5En/MlUMecp6UOVlbXqXrHk9QG++XRsKE1efC5quDQTZo5kp6ASc
qTG4aKa6IUj//MSfM00XMoIRGIQPVBw0ExYnqA4Q4b2hx/hXD1eAQn9/gkLdKGSY82Q3pa7rzvJz
zLBgvhpC/1cqTXXqD+NCSta6B59SH2YsT2LfH9geqxZkafnfN9D7+sazalPVPapeGBwEiWTOHokT
wx8irrFLOiDR+yQcQVEiV4UH9Lb+LNoXWTVacSBFYO+IqB6cnfRCEJy/x/CQ8LlcrPLb+GrzSXxV
TrOkkI40e4nhdjWbDJG0LOwyeWRqXbi/tQ2I0vPrmZ5PW8mrU5qr0nzLIqTMjBmqp/160WG6/MjZ
6g/z8WoD6cysmb0KUbq/n6C/LAa2LBWjn46s0YtXaD+nmn/SGuAdECxyTi+KNAf8C39e4nxSN0y8
cS0O1/wupKfsx1v/KQJnCIakl6zsX8fEVsc+Ycqsm4KmcVu9UgUvhYKQJV4ZskaKRbkjpX40z/pL
fy3pqBwIcKgYQQZ8mHNheqpUpuKDiehuYFrw9el1d6YSTmeGB5cxDea5L2wz2s/tGSEFb0Kiw25B
27SZFvb9LKPc8f2AhXrOV5+dX4fTgU6AisaU8izFrC6FaNGyzxgeIGV+ofdRRSTYQEL7pin4Mjyi
dSy7yjDJrtvkpSuFzybMY4z99WsPM+e/cUCVkr0kc45V5+N/IOBjTytIEEy59TshqRJhGYeztHeK
7PV5IsfWSKS2lj0GwzHLK6Xc/Wph6WaXNjS5epzE0krIziuX5jD7FcuhB8BdFhn10ZPNzrf8ZWs6
FIMAxty6FoaLT2WwZhYe3NYIJ17DyQ0kyav+fnrFSrwK9EoqiPCq2Zy8L9gU6qlcjrAHCnr+8ZW0
eXbkUU+IZUAO/x/TyRV/yjI4blZ/yCKu5rnp9RNFJrliNJQHbFWUwSNIp2ZLhZSA5W0OEWLJjIMO
uoGoaSlgCVIQbkF3/VaIFDaXna0MI0BKUd4ZmhyKdbTC/blBJXf8LAShB204AfnQKBj/pMAai3fz
kS3NDS7yuVNsjGuPRDgRT28VOeVoDYs9FPkZuQvuPep4QxKOKpfhwQjNyNb5zSPWrqffzHj292Z7
jpn2FsjHAJ206ZUZZN4VwDtQUcbVXj2vM1JHlQvzPCoHyybCFXkr8HK3WjPztg6PbklsuOa/StQ3
U+wD0CIRiyTRg2w6inghfmAYbV/rAklebZn+t1h6butAoNDtdtivwU0jqJY6iUl1TJmukjPid8Pm
Y0zOjBMHs6+5sJyQPglapI9afMcR0UPZNH067M2pXcz7MQrM7t6wRqiVhPndwu85BytEBydKuGNU
9f5ZFwChxHJ6gpyBggmmRqVXGwjwoW4aN9dpUQLNvJyCJsJPBW7glYuyXeD37qUph16+1KYzf3Gn
xtmAmOe66iEEwAkl1qSmBqeQQvcrufP2oqq5+JiVnL+tI2bnSawrdJ2x2ssXhT/Nh+vmSt/Updh8
W5tLO+gmJtLkwQKeD0q/+d7WwY0itDOTdNh74rwyIAhGUxWMJdpcEQuARhY1z5XCXSWAb9dUhimB
jmQ9XPxQeoXEOTPLL53YnYq14W/K+MUGB7jJ1tTTFfTz0wC4/wwa2MN6uwG00vX1UF9V9OWuHTb3
FjpaAk//RGyH5Gg+q9Pht2y0haUMAqGXF395MIVQyTowJFu5NUgscVlbGjE7F3p4otRtMoSaPoBu
u7bORZ2Yc+efdZNiZGMfumy5T9mMqm8F+pWFVtb/D24J4D+EB1jb9CdTA+VeJlpNgDI5i8RIWS4A
z/+phWaOnPp4nY+I4kK6aw3GBMHlUjJcg9bwkwaI8kSDXDR094fGEubKYUcfuYt71+yAR7w08d79
rPCmUTbU3J3vCnG3LT2LIh0c4IjCOqnoo0xud1RCxil0I8pOVWu9SbpMLyNu2Z0xSJp4y5v+uG6Q
qq5ogezcY6muBFUw1hW4udhxUZ13xfKxJMEwg/tcn6haOlN5JfMGwVA6fWygJ7saVLI0taANPdnf
cAxImgQTmdt0eMqczfCZPSBzrdbCIGlUkMrnQeNLw9KQGa5DW2YhF9vjPIscM+Sg4uYNeyEo5pFq
29maArxtbz0IJ2ZShqll6Q780OPjf3XBZN4nrr9VKXaTwQzJ35BA8qRP2TpOa25L1TlGrYDfy+8Y
VQXZXxpPshf+tUQoFebzSIa6TNf6hdijU0jBa/VP5SQOqbRBV2P5SLBN8CDpdSJvp3T+uGt4u6mi
l5uqiV8bGTcGjapK3+LjcfDVoW55y0fHCWE6nbeA5JZbrjOU/Ir686+nAW0vBUDc80SxgcNy3Y44
N62Wkkbisi0LweoEVdAjdsAAZlFgpswKfX5UaNyhCFU8MJ8nFQDCwXzb8tXptKeAI8hOXhH5zVAZ
vUJ+8ozmfmufZupOEfxHodi1Mr19j3ScDk2w5H2vZXALzdhVI/YDfvOCsWBHXaZnZPtZ4EicIb86
E6M8ibqAmPvxTc5h0Wxbp9VvzvD6ylD66TeCBlAG4c0AIWtghJ5MJWaSlsZdB3fQoOI6cQz+W3WJ
YM0UnhouxjoiWu5ob7vi7PMSXiN4uI99G+7WHjxtBYPRiVJa1yu3lhIpCUl1YjKMLKBCLys+9u4i
JL43HGs05SZ69NQEEGX1NQ0rTe8V6g5Bz1zHSvHNEkAI8CfwwucH1TMJoCmgXl+NRUCdQ0S3qqlI
ZPhKpEmtIdJr+N8n+GbNIBbrWA6gGmqRvTh4JcCZZH1BlFbud5pseLEAhK2XGqblis0xWDlBOp9c
5tJ13ZTgxFzlR+2MFW5qCA3i/T9eOPG0rIh7yYFgif6KbEQrEpXlmoUTM57PDQweCwqr7rlr7Jh3
GPLGFHPaAeRabOA0jL5m6cnt9UyYotWATT6g7uHynQlw5+8JCrf54IVQloGHwRpHWh5sVmaDaQQr
0tbAbBi2LXb9x0KlwHyus/ihbm+LyMgotRpVWuH/7zHY1im41vn381Sd4UWp4L2ei9D0faDaH5Ft
gXVew5GtuYGUsIrB4IzPW8kna30/caPvMsOax0SOt2iK6AHWmbWTCyVaOKH3FUvKdDv0v5OLyQAy
FQTVIsrkOg7S4e1vxzTP1aNqGe1uxGzI7iOsYnvaFnfiVM9BCWCQSvuVuaXGFv1vVc9212XwRHD2
38y9F7kKxR0WCMmw076lJe5uQr0zYlAi1OveJ+maanwroN5h9E8KPWbxF/1wR9fERlYkA8dGZDs1
fYLM7RF6Q7qfbkSq4J/56u2Neg3dVArd92TEIf+KCb8alHcalNrSbO4Uk4FyyOgh2ypaMrmYdCQg
zAVf6KZ6d6gSDilDMCOVYzxcpZTX/kIA+PC72/MvLEgqOTb9g2Gp4SbZSnEo3WgsCmjgZKbNhmmP
13Qw/cbaDvOU3GArzAhmvEVopakcXJCiYnx0TG1antCyQJhNSitfE3CBWoEzs5OSLj3qhILtB5ti
w4wnwcLgq2lyn/YfvxJiJnSiW4h+r3iXsfDyekleb+FWvt1VXlfPrw897XwUcFO3mDHIb/J3ijBV
xXOdhn+PKOQfV32ZMEZ9+ONMYnOUWo6aTk5VCukqp8D1Na80d326oALbrEjFCbzdfEGLaQzdwOkP
Ldr/y4L2VmHAk/Nkt9cIglXwnWZ/ZweCicW8UTmdQYkveTze5c/c/5c2Xq+lhiNmShnDQl1Ke1kQ
mAK8AHLMdf3zD/YUZLKvxOlAsVwSejrTGVs1Bukch+J+R1CMgAZsdu297is+MjxTN5gr8o/QZhh8
AhraXoNF2RaRXrjB7fxhbrIlS0npDmRbbJciHZIyKvn9O/zE/9hwm+93muUsJnb4knPzVBETHZ+K
SMk+bxi1KTIgD9ovaa1zOigi/zo/7HhflOFiHK63JdSIdo3wXg5KZ6lZQ7FLzKd8CAdp0bgfldt2
TeMrNGhB1uG73MijHYHcc6pGtxazR0JmM5ehvUEeKuQ09SuY4hqqWVHe7dZaoBhbhaYZrzs1T2cK
c7qyV2N4cagpTHdGHtp/2CS/f4RYLLuWZv+RLCKfUiXEv+V6o6d5aVy1XTuP0T7+gBlKjWDxMjHh
M6Y9vcXzMqcRQ2XoDx80DRpMvNcAWQyoDfj/RaZcMibS75+9Vt5g50fclKGvnavnqS5nYxhBBr1g
DSQ5nrJ/Ruh+ftefOvuQ2QUWPkATTfTiUvNmVvazptuJMlGPAua4KPE+9MWpegLF3n+RCiSKRH+T
m0glQIoudMqLMCy3KfYMtT8QXxKpna8yhX41ZWNt22T5ptT41fl0MFkw2hIQBk35ADilLye2GkBx
Z7hx3yKq++MJ6GeYfGm6F9uxbkbl7hWzKgSOaDGOrPp2GsP85G26IODwdNAvjraoQfywIaMwOlWO
CqXMIhNVuWm9ajpi4JszV5gBToFZ6+AharmEU95bL4jcEhkr3Wuq0Jkcd5cXh00SxVh9HjW4rDFo
QtRk4R3UI6OCaWwaZGCY4So2MPjtAulODZRNYqVlayqcm2XR+mfuzXd7rUHu9CRxYKKJJtSgyZN7
Lrtx5P8xMlA+wmPIqQKqiSb1yKOsYFtuuJcnX0kaBf0KebVZd/5PLK8E+2puGpPbsZ4Akoo4S6Kg
IpCoOM92ZNpP1RTbJJFH2nO8v9aP8X9IgoSMAv0tl/njM7cIaFAlnzU/1o/deGTCzoxdTiUuMrjz
6atNck0+oTYgiyXcCkvVDTdV9reDTj7JvB8lEU7aixOf7vNE/Pn3v5jcQ4uiJN1pergTd79G1Pj/
uZg7H9NFeQBe5sllR4MMNzEFlsv8gEWD0IOtV3tjwMIypt4WsOSIUAvmee2v8pOYQckTJepPXFXg
TBoaYd4MGNGaUX+e8NzKSd//mfRsWzSV2LRwNWrF0YspeuDWiuLDorsBJpEPm4WYmGjEZ2eu/rVf
WeOjtEMwpT0imRQgMfNZIYfe1x1/5hWrS53LXM+ZDgLJNQmcxu5OavM2ElcCbt/LyWhEYbYwqlc+
7IpQP/Tpe4Z6DLS1CBQhydQzccTuVJLtwpoVdy8Wv/iS5WYbEGZ2/QYsVFVq/ZJp3+m577G4ab5U
YVUjuy1qfdn3tQx5mAfkAKm/wLRISVLj4mrazNoxEEPm3xnlkPAYxQZahbjJhh97bKBOzYbzz21V
1GquV2CfFe3RniHFzpBKXZijAdkTjG+XXoZiOsEBmazs32eBTXmhv5FZU9vGypWlIvP69K2Ueekd
gLke5gVB5kE53HnEYN/aOWohNLcptj2WADhUmkXSXa6sE99/25VjLvMpr2ujPT1LcikRMBzkxO/y
7tpEOjDN7b5+CkszgfqROu1JiCQIuG6zdLC/xDZ/DaQhNgTGW5BvV0bSXQ3qR3vMyUztspR9E5sK
lXu29J9xbTX/8R/9bXJalEMoDPPZFhHL/pHGTYzzPYdak9XGT7X6SgJcOWm9f7X/6CCaNgW5FQjF
Z5PdEqWGylOHO5b9ggfb1ADMbpf15+b3ofAINxF+wDBU7iZzQpeZi7s9fukfGhY8AyFR+FD1bpRQ
KNdn8I/gJScTirHkF+XRGBjFB7NFS5s4vo7l1krXjcEBG6qjGnjCo/rKnhLWc459AfzZoI7Niyx0
QcwXDkNIGDvo4f2SOuuyNw/5pt8VVmWmPEI/XJYL9INmv/6gBUzvWvHMY/yyoJU97KmIfpNGJuC2
OSPEAjREwtjevCFZvj0loYdTPgHV7qfBsGnM0LOS9Fyt8D5ytQ0TH94e94KJrvjeDPQWaOhpF8ME
1yuLBr3aGpl9y9r9eljCCme0zjNloy39mCvryKopWb8gJcHc3I10GXPmQy93SBM6Lk8JmbumknBw
F3Qm1GnxTxIY9SzI+jcyhRMvs/ijeNLBJj2hSQZl4WDNn4IOQYldJrv8n1qDVY6um+/U+U8i02d+
mb0XhJY+K5CEaiQINbj/QHJ32cRNnQNQHc08uea/B9JWluedyd2+cs2JmEnJTkMQ/D3Adfl8nCh0
ZfAPXCHgiyRNzAqxVuKyd434z3ZdC+qkAMBjlU7HmZ7oIhSs8qHcxk3ea5jNtaeiU4mHuBqdbycC
SvVYQX7jq0nux50wir9LKNzBdWfhfwbQegZncAH2eZU4mY/iFYs9wwv2a5GuUZLT7B+g433xuNq8
MCoUMakIIV3T+8vnwJHmjJHyccmdlc2PoCKYVNRwC+M4ao9U1ZaMlQo4MRRgHY9yG4Oj8Rbsr0OJ
nSUCs2uJojQ8ctFw37LqMIFVGTxkHrVOCdKnR0Ab6DjFUnwPtDYlHvFrpthsZkNvqI8YBCtxt9Bz
NWNGOex5nG6fRAmZlV7stnyf/IitE33Dliu+sqACWOoTIwzOmXEGlviJD21k1x61Z31zwrcGGgK4
DyJRYihp3t6mRgOrHVG9E8JAkMuzR3s8rM17vwrlH5KxwQ4eGZnOBfVbdBPBB1kK6cKJEfmVVv40
Kfbl7PQGeV2+QNNXuQb/0rQsbyW6BpJuvA7HaCDoFwIRfv9lt5xUERGCVMSZJlbkvSF4RS1J7KcS
8bpy++XFuGByHhB2BIcM7vQDrcwynIYEcefJLCn+eiDNuvCsWsvymxKO9LzqbYvJoaH+E7B0EOGl
AgkvVjJaK05Xz8wHa6gIaDwxu5YLDlUNMYPIs6TBrqujg1L+7l8EY/qhCSA9RG3OlE2ym4TPL5Oq
mzae+UYoh5SNnHG5TQ/FJFxmhAa9OmsJRvDOPDUGgEApRO5D8Ox+qpSOvRr7A1l1989EmfShtpL4
NDE9rOvYZ6ipur+zOL8rCWpy2KbjrLmWJhw1Oa/7jRH0TcIpHY99B7+NV8djmQflT0CGUQorBTvB
1UmnEMpG0/JOplICCfuIGC5IBL9QmJrUk4DvgJPOy3swn1JlNd7/zjxVkuHbzg4IG9e5hDzlzP2L
jDJ8hMRsu14ch68usyWB/RjZqYVZ/79N6rhS/aTFanEYYeSA9Hjn6JZCwCNlPi8R2kXGe3wZWHsX
sBMMbCDegF9X20P9Cyc7Kixai6jUjDZNPZiSp4TtStmtGgOTOxaB8AoCwm7UTtdlXxllrlPu6QeU
iiBmAuQMY+ByoBhR6GnmaN4BZzfWxY/kCd+zh2jkBsAAQTnZoyF0Jq/52XzfXDFu81I/0/Nxi9/3
v2o73zx1oNbDb09wniR2lCcSYO8BA1j8NEBcGJWIzJR2atEiMIWzox9cd8X/Osjz6nAtBSkupnYY
7pRMS6iENPtM35XuvyK4wP4sJ1/32LHVFJa09PsXNBxgP/Yfp8b3CVBy3L0dBERV+PFJcSFii57N
fRxEP/m7p7/brCjEPZWFte/GCDGbxJzRNBqh7m91BbWVVoLWBOO4np6ur9ksPYtLd5sQlR1zUBKW
WKYp04T/y/DEU8ZtE8Et1XkncMt3dwgnNggCVIqLeeQ6LJUcef/vUaCIMb/9uzRoe7G62bPijRBd
SAMDPfP6pfbtAr9LwoxSaINIcXS6XwR4OBIfVPjNvqv0ASpWvcNYlP+/5FoSThvXX8NviFrh6+LO
fyaLnGbe8PJ5IkRLxvR/smp+8/5Y9zccHdkjwvPRxXT7UikmqaWTphkUNM58fN+KBRp+8+TjmD99
DLJn54PTZYFhvFJKSbYnNis9dp8xR6LCOwsNdaAApUHz98lYYB8OiO4QGd45VfNVrcmLPJeTqdOT
BYdEoHnBkPwgrxztQkBGlVCF7XJgNHjOKX6Q65+0uKNV9ggDBd5zeXp8qgsqxh3N3EWSoId7+esm
quWjhhfLFn/2BzzdwgHUQq/OwebbxTFYuOT5ynCk20BOZCFD8C8rAM90hK+UT/a6+OJKR8/5gqLD
LrSNmSmMMIXaPCOPusKamtpPnLPNIOH1nCK87RrUiHhj3dyekVJLUTkpSKohzrSk/oWPul4GNGxV
y9s/RaM7OhcEHFE7er5Gk4xdz2uQXI5odevZTaviiOxPJXDvxn+OrmRdGOa0Q0afPqHCi84GipNq
EEm4CnUt1AbquYz0wmYIiLevN39MgiwB9IdSPrLBOWjwy9c5bi7hpOjocW+GwMngVuSI3RzsAn0e
5tC4zYOachMhCFxzGLmP0CaEFrz5HCA67wPC/dcfrS5Dihcxh82hH6Ol+wgC4NdL7i6s5zfJJWyB
VIBEnIM5SLaJgZxpo325z4y0K7RkxSExRQi0yw1x3YFMJHSQLBrPOf6o6nO77LVhTJAP3e5qgmAU
PGabhuOUb2hRrY4WRXxDrydamsS9g9D+4EyHNUKTuvC3kLmFJiKreqZvv+MND1m+VURfMY2F//4i
yUS3idZeIC3Ofgd2d5ep1YUDw7rRxFfZ9tEmKsWvYovnZ2px3+MsYOkoOndovsnZ7+pX+LyLKmg1
e0GiNdlXmeI1sg6fB8jMxa/Y0acfcpDZD8zI7N5BhZavP+H0XHU2DZuyS66LMoIF+TEzfTSQwUgj
ugdaEuq4haUYMCKa86YWzfT8SXclpFBn796TYHDDw7FXNCEvPC0tqpQ/Jn3oOfzHIgHXct2nPndJ
njIPAPJ829sg0DLtHryTSxalOLTZgoHTH4DFaLoDbsBtanyUrM4cpSnUtcHKudvMbfLZFj0C0KbI
at+65j+kk9gH7HwfEcw0X4ZJ0sYiCup0RBPfs/QVo7M/iX+f8vV/eGm9ySOwoCApRabhvJt2htMK
J9gMVT1kmef9tiuD5PGQ/Kl7Qo6JBKDvACBvYYqYVoQAhXnbTwFE7AiMKSuHxqKYDP6iF+hT2RgB
OysWsFX0DycxVqkO310DTLH4khG9fo5BEj/0hcNNjzZX6MgGc6uUEfU9ttnZEo4CeXTA/nk0r8/e
UKDqwluNnan2gLmA2lAJ1rT/2I5qgctttMxwxOPsViPgKtHWMRr/A2JWtu3/tk+HgoP5OFzSBe2h
aI6gQAiaajMtY46yq1Vkr3bQH/mzAt4fzZEnHgKaYYSOc+05HeMzBauqOtTjbcHHYEbHGcVzVnrj
BY+S5z5r6rzZiHXBRV9Hb5zGRgysMzTGczrQkUbDIsJAe4F2S/XE/D5Hmc0vPGDWn7tMRcd+g78d
wD2v8pDhYCdURQ8yo2BkyI2rMowWLZsjG8JXlqmEJYxz4JJqRRzxA3afd6u4MzJDeXOq8vNk3G+1
YtMtYGuQRF3nkZQ6RJPptsDdZJ5aQbyJkWt9NImQx2mQI6JJrVd05qsHDauEB3/Ve01+hbDvkd/G
9wuVCGnRV3ZPtMTD1d+qgwSrfC/r6bLUrC8XWsogVaLQ+EyN7Y9tMWt2v8wMecn7iQspgftvES5o
cgp3459qI/cKyMI3E+mQsnLz+SgALVn1hFHHCnNyJHqsr2cl0SpH4dqAjTFqcif3qjESB1GyJssT
QkR31h7/v1aVOgDzY30AzDRUraQieed9AR39wa8FWRsCshG/gsCxg8F56T6/nPrlXFPPLoL2B5NJ
kbVo+ZxTc7mU2soTikcQxMO3iK+t16INpazntm0fnjp19mGO38QxC8L62hM3vVgWeD3tc4sfYSVL
01T1o64xHcU7V7klY/2rfoJBRq0YTSQmh0QdsRBbJVGAsDeCqDad1HO6lxm/O32V4bdqQb1qbIOB
VIIKIVtG/j9+mcWVHeXI3JOViFkxxspH0CNdrE4Xb0KZcDUa7dDMtYuwiUwL50089XUoAMcSUr2O
UdUhLvd89/GwOP8YZmyhETUVEqopMwBtqzMHI28kZk6msGYe8rE5mgb+5xzb1ykXJ9NSRPCuZUDh
66mZ+HmUDPbT6qNVdqOEtJNgZU+oCK9ZMr7kTXNKPrzd9iLUzJKyRRZFQKnjDQcoY8OfxAhRXkGD
0bFw/XMXYac7pLmBs3td70z8DI00V6RHYnjbN7JOWg4YssU5MeeWbl7HkuuQcXT8zEl4tfxHyNwr
yGm4cT2opLfcQ4mSxOhyec8Ivk5J/MSCPYdGVPukozz35erGF5EcxqCRGvu8BVXmHbLFi1OKcrKL
5uElzUakmVws3B7ISNLJYE8f39CAS4HP1sWYniow0FpRhHkKTPEWans2QSh6iSJrTU8VFeRsuBO/
OFGKAlWDzozjmC7MQDXbjuJOt3gd+6EB4xeEZliSRR4X6T5ArKERqgZ4vLW81Rh7wvBw+Eo6SfQf
kBDmIa0FoNqS7KrSeRldA8i999Zw6DvSC/eKgVBpRvqc6kUNMzPWXJ53MbP9i498G5RcMgK3E9tZ
hV9uqtcUAssVl60vP8nbRlUgWlR+eVJHflUwQRi9yh3coLIKZOs54RPigvEtLFzBHTtEI20sooUT
AmpAdeNzMohm30ZBiGuaGErzYbETGvCmF8XTKwXXLdG7h1Xs0m1Z9YzcpdbIq8xDm+wI8agmEPM5
PZzQz9uBlzFuOaLcT6ti7YX/128VeV8aBhCOFLU6ejAgoXXFKr7zhlmBnWRO6qthbx665zNnkOMZ
r0P/tDp955HvXgBUa4WNx+g4N1OkrA7YsljkvLCd5BfDG2HxRMkDVoSo38aK10qVhq0BNoK9wT0z
FZjeiJ1g7dqLA+vXFKB309FNOXqNcycewyDQGzhCjFKBDYa+DLcVQVzHhKEmVifb/bA8q+AwVQNk
g/qlCrsfvGrabOyOEnBlAHBnABu7DxskJKFC9nAyXgS9/R62JfWlj21JyBj7Z8REX5Co957pwBYd
DasezrXpsCmZwkMmxLyKvaLE+M50uKo8lB6uBzUdUf+sLOco7zcqbJ9ltts3MpscXZpj0ZDK3gXg
jnGo/4fPUMPvlNjP5QuSf9YUFICw4dF1XRBN9EP0A6jafAiFXErHrOceB//uFaLz9YyvIb1yStKB
1AWZpjqwDDmfZVlVG1s8ICDPHCayvPqzuPcCTYIfcnUVAkzLggrnh1DKXpA4NCMYDcHC6YdvbKoe
wSikTg/w13KvonmuHxyn+hUvpoYWzLyY9T6pSQumITABSb3afRqQMbP2B/xlbhSRUxykB2pSHkLg
nknur7mEWZ75zItXMlCbZeCbOttIZ2VyqfhaFP5cddnhaoPyAFuzIrv5wvGKMeYyNiLG9z7n0PIz
mp7muuFmFp5FVD+0wNUxwq4BQpcU0bbl6LZVoEasEvsP8uwZ1NrdLlR7uwnPqLHygOyEWyv3DsUF
tnNwdhDKHv3Fk4+gOcynByA34YtRtFMwls1/do3nlYc+ZDF5fM6nZ5lZrzrQ0TXZ6lIws/9cBBOw
VYZMb0jG8ItZ1dwY22tFyjRzh1jh3mf+wQycfahnCfZ0Dhd+7F4WFW/0MIc6gOSIAIJluV/fgmn8
9GNSiIU6Mb8FGGS7NmttgBHkP0Dp5IKuvWlhaF17PU+E5jnuLaqm09Y9740HM0Am401IDOi58gFp
YWOM4Fcr5iOsnb+FAdg6gQhvLLjRpV5m/UJ5clt6DgxXr3ETuHQkgpIWBp/mFxuobmhjKqviDLDS
g9niCFFhtX0qbeE0Q2XjT8hQkwgzl3R/0BtqAsL2s5EkIZI8PaPllPJGs2FF/RmEPF5D1owTXv0n
dk2s/OZG+14ejVmLwxUhjhP8RYS/vRk6YXKLWcw9W/f9j417n3yiAW+cHGIJywucWOZh2JVodTe9
sSmzGXc5V2rGchpeA7ygl9fxk2ODrmGv74zowUl7Yvga/a9/NkFwB/Lw6eO887rFon1JGbN1U12F
0mgh3HfCyCffMrxAKPuuc+q1sJoGP5j/E0rsGis/ilQ0UWpXaslMnrwNycogg1hilbMTylrP3TWH
zE6loAbrDqOBDWA6OFn0Kue7ZVbRr0MaZfF6M/FakojYowWLz4z61nxfhQuZ+rZksXR2yWUm2V62
JU5Juk42PW/37LOuJMzoUAkiSgsGA6Ff8+YJNyrnONjwMxl3HNJMHYlfVOF9NsN6/Y0JWRnuYv0W
2ro+xphufGSi6yWYHUo9opfwWjSqh8m/tYUElhnFADgDUBmpnVydskSmqYiLX4A9XDyyxmlIz+0o
CTNg9vFmwd6qLDEzcc6GS4UeWrl7n0TXz90T3ek9vd6YGGTHmddssVczjQupwHj/CYMEg4OhL37F
IQ/hg3b7qeQtaPVTJwLEzBFPTk85dyrhvLk4lFIGQVRtw0EGMCMJYTJPU2qz4P15PNHQzWfd13Y9
gfBeHBNsJ8JstNdY1ynIjUsBg/pGvD5U7R0slIO6j+BIARW4BBNyuJSwyMrnORwkCd7HN7g+Y2gb
5EvvODFt5/vTrqxR61jN5lpm9nJCEQibXBaDTu08STjjdfRvUAu95loByT7BOFJOXcZQPPmkx4jF
irp7jUN2NWHvyqlS07RhlYyB5dTgQpDRMhiUiuysPLxwfxesP6sXHF8ob1kXuFNc/RnSZu2ybEZZ
1XdWPuyY1n80ASaEW6kCJjr+Z8ZjtM0q0FU3Acds3z66eX00EItBgyvj10OHHU60rXq5uAvj5kQK
69/VRQORwcinNVeIF6gVa8AgZdWricTzJDygfsFAlsZWiuOgIP7wYVPdtX03qeHBPKqx1I2pm9wG
TT4ugmPvHjXKN0YzTKJrTVsterLzNC+kPjBQhIeMr2a8Pkt9mWa1m+AcJtcYK1+6pkgERKsAGaPe
5pTkeSPPlkIfNLOyriTbHpb2/8QoRztgykOzlM8q0+2v9QGUfzS87vXnbu1MrMpvvfv5Yh3S24tt
oPTcHXaTwsG0E8stXwL06vcAAEoFjONl3x24O0kVEIY43qrYKUVaxEp8qiMam03g+wPPlAoB965f
EZUGHi0iI78MTxuAzBaxrEMw5JLLXu1/QNT649nAq4y6s04KkVcz5HyO92fNYolE0rQuqYDuWxEV
l31p5mMLpIqGuuPXxK365f0EDSfNSJ8M++K00tp0FLYAIyxeHYGP9haITAl7K61srkAcmof3cErW
OdqzJaB/HB+ZtCFBtY12Znp0YnXJZ+cuNA6rDg92/Li353IkX2A0cIjmER5ZF8pLrez1f7PjVqx9
WjE0yqdq5b5Ofm+MzxRtjy7cSqyEptWuS3Apd15AjHW8CqgvO6JQAYQSU37SAMA0LHRSG6WcXSwY
O2LkOMPXlkqRGFGx1OfscnAfndiS5lZC+x00nR+NMGMZWhI0ELzFOOzEzKH5tBClFRvglyJQInzH
KsVb9ViTlnK++F75EZHRRtGyWSyA/raykF3bE7INll1QugYVRViYOyfTIo9dVB7jpWOciggf6yjI
hgP8bU3N48Pm7ci1iHOPptaNTO4MsklzugzDQvjTLYv0O2Ck7PgmQYoy4xM0HIvwV5tm624AIMc5
eQ/2OZJiSzX0K+gTuIN6/KxbsFJE/210WojlIxbjbC4pXhs6ulqQiG13IhCVd9qwgLPTeCsNoWUL
6aWCO3d1V2sNQ6Xj7r5efRTy/vzHgCbQ8TB/KA5JRevwGH1G6OFWfJ8AKCmm8j3KhOufxX47bV7X
047aoB4X7816jC9KvIi7b2OikHY1kKSTfdr15G2ahRK7ysTIu15/STzoYvbUilstjZyosUaNLqBQ
SnpDaQxpAV7COR1X4ERTQbPq29en+SslyUkjGoup9py3fS3vudeSzCFQPw8IRDfbl7ROwfkNBX85
1utPjhwy9nI+0bTiZraSaPdxhm6BUPRoUV/qCA6vvCbJS/b2gS/cbpVOd/WiLeOLH6Ia0Iqtk14b
XCCsKqkzrnUsejC8u++XvmwDfilP4bs7wOgYyOs4eo4ZhJ1baaFQ19FuR6MqOmnU9rxAtinadZgH
6bFAthGx7aCnZKVq0LnVSUmzqdpxPgRdCRQhiH1fD0AugoQ4lrX4GpueuqR3fG0Qhhzbf0I/rnDV
aREMQpJ6174Egq6zvlBofp/r44eWW7KjG8vEUroJdaQdoa0zC79ndKH7lmh8Ac+aY2GNPZ0ahLO5
J7WqDj1DScT8mjtOgRrd928Wfg7kMWe+v5EmKkGKsUJWZR6VPT10G9gxmM/aRPqRe71UCRog68Py
aJ77ovASqvale6LrhRjZlXPvzOnXqc8hIUHFWTg4n8+bGdfUqaq3zr3+n+bnDFnFqDq19bvtIhJT
BPDEYNGqW6Jkzii8OYpqSbkGLDov6nP655GCWdrIdPgJp7/zjOJTcfD0QVqPvapyEyDcciQYQLC5
Du+ikRRURGBGVFWnNrCodCa+7WBlykokKYw9EyFPzHwKc34hDYjhI9pwZol3SynF0/9zRhhM17G/
1cSeYhYEOcmxUVTilo2j/hY5YKrDmbUCDqkzxnky8AAD6MOxuzPA6HBftKIbbjqhdd1AP+lYLhQL
ZG8sc1nUT2GdHzd3zCekw2fv3SXAEy54zMotMW4EQyQRRfihYrAMS5cc4jNk8dQpQ5+TMYoRflvI
C2X7RNTwRhmKj0B+myhlp7AhqcEK902x1SU+w62cjm465hFx1esIBnVE6Y852kLRRSPFNH64L3X5
boBtv4fjOeqcIcT7eEmJfctTH2Ejzmm/m5oOQOzFvVWoRjjIb6HXoNNa6pm2b+UhpNFsmVPvgzJZ
Dll2MQytxH/p6uryX6q2WusGTBe2RDacHU5n2s8HeEsp6v9Lh8aTm9er6JXFOVzhnSXeD/rBchfI
T3BaedwGPpqeg/7CPcvvJCvcEGBM29FYZDcesThmII3vBcitPI4EK6EVHQy4kSStePHcjK5lAZXo
V8WtQrrhyo61s3HNDAS4LRtpVte86xwqU2ybO522H3ttXBlTbiuBgUdky3zX16ShRq5pIrh7YJNu
h5IJey7M5KXRAauutqX3TTPu89wLyvklPq/ogZIxsh08xoC/SZ8UtkcorcZOn/GemnflziC8fW6y
VtwYfHNJ+lwpmxZC8oZ9916NewzqktLAwz6H6Obu5yR1hUU440TxIHYULUvQe3JTDG/x2538PUxl
4kU1fbf0ZVgeyFGJgyOO+3WbWu719KiAt7Zh3NkejM0GQ95uqjlUjv8AdVxjJNGHZftvaDWZiyv3
sSio2c14equQ+WS1nooswsxTIcm3jMtu9AHnNYb4y0Y1j56VmATUIXQYDW87Fkvam2nP92dzrPz4
zcYYq4XigdA2GzNL0urIfDBPam96o7icZzYUh/r6AplSVe+szoAO+G9AK7Sp2mTSf/mHzvPBuLO9
Gow3L/wpvRRCXb+NNQKYYZX8KOhilPRD6KVh6Dlphm75CbUhnOOejyhgmpcg8HZVUZ3x8BI5wnkC
t1LA7/uaLjwlqzDTA4mRWxBNNol9dZPONivICevlJrPKYXDe9ZxD11poNpnBKTAOsIwwcnAiQpav
uCBi7Rguwgb54CX6Y2k4gsK87Wmev+L0t8wQhr/1D7hLC4ag0hmPnKOEUnziheS2yG1qGc+13kOf
Ksz9uP3eRrYkxkO9Yb27JKi1afZZ/8vfxm+avh1WpbfVl9UMfmIOk4tJ4YMCIiQwHOGiOXb0IJV+
2YM0GK4fZtTNn8UQia3GYD4yAam/DhVDsiuMSiSqIojPKmkytTVK4jNuJAShFrCow/gcUwd/FsE+
uS/cyUiIq3kxSJTQ/pZRB6i297yU6X7r7rdXEOciZ3tp2DMSkx9LbKvpDahgBuslh/YLxaLo+q6z
9nlRR2YKSll8xPZc59kymPBUiS2v8GIG9WFG6Nxqf3VK+41nFCQuYkachGFPVo6UWTmqkEbh18hm
T0BSPpDhgampdWZiBpO4rP5OzvNuhiG62ofWuCA+OVstoX7xN6BDutSZpfghF8yk4EbOcnAhyTc/
S4VDOurXmGVpmAp4HVEI9xUHeCjTajfANYyviNmGUIcm8iE9CJefJDV/pIWWiKfdkCQPwdfitJIy
XX+rZKTiI1kg9gqPLhguVV8Cx79ZgOEWy6kk+Lp1sq4AWmcSJmJu1VwOLebfJUMyxUZf1R7nFUPm
QIS+qlHaAIN84nSAsK833sTos2+ykZuCRAY/CJDrzf3m980bKvQJkIfeDUZ4vu/L50Z5T+TJXdfx
bs/RaUNt7y7utqMv6i6P4aZBXoNouIrI/ziMlAl8HqViK/ApIqeE09+sgVB54EwnCcK0uqNyRGIG
8HnEV0LQA03yhpC/vd8KVnPF9WxgpvQQfr0Zv1MqeDOJGBY8Ix+LNTNacKMcUaZ0tqVr65Nostzu
AkrwB3nEcJpiCSCyyQNjIYFfqK2gFmZ52EGfnUHdmDcSWk5Bg+sjJDDEqnzrhz+AeMvg83l39TPW
q5xyVt8TTe9A1BEZ2cXBcNUkohqLt03iUyTBKZFnGMcx8Y2cVuRVY0wYo99hEmQsZP2YexFWVoUP
yHWkjGq4HRoRQWiaipWbTVvVpm4PK28T7CBLMr3ha3O+tCAHTUlwEr/1auXo5YFztvSy67osZ8fc
VZVeWwc0EGiaREEY0G4WNFLi6W7nA3sbYXfXlXM+MKYhAEBc0wp43Hl+SmtTmpFHciPLCt0g4+OB
xS4t8ycuIp8ukooZrtR7tgEQf7W7IDmgKvOwUeACGYdT+NHp3QQLNvQxLNdF7V7ZK1/Ek2pxafnC
LL751UEeDSCBAyo5oU8/YYE7gjSKhFkethsOX5gQQsBPnRSRD5sY30q53zXhKvFAQ1Fjz+WNJBDp
fHU7JJq0mPiBwALaJU20EDIVZdXJDl0MtiWUv5Gw06vNrqsxDwBdVIiqQAy/tTbMVWdLdCryIDeh
bEOo7uv0eRnmZCL+Ym18NlbdGMwbgWXWNMbkIlTBXjFFj5rZCalZtIgqB4JMY1jen9ztQPsR6cae
buk6PoQYAS36Hx2Z9Pp5nxQVB+qWGf5GxUnp7ydAgYcbRFd1cvCyMvOgRFBF3Gr6bdVErhw6Wbe1
wQINI5HdWx4N15Ja7U8jx0omGbducdnrOJbQxQKs2zYc8VWpqdsD5ghnLqLo/FRKLX+IVTJ7GJ0g
GLienngKSYio8cvSywdADDm43GWLj7gwQYw6fmw/5wVAZ0z2HPR90KBMtviMVCGH2JjturRyXg3U
xt+V0iUT0m2/ZS+1JG/fZStT8hbU2jAgGSOOqZMe0OEqKmJa1rFfftKDd3fd0yFJX/BUqTWtGiEa
oNPrbO8Pzxt7V3K2wbLpC1uuxUhkMTbGlHNeryqoIKuNzWrVEUugzHRQAQV566dO23PnqcMOhxoF
qm8D6VlRqE/3oLnuDnyMTWowWf8S6rAItS9L5vkQCzn8XATJdX9H7PcAYAd/bzF3X+gTDczeAWZh
V4vTFo/gCEHnoyp8jA5nJzSZBOCvN0Gyvz//WWCal1aJwIDZ2o8pHAnzToiNv4IMc+qNWRwNljCE
7PgNpb3c/3ZGzil8qokl2UW8395dL1NC85xxkcnZDMiIJDiMzkTyvpAlnO2gQBmIqvXmW8zBIswl
gDJi/1R+vhYSRv7MoMcYnD2gjs7gVcGC/5nTPvXQ9q+z4nVtFt8sk2HqsL5C89rpH6WI886vZ/lP
fNKR3FnAAmyoWn/mYsGMyic/o3yX4r74d/X7nrBrljD/kx/alFnjoTjp75O5lrLu49XrZGD+b7xB
iVhbeEy9yPeEWizddVtCrODCmXunwt6mA3qc566W2i0qflG4GepGiOJt1waz2W/FLlAevwXP0OBD
BU04U/XeS8R3dPQPA4TIsbFcJQ4qrFcyGuh3HqACyVaQ16BLrNMGiw30YmRZRl+bdY0LFYRp7wFo
B3tFiglsniu2fQ6HU2V4NWGUyoyGEXlPZHCVxxrKqYyNlBoMfi1hdnpQgwwQkTJnO/AznjsYl8ET
R0yn0NgpMZgzOL3tjuPo6jb2nJv7kjdLKEjVhH9TmUScg8WLnSn4+2Zq6H2aSl2Psw6gX0KHLJ45
K9xS+Ek3YyX+TepcAPgpxDdoUpsGnWVOH3gKLiemVD+ICxh54YrZoN3Qo3dFTCet76JTPRsEVvCC
wr8pzCb+aGbgpAAO3fr1X1LQQ9BcH9oaI0G/8u1fIalLNIRf4kw3mtnKC7G+Suuo1sbCERZ3+0V6
Flt+/AD0vS7I5kqjVJiqpkio65JKgQ/NhOQ58V/z89nOOPDfwpPCGv4+1sy841tot/9/+gHyn1Kv
ZJR51EuPGvDr/S8ADcQ7y3zwyDbvVK8VUDaCZPjdOO1rgeA8VVk7lPkCZGsGNd6JBWmIQleCFcgL
9cTUHMG4dM928SVD2AWyVL+jbuwdbST0om85/q/mapmZ9xW9wM5ZRJRsngRk0130rnO+3pBq1j5r
p3wErQ7Qx06E1KmznzLLrbtADaa5rqk3vfRLKmiTPFObzMPAIOh4mmqWLnzDSPOvzAhqiaAHXj3l
JBdC1ORQ5+wuDOSV05sopwJqIdgtokm1/JjiORX/fR5it4IcyQuT0gsYnBiR4+pQXJkDaU/AcYDN
bo6U8uJITRtx1fNUd5/8odYwP/CJAG9AaGeUX1mQAa3w5CH2zBn8+gSaWU9coQUbjhz13PCgsunF
dO0AGOfzgs36y/h8t20WoJNHJiOwE3myHvfm+nOurpHFHkJ6C0leUjsPw8UlF3EA+T52IAhaue6g
yflme9aB40BXszEQRQxEN31vY6Q64qoyMPlexWsTZLT9KkCjUckQPcVfN4EaqY+VPmAcGnUAIa+k
370KXHfBfsKESFrg/I0TnPUtLnfKH3RMJcUiY8wDQCl5+1P5pbcYJlwwKB7Md4NCDf73gsjpcbog
C9jVPHy+A/nqwFqX7ITVBhpxkImQBeJvMx1NcLel4om5YIAlrVNvKuRGhCTkHPbBCxq1wP90NBX8
PxBOmlJktVqzpYg4HjBF9S/rVeogB76JyLk/aT0VLtDxPDMhsdglvjcMky7GFpdwMNNSSXGE2on3
dEekS5eAqyhxuMMz+EoQunJmsgMaQxt26PJsd/f7+2hb4GM3BDwjXLlpZ9fnzuV6enixQsuMERtQ
NrEZx5du3TjO6t40w2GPOGgsHSxmh42myZe3yu0b7Tpchv68uovPpiHCv8W86o71Aj7HrNS1aur1
tOVne8Bcdg/S09DJafPeDG6ch6lhZUFmd8/nWJOVswVOWN8aJ3sug50PdCH2LNNUQUbNW7txfEI/
BXbH7rqjbhi6yDAqpfGRBTuIeudQXf8DuSL1dyclLA+MYVvpHTM8aHJjgF9cncQiicL4S99DI6EJ
SqIFdRb2lx8wXgSx7rKLPpSnRHKATOYTNgA5QUwq8cfnwFo9rwsvFmNtADRLbUK4DpxQqg5A7rGb
REGwVsSyXis5p6UD9c4mzgkRU/9C19weO3yyBy0oCAY537ihkTY8VyQWvE49+3Tj9pfY+zNadnzR
Z6ybnzaXjAPDB4ojlMa8LW4dh/69qyRdfgLbNKS1aWFZmp8ruOBeRmeHaXGZ/k/FEsmT+MHCebKm
6108hc58bLqDq+AoiIDI5nic19RgYHoNjZZpLx8BI6anCSNlmWghhS5SuV/ak5d+ccH6XDXZybFJ
o74X3qQ+sTquKoLx2OXFkPbXFmiLKLqPxqEu8AqNPsmKR5VlY5oMQVsPt/ZX4/5kLaU7lyX5UEOi
o6Ic+t4dav285ChJOo/HO6RRUo8PANdEgeOPrB7QjpJ3cMv2lVb+X6a/d1MfBJfUYJ43sJ1yOwbq
2ElAtgl8dQcj0wwdGZ+Qf8jB+0W/9QGLj59ANfKzPHFyyxw/yyRHZTxWukfDpRpDVgoPAwhHLpyr
1MT2tNVp6oDRLuBkYSD6GpiZsofmmEZD1EJ8oB9Doa3pr5/B/mT2TYB+kB8Cf2KpnOsoJ8p5nlrQ
YgKbgR19K9Czotss38ONlJMhdh9URlyyGsURdmGQAMlLxmdH1LdEZ2a/V3Wno9dPHUHgn6/W7Rj5
SBE5iAwllgUd713LK2PXNUAsz9l8yOF7igqz14hcBDS9743ZrDIB9TIuC8qLlUZZToCY22UguE00
8zkdkA88moVRg39xx4+bT+7hHHmzb/4Hn9BYjLPqyAQAlIGO9oBatAzFsRVp4Vfr9uOrCTSZDj72
eTWa/nnDcBauvJbD2m9p95odklkEsQWg8yHctcap8iIyZfsebwfa22N8ATK8mydX+fy5zUQliVpV
m4jOd3PSmnkKci7qc9o5zHAJwUPD5VAJhfY2R11uicHZy6U9gISZ77BTr7xAxRWydVz38lsoj2FW
AxkLCdSjyFw1g9g/jcahiky2D1ELAb7f4he3Jo6mgaY7dzifXjSwqh2jTK+HgjXiG0QrqxfQhQ5/
nGk5bGr5g5KO/631ZhaRhzIdhAU8K23ic2nDObSkNgCemyM2T/HCu5NWF6u1ZMOAmEbxO2aEPsiR
QxHoIHUOpQkwYtxNcj6TL+8s9Ym7GsPe8ZXywwllXJ9DdPajJnLJ1hiJ8urKGDvsz/eLQzUSSIg8
mhvh6XDYdNuDA7l8dchsrQhdmTzkmeOQHICY6zPlVe0xH5Juh05iXx28Q4HvtnvBjw6dRF60IfPW
4HsyPlT6C6ZDtcNgR4BPYq38W4ZEyqyozQxN7BhxxcI1YqMoXJAC+7CCR5ovKRvRUbr+iIaGOw7X
kRcgYgpfHb+BVTbU49bp0S6FLIge7uhSbgP8gyQ1GHyejS44yU58sWQhwwkdXom6CyarZtzuRKvn
gHhtbHWfANteXo3MnePYm8+K98VVrIMfhO9D9B0xWoVtPiXkHlJ04xAo+utmYLbsOWrnk6UwY0PW
wrQpdAbKH8DbHVSNJaMR9DwNRkFHu+QlwGjeCVSfQV5qJhAWrlSffjAYIxJgjtj9t0GjTtaGugwY
Tet+16fIzWXThCWE6gzqM2eHmOXLb5J6aB8+KIm+H7t9OAmkP6ffURG5D4KCsUJV544CPhASieZt
omnP3eatw4Beh42e2Xut5Uo2T0jald2K1OXA4dUnnlY+BTSbeE8a6Ghz92WXHpGoL6Olvaxaez0e
wk1bs0YoBsKaX5PU54uT9LeDmzp7hvWzEB7XXbVjRzZorLvACsncZTobx326Wi+Cd4WYr4GDv35B
QSjX6R4lpvvza01HuPfrKvJNf4V/NMxl6/1v824Mca2B/5mt4QuJwi22ruf9G4of5vtMZtzFITI7
NGtnMmQaeeUNEPDNPA7gqczez+UDd5TjbrJqeZsFkqTFayrLwInczi3ZdMY/wE70bvFJQeJmp9Yg
PyOeJlEM/ZFzsUme5K5wtDBZJ1vbodzTFfAi4DkI/KbYaiCPUuAVSJMazY96IA9koBDCooRiqmAF
TTjYh+0cSgkfwzUxfel6YWQ8Oc2bVIAnbbJvkUNuHAcj+5UvlvdXqfv99Nb32GD1afi9n9gQYtGE
pRu4H5yteaXjw5uhXoYLBQHSbR08CC0CLD9B5Oon3yoUdpguFbf4jA60w9eMgkuIKzymbxaGudw8
7Mo0AUZSlD7EkoXaIp2pU0i0HpLPoV2oB7J/Ao7U/O/qNBgo1QslBcg6smZkvUA6sCR7+15TLs+c
QOpjJLLKqGPj+qxuELq2iggMqsY1yvwWnkFJ24UreVSLkoLkoxaqjHBTCI/wReTF88u9BORp5Im8
8l6rdbX3DpvdtX4wI08eeUq74h1L7fIdjTdwfpBQrJE2RqUg3sHxvN1d3KzycRP/EFop0RpdFt8f
h6vRaoWarU2R4R2qn48Me8lNdAxtL5MdvMGy79hkRL8ralbjS55aC0mAr5Y37TtzSKKc8hpi5q3Y
xWFdLxTgFlWGO+UQLU3cfonvN2EHcLlHWoxLk7+BiTu6k6T2FUgdZXxoqg9yTXa7gaUsW0F1iV9E
MQjtMPgWMIl2yRyYMKBrcT1msMq4O5Y4zJK6405POhdR3YeWAaYJIaOzxdzfcQbTrRYYMKPiN71+
SiVitg9FxWh9l+LR4T0/lfFku7ED5jERa+H84V65FRNHOj7B5LNkD8F0r6mFQCyRZWdod/kXKvlp
+/++IcQ8ZhZR4t6ryvhXEcLqro9u3LU4l3Gdk18n2ye88lIInuPFDZt9ITMGYuAIFESdxJSUt7sI
7htf+0yyX1Dq073aTJNNrfnenUqzKSkYAhQFknbPhEkU8QaGHLyAQG7hmfyjFIUpvOZI4WffRAmO
/+E8P62G8+61mZ+qgsBXqaHgTzbLTG8mjwOpKaVnfkBbY8Q5JT9JnnRfkQcPV/QUWeFUDW0OaVoc
RfnB6inR57gXg0vxjfOO42SBqF+4kI18Vkcr/TerlSYigvj28smCcz5NadThBElE6rc/Yw6iG64e
8oLe5uZV55pdJfT79SAdTqUZM53+lUGaRHyro/pYzijuvsXVVHdycVJ59wez22Sa7Biv7cHUAmdq
qsu6f7uaDXyDiVsw3Z1HSracNwdK74T1Yi5j8qm0RGDXyHpL8moHpleCFmyYVqfWG3u0nvaXVyAS
YcVlTQmIclTBY0nLXbbBQzvnccm5DUFif1Ku8p+gmxv8o6q2+YMxgkShh5cqEuI1aZLQis8/rWCt
0oFh8KNjmW16vUPmzuBgIsRdfxJxFO5e8qEJL+1DgsK8fnh5zlHjQKVEB0VbTuHvP1/VHW6qUKfP
Tdf6XtuJS8Fp0kjkNGnQtZKnGVWEq/MLkAhO8BTsnZw0AZXtz8KRWbRWzc+vXTBQfZm5GafuBnBj
bmRIvolJdyJS5s4Q2wxDb2nI7aqEfFOO1NaGyfvaftmLkp2jWgokgC3ADgscAcypMpGYj3h0+HZ8
cy+xV0wUJd87BieCOJyj4ADsJBwSXYC51Furg19gxYos2xqF8HI43v3t0MJ+QjJEYIuFZ60y82E1
2pLzO9mYL0sZ9YA3BY07C1EyzvcAlu5UFTVFpJd9HolNpYHpHL1ZUF46pFqBpJRcDOAM7j8gVMOJ
JbgkWc1Tb2Vmrp9juv4DcZuj1diRlvSRow0NyTq28vvLoDEHxr36Lbyoc8bJv6D8y0a4u/FpqTFQ
IsV7Y41uP3N2iGFlO/4SCmWTg1F2HDZi3dDFo6MOLMIZEOD+81W4YvZwGyUGmtyeLgAVhVeuyzyN
AL8yF/WmitLNDphPFESB/rtYHTVNm0x8OrQQL/NurONTmW478I2BckG+9deAFpt6d+W+JcOZ70IV
1HUqBpmAgvyrHmmR5SbGBhkgWIiKiP7SH/kX2f76ojDRBi88Ec2kP8WBjysGhY86aI++cxjJ5Lyj
AvKGHCDqLQgTnVjmOzyZkU76SRFftXxe5cJS6mC2p1sgs3IJQ6+cvdgw7nltyDnHSL+WBCTxugU6
Uw2dXbi0MIJpZQXSBusyzmxJn4CH+nQCW+HwNPVlJe62akYZA6EiallCAheXc+90vMDFUOscigwR
dyYbtU8hQ87RveFNSJqRTmejDRN6ByOjXWk835AdtoF87iEiiEwdgsTDRrSSyglULPpCiZgPSb3X
ENp2sq8dbwqNbZs7Trb3wbRvfVgjyBDq8SU2fNeTFhWQKIH0xAM+UZfEV4jksMceLs4OcXfpu27Y
Nk2IUpPxdi9imbNsU2a8nq0OGxcAifsm8ZXc5aTYNO6abMl7uidD/B8xF6qcmxUkLpXbEIpZxMY1
5+yAMggKhszkndgifWjx+P8u9a2FtyE6Fj7uxRFiVxFqJqCd+9tHNJCNdQXq5ZHgaPMwtr3Fm5Z5
LTnkDnH4cK9kfsOou3eP+cWYsow2Pily23pLwIL8d7D3aGm/j2Qnjbab0sgJkTt+S5H3CB/5U2Vo
o1g1EromNbfYczu7pyfKyzYgHaB870EOajc0jdHz1LEsqjP9ghkON4jcxPmfIJDhuU6iCODlDF9p
a+DEN6oiuVlM3mGsdB0aTc6M+WTMKBMehJOviEEYqIslo32qTX4nTOGo18U+shD52wn4LWS5eZao
GUpVvTHfncL7/dAZKL7kqH4KX5LXpANxQheO1wV/kgaSp7TbZRuQADgHiqIuBrE/wKLJXpGDQnVi
+l6rm6Ipb7kmI1gAU9i5p6bt04UaUBAli1aMr7xpHBwskShOujKbBZmFjIMwDXpWId7BC1KzPLwm
tziDwHIW9+XWWUDT8xqSWFbVBL1/pExq2c+fHaoj9SWetGxm0CoG574VfvdK8XyclTS80Fvtz0Zb
jHAJLKs2Hhw04vBYY3vruj/yfTGKzMBB435xIi9rZc+WPPrxQBExyKITLxGbVxSuM0PPzj8H3dVV
Z8GXShRqISujI/FAuGOIoas/tTHHWW7QFrgG2+gx72FK1cRVyXeOH1c0buuJh8s+Gddfcq3Qmta+
OP/xsSMD/vguKFCD6u08zz1djmvE47urX73lisRr2eQCP/e8Cy3gpQWX0rYqDF7nXTgUtPuCvdOo
m3v8tBbzz05L6fq82nSzWVRJAHiNgE8P27R72INX8OqJjTAI+byOQzet/M3V22ysYZs0anVn8cdu
+T1iuGahuj7mY8B23appK5jQL6JQOq4CGWULZQvcd3XnKVQwilnQfbO3NLHL0DS+k5iGQyhefvim
0t2naKUvPrXTL91dyBgc5QilX5niLmtWizOfZesof4QdEWfL50Pb7Jy+MhmZ+YNTgeJZmObmAuPX
Q7ZYlrZ2vCneB2UhLA+F8+1vHt2ed4T0YaHRh1ONVszIoIBQk76bNjTF/ZNlTHeMeZiz4kSqCCbj
b3svLfGP4kH+Pnls1knl7jAJwC95bZGsdyv43JrmDiDXiX6a+saPWEKHIghAngZItnPTlRH93RST
FnrfPZMv1DqPSrvBXlGBU+g+oFr7FW1pSe9N+qFlLD9sKfHvDQW2EENbtUajsjgMoe3mPHiID0QL
xHXKOAamU1jHxfUOaAEXL3qDSu42sYR3ZK65A1sro8fuuDUFSxFUIVS09X7GeOjYiUhtiQVUX9/L
ckk3oeBU9DX88cynBp5pEIycmDTSNKBCcBjFn3YHHOQdk/6ney4t24C3PTMDrenSr78CbNKj+tbv
Tg/GVV7adSYuNlIFOcfyn3Mt6soxjn2C8GsDg2KoHR5Mpi5pA8Y/i/vHVwQsrFianiRNnsvyiYLM
3DkJ3mEkPL52IAZH82OIz3x1homRjmgtDdc1HZnKj7vfE6idoD0fVQGxD4xIARy6pSmtkm/hA9oE
UECTRtXkTdxcf4L9qxzFiEotJbaMPqF/mEMQWW7be++bnUbJBmIvjFHftu7iir5abLPB70tITMVX
Te/n33WBYYRe5dyuVBvogyXVsYoRoFjrzcoXd1v7emvPYsR1qf/eThS4dRKVJr51PHXHmjfJcz72
OW6vY6dwfTxEPrFtlWCFqk2hMNvP8bBBnjstbGmSg+nMIPgBc/TgwsZ8Nb2Jo4mDwMvfZ54gfeQb
FFwRKwC8Lovp/IVJCG10J/SD0iKkMwvkFviDHlJv0UKMPgOzbEDOAU43SnF21CwnUmSlVBlQWf2m
vPgOQJhBJm7/6N52FpuJJf2d2fmXazCB2Z92+wHg0+DZ3JAVkUPr59PTPTmXyFhj59XUGTSt/Ivl
iKgb2qlBRyhnrcQzeJFC9jsHHL4aSBgmz6E+SaP5SR4KqLStIn+1HEqHZ2+sBS40pi5cBAYFpLc6
6p+KX9MRZJBArSA4MmB2zY2n6jcxoknmP22Re0aeqkDDqJkvnepVynTSu5qQIWOksIe42l9GhBJX
6RpmMJ7uwEjDQsB+G02/rfg5ZRNo9u+Q3amaV2VAynPEgkKvKlOBu63Sn1eud97yIblJ0yizB9h6
zZvdEKKwcoBsqZeYJRFrGpoRlqqDTNPIKA4EU7zAQF9VDb1z2HmvJpKQtn0Nk90TOHbmY3K7sVmi
+DCPYmGCUYXVp+lY+B8S9z2mGjll+jxjyK4/izg9zdrf1JgcKbrmBshOOIZNmloQC3LXuF3OEdn2
546apI5NEN3iIFJghvgiswSr7bUvivKdkinlRrgaPQW6Turm9pErfbd8/Nn/q6kOv26/bEaXSzRZ
3bwYHWU+4p3+unQ2VXBekcRRPTxVVTY+5+DNqnjYoOPwLz6D9gDY15jKZrNWDCY2oUfen9I47EF+
KtLnag5Vc5ePaRtWbSwX+py0hziq3J9YR96wrP54mItESKgt6v1oR4h5KcGiov2qJKZIFE6NUGHi
SZKHN2T0sfeOzQH8rJv4YtR+qaqdSNScWsrdzZHSRWrFGBZX2Hg6QYosKi7rkgk2GR6NZRr10OP5
SLh9GAPyt5LB5NuEtZIp4jsIcLK0yKPDF9GeM8R7Y8gRy7Km6ILNT/eFc1h29Y6pRuXjuMGqzBPX
BmdFExQPqPuyNUcEnK5B8peGuItwRyQD0KVzbEac0r6oRJeLTWPJM2cIlVrZntOXHxo9thpBWHEh
g3Oui5Se5BCOQ7J17CTHLgbLjeblfSwQNh2uLVwTyci2cZvxFP3EiHDYBAoUN2zTtz0iwj0a5fBj
gKr2P20WxfDI4uzw+uSza0kifYupZfAtOxCRSu8l6/NO60BNJo0444fm+cvl+LY2PWTEJMf/7wXb
rVvywGWApcCCYc9xFa+Zcq5AI9WUQ/5/ksO6KnivDaj277+ARi/yJmdYTkKuHaEMIRtXIUQO/e7r
C2F/XGB7kQ2eELfcvAnq96AH3pCmuMR51N6JrNLhq/rQRRtrUI+Ev2yYlL77RUsz/gDRmJePEe0c
iy8HvPXxxRjcGzBppHF+pAwJ+lUv5dI47cvPwMiGitUpTCtob7wMW6A67GuLTe1VY917ZjwV/L5k
GQmHeOolBjZ07ImnnmVDmNRWouaR3WvuFgtM5+ULBvcDx544nNSX5g6IQswnhTEYiLewubBakJC2
ddh6O7bdUujZLzhbLQGMhr7UB+/LwZTu+MmeFcqoi8WyTrMCFAFewi+lnD9dEh82ikdhfGIUvFrH
PC93TeoA37mcqFib7tUZU+NYNKH7dS4aRIs5WQJH/bFN5aCnRqgZsg5JmJVg4yKWzTjxO5iJNs2i
r/Lbn85lk4n/W6CiMCucAUYQooXbqurkNr0k7VmKpGj3J3DN+AbYFwL2rUAogHJbrWMckSEuOFhE
RcSDE+GtuZXMyHOBGwRGPWc8J2NVOz2mFt0b92t+6Z2Vlfcu8qNDJxq15uSHERIcHNrcpuMTkC58
UxkJaw/oJWr4LE/91VJFZHD4daKOAL9j1XWcFd/yrpwFhG6SrbRpGhSyqt+Q8qqAOEOhsGa152bB
ystTRiXropxUlV1584bozfTd4EE8rYR1gkwgLkpABrEsjnh+HlyUAeA+padimv6V8jDw355zpsV0
LG3bhnyvvc2Ukraj3WoupXgLetFpIhYFjdzWeDQy/KhN2PwiXdhv1jtMFj4vJTzG+XmSfsXS85q9
qpW6toubThvo494mLzt3SmGdj7OlBr9v5/EyyEjERO753SK8K4LXB0New7pN3dtp7fFqQUEwnmhd
AwZz8KevcY6Tld6HBPPuphxXVLZmumL2ciibU+TR3CDGqNYzqZ1gcm7QvSFUK/cpKc3NwdPZHi3D
QNk0ZytcSUEfUqfE+K/HfGPiG0JmyNz0qRIwSzAOC12AmflWdTm5IEhc534KtYiLhf9+0woKi+vL
nUsVraVZpWtuj7Lbgobk1FHDG75aDx5lbuzmHM5JgsGgm5BwXO4R11GiMHW+BVJ6bm7uDeZRIW9x
BSJir8gNZIeDFkrW9YJ5KZUvuRG4nPv5JtXSQ2C7BPg9Dswlllll8NAaXa2CyQyt4zPjNnnlh+2G
ms87jj/PGcwZHEsIWGXn6HISa6JkKieykJkQa23RXZ6Z0FIi/iB3vGRCJ3pUsWdpRFbtPmr0rMeO
IT8yelwBJZTLHyvhoTjlZO3yuy8ddET8NYxJ4iQ1G0qDJPUxtw5qXHaeI6xk4ySLA/SD/ihD6oT+
SXaElUXi2YJKqVW8Xk4+ND6htkTu35/6+HITfmuDO16Cv52wfj23AN5O0yd6IUCNU6dfUcOLPpSy
k4JtRnsEBdqGbA4C3fyHH9BK01FOx1z4LNwvU7erDCoaeW0Z0triTZGdT1oR7tb+Adc14MvBKVEr
yf83dqh2HdvTA8t9Q8dYPlc7LCPvFhBus23hsuUBOcOPtsfyC/YRAe+fT3OefqMjKb0SOyaN+R25
LFkN16kT0m/55O3ixJZ8J66WIntKunrr55y0hAZhcITzghnEKAMi+zua9I3N3ZqdmeY8GdHcVdtc
lDkk3Qzc6OvNaoBUCYx4+SNJmAFs402izi3JLS+Rhf/ql5hnLMQIcrgXvCx20Z2qfZLz8YWkiwTF
vBBvW7zQMpKbpqSRVYoklpWERMhAa8m7e4M/tDIQC61k7Nu+UC+l97UCYYtkYRjDEl1/UYH1P8CE
D0Q75TpXxXq1HzQfW/1yvsNNfqEoGfBIy6L6r4ssSUmZUDEk7p43O7syb13dGFHIN4tN0VAGCq7u
H9Qpif1n7+5RPCWCXaT1+o4djlO9VMUPXMZtx9BpYx30QDACKIvXaiGTV9+K7fQZ9nZdu7kHeSXn
1rwY5SU8QBGdjAIiHOriB2zapx9W5QUyMSa6opycVloysoC0KCK57Nk6aCq3gCk8F16SbOqznjVH
E6StUCG6oc+lsYq3qWFWGV/WtIXGc6PiMIUVVl0Ob6vg9gUwH/iy20Mqbq/6X6slv0lWO4X5P3tv
K75Mpz1Dsye5SQNnGg+1Y1hC2RevxIGpshEVdo5JeVhL5IpLkrHCK8kFgqWrbVMEypkICyLpORg3
L7MY2u2Zxov1GIJETK+7c5kRVoUPOysxCEqw8aJ9DRtwvXHklHetdmGJn3d/0GzYdlsoYreZpghH
BZr0Q+gjzljaZNQppBipB4Te8APHhLZxjMZNG0zs+p6Wp3lT8wILsbe1/xMCN2bbBjPBPnazP+f6
Oyt327wWoLz4nLpIAHjXhq+s5GFSxTEL4+V3QsKDO3ZxkFkVaUBzGQVoZVLwGrxTOpeAnegmJq79
NhmTcfUCudcajSvvveKrrkZ1JDu+Gx1rA9EELNTXtaXWgjHtqaSaUCmZoqLmUL9oLhDmIIH+A6ks
2+6o8NViY+OV/FFYzsaDA5B/AScBm945Yffv9CUnKRPqjNLQyJfOcoZXxpQYWXf7Z0usFwPPtp/o
iJ+p47NvfOTtXkfqUg4RbSzyZv4PPSnQYX0eG0Wt2+yrexj0awZ3el1zY6JC7b9Yzk6NRMBAjpTN
VjwEfYso41yM7iOWx76UN+CKwYketIoMu94pnhAMNzG0hzQ+L/XSLxkbibWzEoSaCmrc73p6PpxC
Nv8SG9OPnWj5XoUB9qPeEoXKEl/y6DstxholZVNYWy1MzJdZq22L+2Yv59CKTPTe7cagioEJlvh0
8ObX0Qy9HyZBjZ/dFDneVK/AMvJMm/KBnDk7f2vOOEvi50GR4DwKahQs6tbWfKGD2Z3DKZqwqGR/
ug3vVu1rWPQQZGfpquTHpCPy8CQFvXYCWZDq4uV6kzA0Qg6clQh3otapOMn0cmWkFJpF45ilaQfD
esxL1L0O/EG6iFVah1GYPEI+UYgb6NXTdh62G8hnN63nbFH2uIZ/6Xc2GonGoqJwLeu5YsSnjMF6
gssYg+WlwG3hzH7yTHmGfCAhFcQtnlqaq3Kw1ef5qNy1wvO5ocBSsYiKutnJLd6KjlZy6Ih9O8hC
Shm29/AuNrE02EPxKYS6P7rqxcH/pGqUVvvsa7GmCCn+2WXZkHv7ye9Qh5OT6pfVsE7avg7jheV6
nZLF3GkB46KhlnxWEw1gpZ6zmU8RyYsXAiM3ejL6JMa+8WwsZKYSG+HKtOBxfr5v0sQ3umMlf6Hr
sAVPs6fCMVFrmMY58YXucww2kmnOxMFxLnJQyluQbFNxLBgU9TVnp13AkH4+eLE4UlycioqqBAui
XUZqSI+387UYtXHeyc1twwKVm+bzbrB869qoD4ZpL4Yc9jwT26J1PUrERvdmr6DC2MJttgHQyMyA
SYn3PRicJX4vaRYpXTdTTPS3cxl7syBU3r4bgLELnqUBi77pTODqekgWJ9Ke014m1zmjXwHg0i1t
72gnZSG/S41fjSenZ7UuDFPEzmH0qSc1a84d+DWZE3x61QDT/BU7X8qr+kiwaeOpHWi7WuarRKZD
T5bZKzSPdbcD7IZaOGybgIQ14MWzHEarhef7ZbLckWLz5RYlZOM9RGBYHmHPThiV/vB3vT9yP5Oj
jEc343/BYsb42l5Tch5IyhZ8g9Ed/Cp0H1PKPcqQKmmw88OR1H6Mvsh8A4ymfCorBhk8tgEmYzsR
v2a87bAcOcg6hHt3bcGi6H3RIk0Qr6/5rQZiAgBIiFHEKFPJmanobBH7bGKnlFQ89stlQ7ABnaoi
MGE5Hj+bX3VzzcoMVPE21wL445UWcS9NKSNgtpY9KH8G9won4BDCQ7O5//ICdjpW1XDqf6VDINjv
MW87v0fzjxdw/xKRBTo/4FCtMKQesEwa1QVuyzzexoD9NReuThWAeCveVzfxEaPO2al/oot8Mqcg
w7S3ERdVnHAp0Rm26jQSvuOyWWCLl22c9/SgR4uzyufQZe02BZ1U+hGeteyiDOFnEbmjI9VDRNG4
IGB0L/yRQ+aBL1JdHlAvWzHeY9Vwj0sf6NMA7PQ/qamCz3JuiuTv54SIZncHynVq4LhEINQySywS
xmUNe0Rpr0Hd312YztJg4LURzaDIea/2IIN1UOtZMkYoaS2YuZ9IopzCyZaQsHjnR2/ax+UNJQBV
UQQw0rZ7WZwcUpjTmjRmGHrhCkAXzX2E5rHDd4vpJgYdEEs2fqjq2Glun5ckuwFIWuz/9qPD8PuP
lkLRMbHIQvKzxBLcpUWPBisHF+Q1+RUAHkER2DNPxQE4A+myo/8zrmB9OQbmtOzPL4LJ8Y+IoIiy
RbFHodr1r2uwP+dclDv3tLpNUuApDSiz+Jd0S9vgnHlYghYKkspcHgo4TpEPYvBV9xG3wC7LQF4b
8oScJac898d4/CBYjfbVwFZDBGL0bXw59VjSfdjY19AggIdDFsJ/ZPuyfcAZlcykua7zkFjvDNET
XoTCBzfyXOBOdv4KAAjsXOlCH8nXBxWXNz4jM067brHE1mLsxjaH6dhLNtrJCGjG0IQScTGitD0B
7OyNw6UwsevIkFpI11HuORBKkElwqxTZ4pv7XNae3V9IY8DyYR823K6d2FvyfRb5h+szPNybXqUp
kzgI+rpPxqhW7sXfn87QxeaFQQDAXqcTitGYNorBQoZ68WdBOo/0uN/SsHXAVsg4zJ78ve/uKERs
vuI0Lfcsh57F6tUi0ZMW3+SC3WgMeDcq1X1XQ20OFN8P+QpW71FYV2kKhX9u2CiCoTqMZJ1w7rLu
nkc1QquISTrWhKc5fdUPjb0+SVZQstnYXU861A8hgPsIvcZ5+WufRgYdPRNfTeclDhvm4+WW2tHr
9TM368c2XOxDl+xD0ySQhZV1DYjtUVGN1BY0LWJ5ONxSDELCHkIgPVxV+iQiQi4R4Yye3sRaPIsv
gfR4jtP60/3LHOj3mAAvz0Nx/XU9cEVbbduSVExtzcUy6DYHWdJvWK2rG2ejAxXNuemUb7lggXtq
8CiTkg3JsFH+t8Zibr5m+FUaoK7rf7U22d5cYjw3wED7mQhKmpoxDNAKIFFLXGGZhDfvs4XOhdgi
+wdXqJ6+D4TgYR+EKFIuVhp3lCUes9Sp1ekP2o0BP3j0mb04Jyuh7Ui+f3aMhfBRoCSWury5Hre+
vuUtc+PHfcs2WUt8e2QhP5tafrzhUt5Q2W61Zf7xsAn4TjmHhK1Eh1pYID8BJWdBZaa3f7YmzsTP
kMp/szit0WFYVUbj7nfTXact2YGjLWYpKGNjqI94wqPONbZw37bUPyGZ/AS1S91GwuurX2n6NsYO
XQkcHqYJiL0ct3i6fErDrTcuTpu/0CqV9fGlAcglnocWXQq8oByW73eBVMT2pRNTyGK+DCYe4g13
CMRFWrOjsPiWrsBGPKN7UfC1HidrhB65EVL1jyyE+BnxYr+DyeKzahfk90Szmjoh3B3tq+00G6en
C3hPB3DDGxYOYPLos1CaZy7aMGUObrwJW60g+D5rIuLnsoIbExKwTgjqC4wzQP4JDL1iH7sCRhq1
mclU2xZChKKgG4+IId52p8QsrNyzm83sQt5N3jJ2UL7MCNWqCw/6Dv4QfglHE/i6FTiRKKkjnc6k
yZmYEIq6WJrNyNp32fjTzGOZK83BREF6BBr/t4L/3ncDSfbL3wUDBdqTThzOM7g9u65rXUjqWzfb
fGO1sXtevDzaCQgcqRs+b0NrwYYuGL6577aUngYqe5McdxpwsT8gKEU0mUK9ei4WjHTkdWkN1dYu
QV8HSxW4ZXDcP6GmCnG18QhSvsz7oUzDye4obCFiwwyiRTeihfZHsFfCVfwxkzq2hKxsbVNutXf+
S0zyGSZPULQEwNLWI/79sxQMmhR4zaMMjQlNyshUx8cqDGJqWFlfq5Cj3zZvI8vG5j62+2eJl4JW
N/GMEFyuu81+C6VNWLKZbZxXLuDT5FPQH+ZoBp0PVteXl9dhbCfhGMvyP1H4wVlA+84evX7IBV+s
jwS6YfJbY3h0QBsolfSrhP9X6Tpih4uKcWckhD4Bq87g+rSRYFn6o9K4axfRvQz0GLZ0EK/SCQcy
NXNVZyZNmKqIEtJKajt4nwgCIdZsWKuzyaDjGLFBGMGVP2UpHpIqMpPPcnZMmiA5HCjUf9IIgnpZ
UAtGwvOukGlG55pMmmgO/gQFxaa4oFTp+xbdDYyQyonI90x2qrnWQ/TejYjskczQkn96Wtg/aSXJ
LG1bCgUianPwLfDrmtMKy/PvwHalm7VAok2/Dcfq4pG0Z4OnICehxOpMrl6ne4ggnnqW4w/Qa3Z7
nLUmpECZvxRco2l5bhqpPri5gWfotMSyFX+JxFW0/sauAI0fgUzeKU5tlHNRsVHUsRkaE1/sSeK7
lQ4OMsroceaGx//oT382+RbgVDei2p20WAicLPpI0eHlUlSJ2AYbzdpw4L+wk/N8bPfDAztomzSH
9ZOqG8dcSSPpxYFBUv9ZEAQi7NYAu7Ru3Oi6zUZ8YtuUlGsjs6+oeHk4QlrkYvvzpcbkofatVsHT
XYdzaeMRN5LBasBAag3A/88BFJ2/u9LxISYokLwMw50SesZhoM2PGNS3xgmhftJMVweBj1jI8UXw
22otRVI2En2rYfzDaOVsI09dA87EciJFXZJMLktLoWgr+jqbCPUa/nw5xbJzQb9aI5WMCjve9DMK
o3YyVtfPBPgodQ8+g1FHF2vBDoeJ/+v663nP40oRK+Ols0WYv3ApR4Twlr/sm/c+teJzKFL/D3TC
zFuUWZwtBRXXxEBL7FbgtIto/t4QkfGzjdGZQ2TBWcRACXF5CrLZWGBt/oYzd3FerTIxVMA3v3gT
mpXu52ZEGNY9vD/G0QS8AE7bj8Ci5wcdfTFTarS952uCfrreUpVrDGECXy4GN4PN1bfz69+Z8KcD
z8/wKVnJBEpOHNSlks7VWKkMW2Ca+YCnxKTWtjfWKvVgg6A32JMCKhacZhfbHhj/lTXwQySfsoRl
RosWCxUGoi8/zibPeWv37+17DLDsYvKQ04y2zFq4LCJBPjLs63KLUBI5Pdi+bz4y1Bt5qoOIKncM
8VYXGOilBpeYXi/omLZtiD8m46COLLkJW/CauTNd6sxqbtYJv713Y/RwBtDD/UEtkeF8LwDY4mtV
PyrlsZMbxtfExn+IaiXYfBtRwpIp6FYIGi7LiwRVl7FqgaAtVJS+D6hMX208/RlmnFViCNqHEKiG
lb04iHbHwCBkxothn90fF/kfqFexQEyRPhTx9MaI3z4FN6YqNlBiC7yKlRmC+G8N9Ut0FemInkbx
ySK7XNlgGNI8NjedojZMmx0se9V0Fa14xLl23QAy4iexu8vy/025IDwpRW5srrkDuHwFm2Jhi/gA
3pbjsv2phN4x0dfAdKq/ZQXvTKDdCKd6RiNcU6jB6oEY5BC75zAwyla2FsnKFltRyyjip0+PvK73
rVU0ELCC08M8Yy2/CqLPHB1rIeVNv+mXXVFURmTmkF4aqqYg42G/49YAUUh0r0kTvoAlJ9YwWTqA
dBburuSKTLWGnfpnJb/2YenHpH4PCAIPscJAIRJSV/HCSbmNUCtNCSOs+Jo7OJmitPi5i+zsj89B
9RNowJcip9z9ih4Q1dU/l1rVE9k0Al+4tDj7kwbQGrx5Z5ZfC19/nNqixJ4JqfVLcrGcOfVjxo+i
k84xkR8ABTvObBgshrq3ZTVJ8h7xLtzXTKlwO5qi337doR5xxCDtOTQQizRE6j6xxVHVDzghc7gP
A7pZJOVvqBr9HYy0C1z5JsmGFNyPWhBujFmiF7vm0R/sUaZEo8rEEKk2B6Vsx+CDiOVL0C24zXLa
AF4euunOD0THT8tib8rBUdQc+XQiV3kP8Mnf5AESzIc2xzDCrmWx5K7momSChzBQZmiRm+uStFPN
chRPCSrApluXcek45udHRc3LmVqZWDP0HdZn29TBPLpZr1J8avrUb4msKZgGkOEJi8MTMU85YYbD
ALgmeLxHXGIi+gUYByra1DcE8cFznhGDp26ZQpMPvRfTqpVyCzUiWGst8ixDWhrbD7woo0pydzgK
zS6rjXkULs8FkQv1P5/YssXjUdWudA4zI4xGQ4TSHe1n24TQMWY1pkn4DrWS4gFDLbswuc0+U6y+
iHjjKLDdLD+1ewaeyPbvQi8M1mY9xDy1Ps6DYKk782zuHO0NBQ/thE3wQiJ4OEKt45vX259WjHlq
6jwzqg/qcLHqvboBaDEezDi4/g5icBqqNkw6MgjANkzwXm/M2DNGsFERDjOOlCWIMTi1zHoVeNbB
u18MquGhCtZcd0MeecUToxrSa/fr/I2YJpbrMrbB2E1S8L96HCjVGB2IuYvN5i1THIW8hzGcVJwr
oIHgcuNDVqdk51sICm9s9z+QBxWNlNn75wElQBaFhXJWHemoKtRhcnr+CnmmHYlMN3jTTtRq45qx
fz+twJtVlv/D1KZeiKcONkNk6lXBhd/dSDB8L3Tb7V9mcnVVK06uLxqxgRrWRwfazND6D7uWc9r7
Gts827O8FCqY5AsX2gmF/X3mA1NHAMczUYONaQXLlcRtMgy4XueK+d+kbl7ihDzH/HlIANleyUkq
BKNoR4dczxR196ddVT1XnBH7IiVoItlBmGJurx7j2e6UdK8NT52LEr2xkyKz9mZC4Zy6mu10TK+C
jT21xK1qx0OZzhhjqhJvLz1PT6cr8cBiJEcIEO9xaeV3Rffvmjc/vZshBrzUsIwi614JQbZ4yo7g
1lVRmUNrhBo+jtaFO5sVzjm9DBdoCpftwDgH3wW9NG3H3WD5tJTwErB4YvRE2dN7WvyPMViKDo+6
0AQ1wgJyusWZi1n55tEVfhm94RsbKn/9NyxMI4v6bgfTrXlxhFZcgubXI2eSe9zN/any3rN8+Upl
eBiZf4hwu+x4GvAxyq2dEQLC11l94+crgdqKNWwJzzNXIKGBIoo7Vtp+GUbvMlDc3+UhT3taUEsK
qHwVmoK4rFEJIz3oMENzMfhXcORC3IE/OQFLD9Y84lYHpGuQyjDmKxYpWngxv4Be/hSlsgQDgxId
r3V7Mf+/OC/AekLh7KnDJ2SNKSZjmsQcO7L8lxHuP05TWcwbzSOKU50gIuTDrr319pp/Q+UzvZRa
lKvev9t6heJcVTjLeBQUpXVZohQv8vbs89tlFUMmLpEA+w/UjN5li+zwHafWuTnJSL3Qg6DtZs5u
OxVu2vq4RO4D0NDjst6gykMCKM+/aETgFYQVMJPU6gRZsqavZ1hMTy+K6RJOx9tJalZD18rOFjyn
pNlVciXWGkhBHh0cdt9abjIbNElNGJliPk9z7mz5QR/mJWPB/1zuSspwhINTDZakIM496J3s4ye3
nBJJhJIt39A2gPu6XJ1V24se1m7cKB7dQkvXwwmJ8bZTqZiWr9+5pi9ZxMBsA8q2tKMmKSKuu/oV
ly0jbwxvSNotT1Lt5bqkzLviXeLXXq32sd4GuKaY7jmlnkCknWn9VRVTsT/838lWbN87MN+HlhFi
ICgwoIyjyqZ+JWK5dD0Ufe4W5mAOKgLK/Qh51h5hIpSXQPjF7u2f/Mv9Rpxl/g8PWsiIsWMSduL4
BW8QsrxKfiA9GRy+mosTnsytFGJr5QMzz7N9GxgBwPkj2NgZnU7sj36RbA5S2aIClwDLSR2A72rd
xCH9DHGwkdMRPSa+jSDKjOcJU9xyz7olRH7P41d0I67WZyAODhiE2+CNI8B9stMnFOqvzWzvsL5a
t6R4EH3cQJAhc7L/WuHw7Gd7bBUd7irx7qhSjbu+wTal0mgok3Pqk8QL9BIp5XLAoJ+eCmkgo1Ny
b31pDyKQ+7kOo99maj1+x8fbHcrj9iNEZayXU9dFjJUOYIveZ0WyY7pE/OC+fOBmsAsJjbzkdGtT
TrDOO0gEsRw58oSCbA253m+bd1+O6d03RluGc1FxMYJQYptK9OJG92ShHe9Ap6QGqvzFPsthZU+o
hI6ARbtDZU+tyQ40oi2aUo5aldl/oGLCbEi2USDkCylCX5UtzjRmwnCz3NdD0NdwGfbIPPufQod8
vOrGr1SZoqGAW1AdDQWtrAoUs/kdS37Pg1Wi8ZnzpF6oaGa5BMJDWfXWQkSrztRu6BDFedNfaiPz
iJtplV/0MX+369lrvPpluN9aEaMU/gD/t8avyhbsal9/50MS146BZk4bmTAqU6yf6paseghLUrob
lDn1HsfGrDLQ2WLxyupbq0KrgJle2J/3H8fCakrJPsrQL5n9aRvOSJbLWogW3AxGcNCHHOr7HJhu
jtecjJDa4Sk6DQpS634Debkb3DA9yRGTGHFKY+dI0uiojJlz4oAyTxdJu/z5KjBnPHyOsy/TLVfD
eRgbZ4G0j9snfvtgT15wbGVsxXfaV9KHXK1PO61HNXsDRFU+hFI6N5a8qg7asqePGTrPr2Ykf6Y/
D2KDDuSELkARpJ5eLCuLpfNYhxCR/2j3PqhzXDT4yWvK7ucq1I4cUxpw6X/LQrBwduFCwxgd0tUL
yN5kvmHkRVD1HsbaUL0UJJ5xakSBg0JjCt9Nn+0TH1CpLW+7V3FQAA6u4Jf1oIeo0JmsYVRoU2kN
dO48x4iVGxzCv4AMIAmSSVP6KytZzPBsxSMy0G+Zoe//fJpRbN4nneQCfrK39yvT6kFIm2erUU4F
WcyH8RmkPCqYy+XAOlpvbVfZ3G+rYFOlpeM1uf5LFKXBvdbO7B9SOy0ZSfCJUdhKycUbwhNfvUCo
Ek7Ytq3mPesEFSqjIQuTvhTYa1LxaiOt9kJobUZTfcq0WOn2wV9gGc/GyuADdzj5cpiQ/jw4jsFA
vTN45k9PN2o/AocBMbpht+FScZpHosyl8Ll5Q4T/KXg4s/ssOLl7trXGBld6tyH7s0Lbe3C7q6J1
D7R9XHjzoBQhwGlFB4vbajOf0ty/mdD3smKo8mKTOhCttnzq12/b7RKDIG/jE2rZOPfffuJxK8oz
GOzkk3M5ZeM+oziezYO1gZdzTol8dUesV+hc0Z8CxpP2kR1BrvPM5uJLuvHZ4AskGNldgAAIzv7e
AdwIaOUqn6SXGV1uMnTmSUuUdreBomzDYqqo+un/9rZgDh0I3XN9o2BELWCW3oWjKOG8opnEhfse
MDgoQit2G9gzf2e+jN7mqjwkNXAvz0OILWmdi2gMaPCgs+f58cKuugA29JmHCfsW+OwRYfIZr+UD
4U+tS3+KyIGulGnpDUjs02A1eGnPutWzwjbNs8A/lLpGw1NKwZruwDsu1yR466P3RyYgNWjw/xxN
9uC+kh+EtyPnYrZwFQjMsy1rdcsMvgpCLHtPWHjkJWlgfunXn4nlB2GTBIr9P38hBv2gzcLioIR0
CL5rOQqHhnyxbhcsPNZabgiIer92n1qK/CKpR0WXpzfqCP3008/X09wV6wEetzMREPYagPamI4nP
d6wZVYbxFrgNfBOd9d0EbpTCTntq8sA81N4zcEysIFtRVMxdBBCWLGblGTcnDqqKZpwzszNrrZPE
pyNQufQ4pzMUUbQ3rC9ZazJba4G2Jw4kp1JnsigsN0ut9KuAatgO/aslMQUiWSxa0vALgm8uDS6J
/VKQygKxH0GyrnMwvlKiDaCWwrq0R7CyUY1nzAgQNRjy4OS1oEzhNZULcPa2AiWLGM0J4REoP58x
xgXTewz/Y20arTFugN073JY+qKalVz7rxNqncNHpWkyVsC/urKJEGjGX6/BkRjH5vy7HL10mSmoo
tii/xk27RnvkbaIPkMmsThZmpKEITuuM6PeeK+24l1w/6MQb2VDDyJ8zRq3FMjZyQ1Ghp9OMzhKG
Xnd4vUp9sfqTAfCgkZ+Gr0Fz99OJ49/wBGCT1tqaapQVHweWGQCJZKb2tm7cj+3ewHcXTyNREZYg
3LZQXrwCLS4Ka5T53W9oWllcn1iDmQ331K22nuM47kUfuPBFSSAYTwSdqdH5lF8G/KaNXz0WPka1
jFqv390PV0ZGFcLRLomdnilYt+sXuUjltQi3reXGf9bIzm4mmJ5BuhQyYvBZx3pN9fe0ruNMLRrQ
nUZU2h/8C3h6b4txqR51J+vZFHlT+UfNPhOT/mdEfp3BHOyQOvHYTEbfvNyQMrCtntUvfCCSBhap
ewPerZ9/bXss23+nVGBRGhd7JXmynbGMtYHzL37UXo2NPLTdQSLu0nX71NjsxeHa28z9UqsM8fGp
n5mh5ainsY782NZ6CH48GRnWcRHX4zwZJyqPzfX2Pk82uEjD7aynunukyuPMTshYJ/XXn3yyyDq1
3F0LVNTmIfo0Gvf/ZwsJTE/ys64+yDCatFotLGb4mjNetW39JklWtUEXZqDA54BpAoBhSE47xs6R
JCF0hh4uKpQvF4bmiSSD84Revi5LSLuLVX4zKbbCm/lznBFRxSPjuexS/ya3CG3WSNZpSudnpLCh
eggDe1XXXuTyj8UJvJHR+RCdehxDaUmlMukXNe1//hjnSrO6Bk5egLAebSpJ+/11CwVT/ux8w62b
Ibg/2Os3KV2i+8LsElqQbEYvhEgvPWAwGzHndxshieErY3ToMoriulrpT0CaBcZS5gJ2jMD96hJq
qonEJdSxMZO5iTd39vxB4BRfIE0r3aHrS1RwhkhXUlME06dY3lgu6QOr1RQjq6/5OuOjOYmEBUIf
iiK7Djzza1NWwaFE1+MmpnIPfAeXbkvw++5YMiGIQRN9EvAv/7ogVddlq8zLLKQZ8uWnDPkPik0R
cM56UJ4iG0p1R8v0jvecSz4hDmDZodEFxIa24IN1S0LM8KAjdY+Zc1EbKPWNgQ7z9NbBMvgR3AsE
FZs01123JEsPAaaxK53S5dfuGCOWkrS3k+yYarautCNnJiGX/10Kz6VR1mAAt0mbDij9aBHXTbDS
+T9d1WH6V3GyzZKZzsBseX5g5WgGPjlLEeuuNUkPS3H1wEQ8n9ee/WIBaUUBXr81Yl8ILuWrwD8j
qdS6nO8gq/UHew6lomZtzedhk1/0Xu6UbygYPjlHGIIYLbQH8eBKpAvp3FyV7cr1HAsYO8rqHGIS
toe6x08B61XKMkJAFhkVlxyJHRoXVCMFO7lG1fhx8SKxAC7Qt92LjhfsXjTgkAPjyXw9rsAaLp29
sbvRfOpncAjybjBRXepeBISFyOya06zP6HTCsXQbm+9cMLo6gGZwCgCJUiaUcU9MyFoMBnh7OW6a
Nbf09TZRpNEtCPH6lxL7IIY/Yk6z+0O/xltThI2IaOqgYU1r6cqCxBHdnDDL6gYWJFSRPxjXXNHl
Gjd1rVv2uW/dQvu6St2HmM3SjpQxuvPovwfzsuaXdj6ax6fIdb0IoWQAj0x/A7YpOQiOyXBMi8HU
kfsoWTHIUGMjBv4Xan2X7LPMziuV1JLux/7dEcVJkS+B21kdIYNWWoU5nQWuRvyFT9/JE5ids7ko
1UbhHLU4WipFT181L+8OvsDHNFgUoFZIYKJwNM0gZl0R3z0p+1WzhxLPNWRTOAp6dtSaD38YHXgO
3s0LS2uqeLt7tvnf1QTE3c0b1Z4RxNGtPvrGfkO8mkvCFtXU0XDbB7VChpyWGcH3WM80RqQpq+54
Ynv5B88LRxyv0AwnOtNdDZgxcnt1HP50QoFQC9CcMv2HYgEvqYr9yCl3w2jmm4Ekm3JsmjfixtY3
OxNX31hhXLfZTuufHCW/ByihX6F1qJjMHm5/oVQWdx8fLE+tlpCdPqa18x/KV5I2Uo5NhNRf3Zqo
wKl2QBV2B0JDPSl6VlN/Lk71PwwIO/1wyY4Iy/FD9Nl9vnWDiuQ1bLkNztiyQsukYR2eGNXQyl9W
vtcu8iL/Wjwz7muM7lAGmiB9RdU5JKiRXpLhti36nkj3JQHFLcjDNQUp1Ilr/xZiNhPxHLth4DAM
1r0lxINjHKRcsCiLlI2Dbmx9uLwGeQMY1zqfTeHt+BBYK6F5SdPd7/hyeWzRqVFy9Kypp7dp/6gB
0Jq+hxiGKckN6/O6MatrLjC/lHFn+a61VftFPogrHxbSrePjh0VaQLSGylu2WNNMV/T9UzjdeNFU
MxeYDv4+3QAEtax9XYaFu3PKCUkacRySDJGAdn5GIFshJTg1WWY4KCEcMCnaeWKplnRboaG7fzwg
y7LLg0zz8atY+hENDHyNByecZzuogUGAQ9k/Vxz38vp7v1wulixJ8RkYmZta+shQ0X45IvEdanmN
wMJCvZWkgP4q3h8S39ol9HBKShYcn06C1FSl4nwKkZDOALbX6sdDAcfKBdnRrNvZf/0CGLAb3aaj
0+4wtX6H5m+syn5+4R0RyXbFGviEbamEz4i0bNqC3ELm6yIkM/Ozp5xgmQpkmw4n1an+lwDNWDgf
425z6ynaHwdGGt2ro9J2687h2Ma3fUG54bgmh065dCZgMRDGPYs6YAMpfskaA1Q2j+yv7uPFMPGN
pVtaVS0EWO9iclfZsx/I/zUdpUQI6nQKd7E2oHFOEwq+VUy6nDdtpVkQXU1Pbl560Xa3syqN14Ka
gbNEpD9xXvKSO3+RPyG2NguruO/tQvLQ7BxLCgpMGAz6ie8Z4HenbmS6fZJ5iPBv3Yx/jAkzsSIa
0UD4QSh1Fs5gMfq5FxLW2zGprLE1k8HYDG//v3VxQ2TYSyanRtiv6ZR22MVyCDBjCgFnoHbW3Nv1
AU61/W49CpqsDOqJV+6QX88HyH510MCHLU51TtipLWLQtpF+DekZfhID2xAnKkbCrGCpCN+2ZZXj
9kvXygZxzyzYnyeW9X+9DjZMCkyprQgDA9Abn50BoRQWKm1weY7uelFh/BBR0kPCnvjy0k74NFnd
1ABUwK8jbzYLlyKxqlcAcLcVkVTjH+6cTYq/L3h3N6L3jLWbswFlaTgOBiv1Ek8X043RwlIwtgOo
D/mPJrknA7ub26udNTNfn8NE0CyZq6ymLJcD5R5EiVKbgZqafqoPHCeOKh0lJeE71UfXT4V3D88m
J7hIA0O6Dp03GxQpSwEfdOQSTEMqHBmzuxVzyKnayHwuzZSv6AZW4x8F9G3TFMJgahvQwci9zv5s
miP3fWz0k0CkDpVjGScs0kdUt5X2FJr8CQqLhKJlDeNpMPYjI6WZ0njmMRR6z+e3tRc7Jq3M8Rog
dnFd1Ebpzel9x1btFwSUfOogZEdJMxlk+28eBtq2uawNsfdphcL62tZl4B9H+TRpWtqtGPHhaNTZ
cxsxuft9NsqsfU0FIRMXLm1p8YM4tLCTDedpOkgfaHmwlouWaeaKsQ+2f6T3bvv/Rq4cW9GfLgeB
szyEmmayEjNv8BhiTA6wBAsnpezBRn7jCcSGqIP4GOvvYDl629PBzos4qGsGOqryrjkxXqTyKX2c
XYEd/3AXjm+oqfh63asFbkp4Cac+j/aNAOx9yAvDKc8Mehb//ptBwuCGTvoS+SH0hv9CCAqhatSG
TT7qDxKm5iFn/IfNSulgA20uozuzZbHgZqSOjqhJDibsiTvuZTa1YZwbJ0np/6PK9Hcx+svTTDF9
ADSlWwDnWVx+Ms/tqO+2jbZlI/eqpH4ZnsgKRp+HPTg5/TZaOlbntCfOC6Zci1z7mWmf++M9W+iY
k7YHElBLdGT6ZaGXPDEQZ764SAbHscoj6v+wyKbtwrFOxWxMQ47nUKRHt4clnYJJQCaba9vvSge9
abLYGGyADPFQyr3OQXXLRnmHTDhtVjx0lKE+IqKfESd1O8/Wxfdld2vRsplPle35EA8jsFqcWJAL
f81FpYogfhUFU9nNM7EqmKnI8KHiZx1RJfb58HA6waXdcjGBTv4Htx/lN1SXN6xqudOoeAb+jCms
y9PUw6UdPxPW5lnnsMp2ev+YyuGsni4WVEw0h/zLrnfNUivVDRpGLn/bnIfM5PwmUWzuHiomzia1
5W3r4zeCqbjtYWZED3kKnoqji+9y7o1o6nAyLmD8jt/FA1t/8uxRZQfjg92hiUARP8Ia7qpKM/z+
qTHf4wnxn0hY031K3pJWQQfdGn+Fn5qSvxhnNhl8VS/lfBpfYnp+UZSqiU6kZpzewSdlSelJYggw
AxHaJAjMxQ4Wezex6iaZD8lIBApBNCgYBWtiUVY9MdyfiACEnRsqNagmrQthAsboat+5AZrP21Xr
ySGRDWEUn3v0Eit3zKBrOKYpoyrXvUKhCa3x6mrqkvWBOMh2LgfOo7wrXFfsp4xtWL6DTvRApRqa
YEf1seOYQYTj56TXF9GuRTRmn3JWIe1xrfpTYAcg4EK8WkOQfvFplCsJn6ntxlk2V5DkNmGfBRon
yL5lWet4Ypos7jbXv8hwd2CeFctH8RwcU+DhgoC3bJqcsKCP1AKmBVo3pmZk8zo/IOxHuhs3ghqO
c3FujUe8gxACsrZQVAFZBkxTm01jzlNc8fLHpPEWTiPAAUe1FZ7DL04YVNmWJMKNsx+voMZgPuvd
tkYltb1iyEJ0L8VHP7A6NWirRGqNogHnEO/9oOkTXJucF3mdPCKsy8OUav116HADLgRuSXCXahrz
nqmcj8JI1kNqBZeJzLUUs1EYJcV4sM1U2IOE7dEmzTPDPove7LIkMrA3oBv3pYGr88wSAkXqOqGB
BVPZFpvLmfxBsIlAR141UU8wlVMvcIAtVCUWAeq4dWC9aySOe3ARk0i/Wl0YhnYaXQVD8uW05uCw
vnCcqyU/j0MU6qSNKe3IYISj9YVC1tPqiL4TCWE3QgVCsPZdri4xBHZ1ptIL2sqcU66Yxp9rey+B
Pxi9XVeHHvyZ1dY2dWTNLFD8m7MUtaufyqCBC+v3G27C+r8953MtN42kHhIPhQtfs4xzNgx9i7Dk
yENsahYovES74/eS5D9J0RSi/5WQMu1z6n1TANl8uFS0XC1GLuEOfTo43CfZz1itMHyGieRqeumM
fk2Rf4UKlCbrHcUFvnK0yYzaVeUwusZpm/fWFyfrwkZB5QoSon3AJzyMdVUSnUQl/EdWxpp+fbfn
pSd20sIOsR6jvaDI3yUKWdaEZ/HNvRJacJKVHwmqOXtytymPqjodhtDfuxqyf8iKoqczyR/NRY6J
iFeqB3JufWaP2pB4a4fSpOPhP7cxdYWTWklStQXe0v49TtMQfu9mYgf+eDn0s7csEKEV2Vv9RHkr
0Z4DC6ILP+2wNl61j41O3NCsVdfydRpcPd0ZwdRNT36PrBOPUTTJ3xiFgQzBsRrhf4CB7P343Kgf
dc5xWgbFO+hgRdyVePBcHwkS85wG1vukCHBVmzeXM9Wy0fvLvZxqcFHuDh33SleWePLvZDNyvTkA
t6al2mceSWqHk2ut5NDMZmo7mr1+WRTXUrMqeCHK3EdYWZt2QqKBCr00DJZL32CfcL8JR5E5mlX2
3YVi3RAt0/rdsGvVOic+EONgQtulh58yTJbjov/Ro7JfmrhG54tz/Zsyzo8AIHSU4/dIPbHrIIY9
s806zbWaXDZpo9fOWywjhHXLWT2+VASjSwEZpwVLqCiNgH1WK8K9P0iv15J/LtQeGhYYB/miz4oS
4ZEzB3PKLX6w3ahcwjwgMnI48OUtTdfqKGxftp/wzofJnV1vgtNPyq6jKjNzNPVswXuRDCGqjgUe
7sTou/s0l/AYoBDgZNpba1LWoWa684yHiIvojfeuH9+slem7uJwb7V5vyAM1i2ZrHhZviht6n66X
O12aQdWii++06wTPTxZoyd2iaUVOYGS2NOypxrd/DLWQC+ypUo8W8qcD376j5dw0M69gBpuoZK/A
HYRj4TQm7USTX0lFKbYpmX+3CMBH/ynF4tvbP3YRNNh3ZDEL6f2QWJF0orb8m6NIkiyOs0yRtSqL
EaL2Utsa13mVks8twBokf2bwTfu9pbbTZpMWFsPWPrX1xD+w9jg0uIFfT3JEa4emmmPPdGc5XSfH
szNOhfhRGILlvP05xlbxX5mcIHFwSt2DACXwc2Ti2YNVj8uUrGDJA0nqYxCdvw0G8c7UuTpZP6xp
e8daBSzB1+rZS8E8BzOao0LD2+3Ahxp92RAIraky+4hhy637+COb+i8dNSxsv21Ae61l97Fa6hcl
UNOU9LxN7GkLHQDGsdgYYL0ko7czaF5dMFYsYAd9ir0A/VULFh6JYDr635mt1+y7VEh5dLvdMou9
vV36vz1I/7j+ei4diQV6Tp18m0PAcpwZUUhQFcgfAdnJ5GQRyOaeEOrn54wsMBL4eHwDQDujRV9q
P8AJB2ORW6m/2rGxNXxwos8n4U3EcDDnU8j9gR4rbsY7alFOfyX9vw9Vs0DnFkoIc3YSVwVKkz2q
SGjxntp0vuCvIqExJbShqw4B0hXiLtwqyPu1BBzoPR1A1ohQBV1VUM6ZgnvFq/yoobWStqiym6as
hheO9IP+d/7f4okFZU+mS8bqF2TU+swnol6owcLJ0JJ+XScbqko9PUxS0RVb2+jwOT7kaVwrMRcZ
IUobcYXZTheJ1cgI3q+RK/4mc8g5cDYj2d5xMRgzqofb9l6mh+0mFx8X8EtoPeINZoKYh//zw0E5
fUWsFAGjhgDefayyBGivZ7qac4e1D+/TXiq0/8Q6xvV3YgnKrDr3gC5xqmgmvzyK/B0n3/GNaiK+
deSIR8MACPC7TNulFY8iVDApqSlu7JfnFUpKy9MyIaUtA7CJglwJZ2OX3beSBHPRdhzUEVBZjeuc
MPxr2PY1mxzIMABcELOIUod3RZ6B6MDrwL1s+Slo9Q6yxgsCSX+Fqtl5t4BfkPU/tL5mZYIg/HPq
xWdb35CzR1Hxp1KO9ILKsB4D8QZjVpWVmGq8UnXqPEyI8nvsMfkpuzcQtsdQZkgN2xj0yrKHugiA
iFFcD11EpjgKIrX+rgMGaVv18oyN/dOfEx3lr4XK0tfAuJ+Jv3t9TvGJv5b85XnFUYWzfF5jVz0p
AXzuYgwouzyjkP2gm3VzcaIaLc5sGuHXQSvrUZ67mUm3lFmsxEoJE8cei/vPDh6hQsQldh5ijg8k
AOUAiEstzebAw3jZmRNjAVWaK7+D9rj/WsZJteA+Rv2GaOkL4qvk6sLrIQ2pDJYnrnV7j1TXe7Sk
Y0Jw/aKRVsyBPYLWJX1D8/kClO4aCj+SNu9ymj4xMxAqcKAiJbHuCXbCm+8c5s1qOXLOSPCZP5wx
ojGu64VMSr4G4O7u9mITxi28yJv12jKTLkcjXAAoV3zyMh/mJNDuuxAHgv2vqWC6B/d7BUPVDSdH
pibqSJEqAUiWUHf9i/oKADUeKgZ7r0abM0AzITc9N/htp2SrI2EnYYm9Er9gBUrwNNHMRZ8POsG3
JnhVDovi8pqOD4PfTYu8GOxQw9HxgWWcPchAMCcgU9RrtkpkU7JrniuGoBI4xSWzWhMMTp83OeQX
9V+x1cNLncbk9E2VS9FWZlfSe/+Gn6dow1KxqA1L2iZJyoOft3bPdC2zZUHtoMmwMTKuCvXHEsjb
ab3z3jqjR20+xezaM6/FY1cvscIqNbmMzKGNa+fflJEcYzDnNHmYAaxUrTDuOt+x/hF+Bot2QPD3
Jay02/DipuEhYXmCXmyBVfBuJC7bYA962w76w1wiZFYC2rumXpy2aipiP1drY3LzEOlVVNhzW5k0
fyCGpjrIU5owVR9yiKsYx1Pm5EAsMEvhRQY46VZ6omAAyl6J2o8eJLEbj0FQHFshJk6kc42lgyj0
3FT6Bc1jCb9HjZzKwKtM/BsT9ksjAfJq+rm90JbHPZ1O+4Kz+qh+mgsiktzCagjoR1FbzuJ0YQZ3
IVx5TzfJS+aS/8Y10EUE+orCLylHZTlM7p9VxWoFzNi8+91LAEGgGTwiW0y/uF0OT88vddSq5/i8
ckFgGZW6gpjRDGOQCrjLqJSXZ19QNI83e7+eXRhZbXntprmAAcVdg9r12y8V8wuKRtKftVMuWZNF
vKO2Q2GXOMJaVuqCAjS23dlKTBP+kW4XwtvKAP6l23iB69/yiiuTWxg7kbfl2MjwK/0vhV/htDIf
y9p+ItV3Jr5tGD4OFnMMnjrLAfXpXZae514acIOc7m7gHeLGO/4AMkS0MMR2RRAKXXQ6PtonNbhn
ANF/3su2VLLgmAjgmf7X8VeHcAFDqM3QLlUBpikzZ5b+fB9GBzR2IJuRn1ju2Ii5BuPSz7zvFVpv
eIHyAiwowegnNmG3pjqrzI1FHy4FGHVCPnCsD7dy7+w5TSHl64Yggv/xUyHFKxSfwLb6DpNRKWED
UHrrFJJPiIYN+1rAxuX+xy0pxRe2vwnik7AwMyGNSXotiKsQXehaQ8aTDbogOd9/jOz0Xj4T1Yyc
4hnjvjedVpHGU4EBgKnQ9InUZJXHoxbB5rKmeJ6vXCpPZR7OUmzmMiG6xdMVaDcjKsbZ3diApQLy
4HLBHL2W0qDT+OrhepBaJOunfe2rKwxMIAhORK/jv0idXTBy20wdAdpudZJP+o8RnCDArkX88Ksz
1quZ+nPSgMXwTBh7z+skgA8Q0Yb+2oE7/yry4bIEIgASkoBtCkoNP/vzAoLtRw/jE/d1WzwgcSm0
sWfkB111e7sGuVVFI8GrbIL/p7+/Z9Y4giF9edPnS27Ogd/p54msjbrmA9PRYiU2h/RL5BDO9g7+
cBSDJft5K8vxLz644WzTHl2Doh0i600lqiVoK6YmtLj6fSFTXdT9LNUy6p9JYazbPCkBjvF7ccwd
mO9/zP97pNMQNE03SGIV3Wp41NfUDgPJvryiMr1/js7K/AGsNx7ZMmbQOrJvjSxbkFVKbEXwpQN8
Vjhcg16kYGyvFz08HVI+iw44W8dbvYjnwYjnzelqwwfQ7EbS8Wm8TtaLPH7mB380WTW7Av7XDxkx
Dtefz0y8obP3VZN+K3uXYlJwHGNuuJk1tyugiHGsTUQ8porVEA+tKfknE8eBuhTiS/AaQqemdG8u
YLDP7ayybdk1xEoIVXALjuLNp4om+0jBGDnLrMy4tJFaDqRPDxxdlQCVm9Kpwnyo2jcugTfYrHRk
+RttUg9MD227tgaTXXRtx7JjIAKCvr03o9IcGCG2ol78tMkKoIaHj0DbuKbK5kP1T89jF8DeYEVy
ocLTJH5rjoBjXFXK/WPmURC3bfTY6nsFJv608m71rLTpBuOeGo4CWyNF4mjMZ/Kodez+IRguxK0q
KX/OZWDBzDxs8Zql+BfZDppljiZEXljHO7OcE1fqHRhT5HIp28QKuf2YFwSdUU80rJ7tYQL8YKzX
2u53FEnGg+wHEBwTBfW3M5Jqic1UTgb3hsUBKbXh89wsxmKo0XrLlUt+ChdWLwZ1866RPOpOSbN9
juWqCYondvIHi1yApBE+9TPl8S+XPrKnGxsf8KC69Hf9SEo8TQd8MFP8pic5U75ZbGUFh+jxPNwH
/pzWvMPMu0esy+mYJq5sJJPqk41y8viJriN60JBh/8gh3m0UBTjL2d3vcmVvcbpVyolNGP/gBFbm
mqIZ0IGKr1i03ZdwbiU9Ndi1YA3L9W35nOxcdGIe4Nj4ssnLO/EHZExsdtz1yxRuUaZyfPyWvoas
NUX8Y3vm2bu1eiaFcwMaIrsi4cmTqEhOThbq3+wA1tWAT+8w898LoDQM48koxNYHFLpAUuC4t2VM
8I1d5H7pSipVwhVWs6jTRimiTl1kZirPPXAoIWevjVPIn1zaAgQNzqKo0YQRsYwmPbtM3h9VcXvF
Jkv4PBFgCP69w3qgoZRmIqjw7Rd3X+gAYH+SUTIN/i6Sbnw7Ca0g29InoKROmReTMZBBnjCYb1yD
hNpHblTK8XvygE/A2N2yp5dhmDNG2hLI1ZmLPKFykWgfnTXzcZRk6o8UM3BaIg93IOhjetx4uH4y
a28ienWK8//4YcdRmHRCQl7xevlIoit58CNRyavMlM9M6pRNb1QelVkVDK7xoIF78qScOH3dWTu3
NMRXPFmEzmR1x+bEAc7AtoFCT/77x5qY+V9kMZwSJ3PJWfqtTezZmz7VfDqiBy6oobrz9E/QW6/M
Sy2A45vhz6XTwlZeSLByfoZ3G78WLxxmyJvdyy/Tsa931C/ue4xeVEkU/xm+X73phebWWU1r3co3
gD2ntSUl5BXwczoXZbNJUZWq23qFxkfbYNpd9eIGfhF5ZuCsRjk9l71KFKduhfVfM4wVy4TNZeSF
OWic7kE6VZE0Een1R2sN9j2p0HTBqUBDCVBvJ4GDVt4ELPKPKL1B9xlBCfqpFfSKMicbr+DfR6D2
QwX/MQ2yIOyKEhMpM87WGueKMnMDEqGPesdI4CcLdh9G8CSDxM7m8bC1QC6I3FNOejmvuJTR6AIC
jPGzTnfz0c3w4WGejRjXe8NtSvmxeQ13BbVMl+cunyvP8v1fgHiKESSy2kZ9hKxlr9B7/6UTCeQ/
BogZBzT+5kOi07cibqsoy1r9ZTz8C1LxymNx/BbzFnaI/1OzAm8UQxm7gt6fgWZutbyXckv+i+Ag
9J22r7oTDImTcRzb1AhlpltFza42qC1gRVoW8YHLmFgbn/jW2F9G+RfqrYHG/5jMr0QbnU7nllMF
MDUexvr+wVJwrkfNgAYFn0hPdrED1GF7EW9KirW30s5+eB0tQy7TAxJEYKde309BOjT39weaKcF5
0txAGFu2CWpuBFWaEl4VJ2KpSJ1HnOcdHYY8KdsHHN5Tvfyhc9UFgP5ZhM+BAIkYnB+k5vuMgUes
U9+rrAQWj4GJ4dvQZIlZ7pkBKEJxJWkP6Hgz6+fAIO2sBuq+I/9N/2umZIfMVU7SkXFfWPqlG5D4
9WDElFRmYkDuh6VvPVQiRt776R1CgRQIop+1Gd1gPr3ptZDgfoQRuBXhCzLIyPUIlkCm7f2XMGap
Tl48R5QOjV1LZJZI3LGV7sbDjW2iirlPaaY90LO3eWmylHNHoq4gYO/sk8HB7/K9BWsAZebKXFWJ
GG5ARaT1Lc8x2BfSiCDhUJ8zlEQdgz/tyyIJsMvksC55VS/FAPfIK9QwfwwfHDp3CF+8LlKUrswQ
nT3qG35ZTE4k51LAudU1xKzOrQXwol0WeDQE5MVi03nKsBIDXKrOJSzAZ7dH0eYIgrn3yORCTdtX
0tasuX3MX5XsPkRLCYdmolvnGfELKKA6EUSj8TsMHJlMUibW63JWOvPoNqo/18qRSxvUgqAlpaHz
5+TsKRA3Njut5e5I4nYXhfkWeL80rfjlcZAKWQ4RgzqYOagp8gLakuHkD14gPUzNjBhSfgAnRQGP
N/qU7sAX8zxzDct9d2R+pyBw4ySPaiV08K32/GDkGorPep92lyNyDAb9AI0fN5ULoeO5VqYhh0uC
yL+bmZiSArMFanrW/KUIBTP5sbsL4Zm5r5fJ+KKUzw9YF7yv1u2Ix8WRFKB8r/LNglFjOkWGtOCk
lNhYA/yvkXHn557GIyGun0JXbJ26LBaU13Bktz9HeDQYLg6Nf50ljwtr7qaNFOTYfq6nf35uzKkm
ETzpWJysbNjQYDVg/oSE6UJROKQ34aXW9Ot88atMIhb+1k4GzcAFtDm92Ve4WTWzhUd7BM+bFUs8
OadKHmJ6koyvobEM7w9a4qmY048qAfh8XJa8ZKCq0vY/E+O5wM3PyADVEeksmQA+s0TB+28lJ72l
wpZrUrsOmHvht/0nP9lsY3aZbQ2v14jyAaoI7jhMIR75Vrch6mdBmj7A3KIBImps5F3/iTZhDjlB
p3bqPMMYhwtxC85+sXKiv4Kai20/ejPgWRPtvV7FNnKl/zf5SRdoGuR96YJNJQfzLyAqUBYK9KbV
Fp3cqfJGhVTkiYfBUK/0PE+O/vfTCDR7nAiRJk2am8Z2Tz0txV8Q3BtHq/+W55vPP4Y9zhh/2rnY
ncgBZKdHKMJUhBOSKQfa37aNEzTYVYaa++HAIQD0sQ9y/vbihxtw/3Z+a/gceYAtV+sgjMOw1Hzr
8u+LlMGUSe6xFaoau109/giZX3zJ2aV386Zoh2sfaEd8fy7gvn8rRxSYpzhxnZtX2RWRSNyZr8MJ
UEbNNsxXWKRdQTZvsiTi+mt7kjv2NOEX9+XnaXxAU97FM/Ri+p/nghQJr8SxJrsAO5uXX6iv1Seg
biWOLkK+kqBIpgR+Anks6BsY7sN0YSryXdpWrXljc4iVdZQe00mYlWaZlWu4cE+0gf+z2OIT6k5s
4TBLvo9yKtkyVewWk1ypDV8EM1drEFdHVi6rvY3aUgLDRjKJs2s+bfzMqkstwDa3TvN7XzX4y3L/
vvNPJ0BhIs8/Ft5HB2v8gZtKWzD1YfmSSx01kZldC8o74kIYtHkzuxJNHJ14Y2A8B4D+WSPdSOsv
MN/6J/2KrOfW4gEVH4DfnYRGAxNF0eLdv25iIV4bNSpItticlf8YqIYcK9T5gQ9pi8wfsTFjnaCC
UC1RPBWRLN6eO35Wls9eMI2j77QUz7XtDcr1dj+VQRYnBpD/nx5KjGRkmKgvGacEdbV2RdGFhEUP
LYNdlQez4R2DT0etx32PlXZDN7wy7447i4I+KDS09CjABwrJDIkffWTf60IN4ggdW8eDnep3xZT6
rzju9TwGmcBm2/SyPTzBpfkLBvxqmGfa2BKO2/CCmSXITNemZXSNNL9d8QH4S4c8bGto0s6SMThq
yDYDYyL+2hZbCv1KbU29LlM2jBCuSeWODOFIj40n3BF1xlTONzt8j52wCcY2x52StiDJ9hmKdmXu
BtlLchOWzc3+GDZQGcRfk6cPg7O1N0ll9PJhnYTd4Z3ksX0mV2LvuEl2pr818boOQwqZBxGu2Edt
DGNAPfgQpc/rg44HNUmAWgc60cus4wMBTzOxhDjQublsF1ZyoXVN4KIGx3sr/VNpYEGGHjt72gFi
XwXrDIDiIN3OIpbxiP0ASnAXuR20uAjGlr2uFv+wZuYRnKl5ErMbAmW/iFYPU2pITQ0+/tlGUmn5
BUvl+BH2YgnbtbHlySOugpjnv9MPyCTcQLnpnA4ipHEIcvevJtFXlcq3QkF9dqt4UJq90ldPy3FH
ogu2w5Wk4dAJGvG0DfoncwGDzld5ak1Axck9tyxOH1dWd4Wv+1PBvgQiNos/iihoz8MYn70zZi0B
18GwOggIDBLjCxZ+CVSjVz10O+xI6H0gc7QbNmIyAqCo8kfLBIHbwfdJ8ixSLly2KLlQiGs/KccD
zZgaitTni5wdtIwOJPi5JCLxY7umox8iTy6YblnawOjebZJ+rsBYSQIb7piDqxzuQYiJbnk0apOu
RwL4+VweWS5cw54hPS+gd+hJFQXRoVpsAxlBnF5et3ahNwxyG0/GE2qNqwU1Rmd660c9T45ses28
uPgrbqcGmNfTjmkX0BEq6uW2kTRrC+lh9Q/ppnpuZ5Wl63gzAwRWN/1/qgPDVYAVcobWUDSEzal/
lvm99ZC4dtxZzS1H/2BT3odzLZaJBWGkwA45bSmR9c4l7Z9DI7CktGlyXKon+SO7FPZ+/FeeRMRn
OoAikDTQNXvkoWtaawp62CsHbgU7YJKoWb1uIGlH1ATormqKZBY8AFRwfgMRwLD9hEl8+edLwm3t
hPxrIonKluAFwcVf9XhMDYpZDWtjVctdyN5OzyKosYRSVQ0z94yh092W4HY7uoHELbhEzvJNRMSo
V6YTM6jGWscrBT6bEkHMzG784N2VvcpGWHtfQZsEr+55KamEmKP8EgcCGoTW+qo23jOTVpybnoUg
SZ8MBnPo40fpb8N9G+gO4JcD/1xqd+9Ko1j7S3oUKwnjmCX1YP7A2lOSEN+QU+vegkjPeg0hnlvU
VK8y3u3kzHNDMx+baILHA4QH1YwCT3U4wLivS4NvwXCuHMQlyzhY3IScbD1R72iei2kSyGeFtwwO
sCpzJT4uWeaVSmcYIW5Lr6iejzeXARXJortMWPtdU04BTZF8ryLJaXObsnN/6FNbxeXI4ADAOrAl
vsV8Gtb1ZKyzd+smTpy70dOxLgbzeTeFYtgHuJAhM3Ua6kCSQTAqWHq/lNE9cPtES0q+P4VYr5Pr
p6OvHHl/6hnGrU/8lVmDn6L80KKA+bEBXAHLjTJm+UqryD4xeQkpH/xyLBfkDpnKXcRQYf4bLeFJ
of72NfNLjelyBrKFcFQPfGvbsm24B89xQjbYAqGIXvzGSneOpmaqjkYksDNP8jPC9GBSewojljAX
PTMvHyyxe1qcX5AYeqNrdEMfI4jRrZSF3VVdqtEGB2jwfif/BpVksAmZTIx+WKzG0mrNyyN46t7Z
b/mCsWzgr6GzLSCoZGDw6AVRFk0CtA7t3wglGpF2+iOiOI7IVfx1JRTeR7sEaAiLS/bnkiiazzMA
vSbsAkrTW2ohlef7aKdw+K9yrcKLJ+AyPGRtzzMjKXuxyFbGRlCVzC6BeGcXTDYy1zc0Siv7tTrL
P374hO5+3UlKQRccSKDH6+NSg6P9ff7AZcNoD3C0JlGAfIsyHIP2gwvSf3O4b/nQ7dAgNM9gJrg3
NxuHGUAyG6aABblu/wQQb3nJWoVfobtkQviYBTZRgVI3UoHRUw9zKGrckhrJVQFVDi+bC4L/olm+
IL+XKPgyJQiDxgKoJ4l8h6bgmC2RqNb0IGCN0nwlCDlXTPdaekwp5H2GHjhbhFUYa9JtT05eBEIH
y33h+0B5alaU0ZK9c5YWDWTpefryvS3Aii25QnDOGehPtXLwoUChdeQ9pXIvZDH08o2U7t+x4sI1
4Xf0qCwsM2uj/Nlwy/O1BHTbWICOp8DnmqlVekW+cO2mJkV8jMXQcVTjtf/ErHHVFtjsx783HEQ0
x1YBDjoOpz71a3Q7XqhY/npQzuTLpXYoi4UBjo/a91Kl2BKLsKpZuxunfdaLHHDW0C5TTgvDrPcu
++4gAHRZ6TdGABJ1Ks2Ow9yXZrv6AYCFASxwoV/C1txZZiAmqV2Xg31OHiDw1++dos+4fRif7xMs
XO65QTmsPvrU21PD5cAY2HykkUwgGSLqy1joV35X0tmFModUWmxQNOF7v1zzFCbeeLlBnmWm1x30
lpEyR71Th8bjYmiItiN/fNd1bBYC1LxUBWPiriLDT8gpdmiGcbzJRKlZMNOXrVQgt8+2MUD7fobv
1yLpzhbeGCXRsMRRZ+p/HMSOKy1FI+EkJ9Cq/gbASyCIa6ACDKz3kBT/B2cPJApJo/BQFQrcP0zZ
P2624wPLzuqHAh021a3aaHwBtEZub6cBGzGuYlDOrk/1UJYbu0/A4v1rTYzXPhUTYYbnopc6yPg9
PMsRH6qHJGVuE1zmdSKkKX8StJKuhcGg2Zkg/TY2zt757XwilxPziB9vEXU8tZPWFVXilGPxwXY6
oEwjQdoOwyZLCmhhiqvMpDHuRP9FH5FrR8pgyOjbm7CBYEUXL55XQ4nCXcM1q3oOoJIk8U4NkbqC
yivK7HlRc/b7zkluBRYQDNq1S6deGAQ8FmuTZ4eGBL1hYlsfUV/CFvR787wnlVLn/Ye+B5u26sDJ
Sr+B5AyhEvo7DkB+I8qJ+r/fvgi4yefgLUek4Pt0ZmuKtTsV+4FefE7W9KsRE7M/h2LzJDHLdbrA
72tjn33GIUtndY+99f2qR+L0LqKSvfBjW5JyDDnXE2TYudSN9K4UKvGA4GTGgKMGzSmRfRiqUFC5
/tPsLPPrXp5ohWWIlgSZHnwkTyKEy9/JN5PbEFizFAuigrNX6YxezRhhpwXaEHQKCB47YxRSWCpC
I7VQKt3zxMTnS1dvbNgcIp7FF/pXtRdEvJKS98XMiAax40GcWWk/WX/eIFsRQopyeucMEYZoBvrG
E1HfZgQAi2PyzQlplKUm3J3u7lQPCTwB4Yk9GLX6d1zMjz6KaXknM2V2ZFNSD8Weii+g3teXQQxm
NCQI8KJMyGibFbGMvNDgPaclfGabN6h4wmKOY2CpQQdVNODEZL5Vf60JtKybKOctrkHXDlN4YsBr
LOT+ePZCQnQwtah8u5uASMpKwMxI/hll6jh3p35uPhUix55MIjSc2zFMouoB2okfhfTgNfCisNBw
DFuyaZkO7AYw4IWOvK/eyXwMPmXjlgMnLkQ3IMf5HqTGUDV7lku2gjI6k5+CMdvhZF5ppupNu8uD
LewT7t7RLqxFydjOs5ylQk+rFROtsNUBptCl9MuOZGeM0nQrCmr+q0JmdxyuZPYE3EjzHHGGwk0u
PI0qXAa/fykHX2KhMCvtnq+yyXO6e99EhG9n2BNPd9PVZUirh0mpkHSZzY37CxmHi0ukE3qc4Pqz
kGCoxUHy5rOI+W7Bwa1QtcpKgkUrlCg9g1haiGzgmRkJ7Xo4feXOXWPt6/qruVHLnWaNgwx9mNhU
yAsPaoRzzvQKU2Xd2vC8sNqwR8QRUos8WkFCpY5KB1i/x3GkONeaOh1yvlhpMX8gRgBJGVs1z8vr
af+I/Q70+eLlcmvLRdrJq24iW2jjfYfPzcob+qF02xBtyda7HLJV42AKzb2x4OepOpowJtardng5
gHWngExNqd5lzWPlkMArfE7+sA4+hTFb/KZdwek3RSbVyf+aT0WWOSu1Fh6wHaEHGMMkHkgAu8wM
CotcMHUOCqRYE/EZ3iB7eNgrAvMgWLFvcNlc4h5TD+m7+DwVvUK5bsy9ECbBk5lIQYqh2/2maOGF
B/p7ypzKJphien9qojv7G1XJjqC1X0B1QrpnSn2L0w9ypN3FaPUiLovOJQAHwvvMFbD+UlGK6iQG
h/y32sezUjybB5dVCCNBouW1pRfFOsena3fJnpEs4XQNu4bxeqdXqNvyNQZXBQVnzdgus8pMiLuP
El5qTBm2xq5u3NhSd2XJ9i7JkJVrzu+QJKQgf9NrRbbTgVCO7u51Fo/oH20bQzP64Xwm1Cp5S7O7
wBSPo8q+nya9wc3f4BH3f5Zp5xmadxCmwFSIKHLXjvCq889r0B4iLyHiDunbHC+MRKLgteSiS8cR
IhpZDS3D2JVQ0W7f+mThuL9e+YdJ3L6cnez27VCE76GpaJtdP2H1xnSMkYUScEaeklMtn7YyRu41
1b2+WN/Y5xB6obMt9fcwSXT/lvecv6DQwE6nGQVk4OL26ulnav2K4sC4m/QXjkH3KCu/JO16k+BV
5SAi8ShGWnqD36jj94gAF4RaWy1X0o2/xlLEDSaCygAyUOtVCOYMBC+W9kzGwtTOuO4v4wGG9wqN
95PhUF3PA8NlxG5lsoEl+67Rjl+LSud1pGShdhJOY5sfQSUMV8g1gKIYYlF7Iq9eE937ElNRrpRS
Y2hirsPTmfKaXgUh95WYW9dnU2lyPWFpprFZZfi5XT/LoHiNOi2kYoFRZGMz6Z3+rz0wPT87rCT9
LZm2oGj36vUUaTxs85vEgWjh8gGARX7MsGyQ8q0wA/ZNxk0VVZSUoMUpUNY49aKs6vwtioSiuRqw
7ZqHbCzje3YRKAGA4u+Uh5TsgqeJk2jaSjSiq34lWHUV8LWb4MFvx7RtLlpzHNCLBm2tRklTW4KG
6rUsDhXf49ErY/P5Xk0Y88bdkoCa7cdNA7iuein1c0iVbPweWZ3sZKvbPzaidwoik/33jHe4ECp8
hHYXQVtEoJCmI7K5l0P5h+apMKIrzprF6shG38J/Ksl/jilzzSp/jLfiIO6fgNbmuAElT6MdDOzK
dkt4JcWmM55D2aAqlbKQ7zwMvGzYMHkSSXVaK3lg4zUZlUy8pAuw+ZchKKOs6eERkDOEJU+iLf5b
8uh9ry1O+GJN9RWc9Zn53ukpJQTZ4f2KAOoQ5OF1SVTdZLtIKtfNw7F6GRb46wCgs355RdM4PG6X
f1noA85fwCzVq/mBgSVkK1k5wpGPUSfPNBgZGyRCHDtDpRwUtYgJbaxRcDi1MtePgdFHBKAYSI2p
uX7bqkqAvZQbPWDReoZCOMPHOBR+DsbABjoQOQdBpa6vdEDiuTzbTRwY7VjOP99gHtapDmPjuBRX
HpEPt+T/ENAybD8mx7Dgp2/hRR7Eae83IPvjSmYw9Xup+p8grFXhJAIoDBPTpfT4RsziTiZQs+Cb
cIxSDMkG2H3DkqTtFqRXfqjA4JRq6c3jNzHeZfX8wtwrAu8dxgH04J/ZRjlvqhqhidhmXUlIOFcG
iizm7BTAWBvxdyEtMXEqg9WjD+AyfmxUzbNgG9P4xJhGvWRnkMIT35fH1OB+BaJxzAZDHUTOVbnz
QGgt4RIwhD9be94jADPDsKrqrwaX/0GBP1qPbAGgfihnD8n7npXIb9v1C0XEJVyFFH/9wghBa1Eu
S7BrT9D3JoArJLaVaC+7b9++JBV6I0uKiGwr8myhn4CmpzNPR7zSt0JoqBmOdLjrKdkeBS9qUcvu
sBTjVrJD0Qpvlsaug9dXAI9t5rXHBFXrCOV9p6SjBzh7MP01WVcOqpcxwQpsbgpIrWZzQEhIeNBb
8rcTVtizDK2Ude9FFnbCMLGjy35Fy/mpQLqXxn2tLMi1m9VfooCF/5jJzgr5biwyBevehSUYRcdA
iWRDk3c9z+0+1IvgYeXfentEtpxW8xMtIsrCf8B15eP7sTCA22VsWaJrrR1cbWed9Z/vc9vPztSU
y3Qfn+b+KOXiDTX0m1MLuN+V1TUzZb7bbCo+HvevgwsGjinxf4Zuk2d/ZtzcB2KEkiARSN5xUhoP
UcbjmD/HxXU1K0cEbC1aNhFds5zd+2pAJ6tUR5oP0+bK2O7f/6ZB7nlG7jepbWwxV4kZo6CvBq+b
zJHiCBCTXgIcYSpxwj+cY8ymU4ghSCNk3Q/Zdse51DIkgLL6UOwNmVayS/23wJ6G+Zpi6wAyaNvI
0E/EMFQNhaiZrVfF82k/2wlW1/HYyUGT9G1TxKoy1Jh8/xGqElxS08o9m+KyTlwRXAFJTrz8lHRu
z1bU7DYc8hP8Mv8Zee7eOv2Mp4mLbKJpf3JAD1kI397fIt4WJeK29YpZA2bRdWsSoZ3o24GzjwIP
oOcEw1/INtGt579l47hCw0/oc1WW6/Q6DjaFTJJUqQaOOaraI9t12pn2utPQX79MCEVO+y7OW7mg
tfTMSUsJxThDe9GI2OXJ45cAr2G0TZjIWvz9qbx90am7R8Rm4jhboGwLld5pnKBMpNM4R6R+puw3
dkoOX3hpSFGXw0WMgAXqP970tRwexLUhCda+jf4Wq77Urwak1RkJgpLfvc/tVUEoS/CNAwLS9Psc
0EE5kFoVW3tMArKDJD0wrCDBxxPCC2IrasYz5xKOFLaVM7q25AtuBVId5SYvTMy18Ivg/f/5dnIO
K21k6yV+Tw4Ooh70TjMI5OEY8hqiYC3bkIrbLZwgRkytaG4Ak/n6EVjBYKE6ABDSQIJcHA08cDvj
RMu13H6E/6BtAjmvTmLzGTc+b4MeqG1fdORAt3ABSwbSo/pYZR156q96Y6LYpccZlEZhOu/oziax
qetDeALojX1SfjsqTaKP/XriXYVVJjT1rNRY/Li7lh+FWulefFhiw/LeUWqE9taqnraq+elbFaRa
k6T56SeqE7qFfPuGdHcFjOccF5Le6rixhh2Iofcm2z3QKNv9NXFKri0WOvhp/Nq35PGUAmX3gNLc
ErTmuzO60dtUb9exA6i3FTyaNmDXg5vaaCJXbVhwJuUHhRPJV8Fvlfw1nAatS3A+YvTNlv9d2LvN
EHjMCEJkmapnrpGQqTd5T7qSKfeCFyAo2WUEPy89aC1qe+awyeHJBO1WZYlFUiTg6Rfda4DHOjzu
13CqKfSq6qf7PrGMwlh+BTxuYHxqZ20xHfP0NrKkPLQkBN+p7MXcJqbAktt4L3EplLh1VZZ/2BNU
x8bgL0vQWiGYz11yFshhYySn8bJVERiEWGAJYKu82X8ezH2Q6X4HdXo5UEDJPSyM6kau4MAFTcLY
MKe0xGw6jA3l9n4NA2zup2sOvl7wNcaTzG7FA50s3JJZ8WX2J7fwNgunPz/SZxKI6QY6qU/DKdyu
9RVzA/4N+X1AfwlUqWZPSQKw8lVxLUG2HL4IRTFthVgEXmhHBjV4pcmQIaKuvkUR04wVpZDSaBNe
NIqFRDX5cQqND+KuFpck3dSWzMPRVXXiN/LbvXc6Hdfpp0X//czJXYOPKuuSMdpLKJbqw7dLRuFw
KYAJUOYWq9cCB1mzsidma+k540RbdBKhXLrmoRe1HUXKV91KVynElj7MU1PTVD0PWAuamGF7sg+B
bejI8UwQf4rioSxeB9SWeMtkufJONqEEnHc6T51FPY1wQM2ZctGN1cOqvDLVzv+fynuZUrdBG6Yo
ybuWZyG5W+ZzAxVktq6kXbzbImMmxO8Nv3sDfzNLcwH2VlVeKBkRfQ2v5PHdkzzrzo012+pXpyNU
wkoPbPtJTMWrTie0r55JYopLCoQnBnFiqO7Cr4Bs8vi4lSEApRup7dPEOC0GDVIwa7cOFQBp9YKU
VXmofgMKSTfyUMbuBieqJ2SEYv7beak6FfMYDY0B4PiCWgvym0nFS8158NFVQhW2VnXiq9R9lW5/
A4JMb+BBxVYzgcSGxiascMkvOaB11OV9n2Bh6wA4OnELUy2EcP1uho9DEMQ16TXc+SfTKogO6IYv
PsU3Zkfmh6zP+Y8sBcgcVVnFAmaSMzmse3pASszhjbvUcE9FCRLmR6WhFxe3aqZ7pgPwe+msns3l
twyWaMi6MxI/WTTgdVcQhvkebzDK67ixmRVAyBPkNLxVHBu+n+aBpJAfnnp1MTcn2ImjNiM9gOWH
2eb+nX6bnFxaCtVpCYv6F33nSI5gbmwzh/3DN0QBijUwl4w88wHKG+YdCz6pYIZiBEs/qSAZYB33
VvN4Gtfkd4ho67A88xZZgEPY2ySUyPD4xbkzDGOpmMhMWZ3KS7MaAat5+mDU+FnMJd6AElObq0ve
F8idir6C4SF/psXzZl6u2IiAm3Y8YoEQFPpfQq2Txk5hzmLBHjcmdPR5q+eaNuRAxqE5QaSj1Ew+
WYYC2xpQ4Ga2k3QarS6NoJXINwDNenadCNk9AXoqT+X3hm8K0XwrnOPyJdK6DWSr+OWfdyVBL8dL
3t9Xluhz0plLtGZF/ne6yhUM/iMKAYgrM2pkekR1i1qBkhISyiiSdykZyEA//N4k7qBCxBxx2Uj9
fpG4ZGtZ6FTbePcwk8ezwecaPtZfllPcy/nEXFaSkfS2VnoElQDg5+ASxhNCiyr4pPaWjFuWzcYs
Uet01VhhIY5w+8FTYT7xeey738rWqWWhzGDC+Ut7+bbq4Qlqna6t/2J72fRXrVtgWznSC+M4Yajj
enuc+Sgv0FqbvXP5LtvPeY2iIM06lPshua2xV6KzXGxgejIkNdmSL16Pru+M9ZALQgUwuocwi+r6
9k3/yLzkWWZMuVQYw9PrNc5SMR8P4kPoh6FCd1IQOJ4NI0yLiChya2p7NWOsJu/yeX6pznq751SS
pZ8/3ked0tzOqhFGe2w8LXDxCHczLAByZ3theMAW3y/tlSssMofp1WbulooAPFbbc8rGITQjlSCq
Xma2kt2ZEJZMpfCEvJgmq8/Cawog/MwOftzALI/Eabn1FvpkBJ4iBqxJ/oYA3t0eV2xlZTsAmrDK
0+vViubpQ+rkVv6obxqL9K32jJt0msxa3PN4G1CKHsr0u0EfBtMVr04zZyyPbmgrtMHuBEdk6ERk
k0N/OVPrVfcaiZ3OT+DfXthUUHiE0G596RvHE1NAh2YfIWO8uElfQxD2zkqc27VxKK+TNKmMpDVC
K1BE3ke4hCuDk1KWS6yKDblFaO9UC/t4VYazN6kWJ+kR3oEeO/CDIUZHRFk/3gMAXwRiuxxH++fF
1EnFmJIwf7iXTdToHGcMmDlDk1gfLNK5lQrN30itY1zvwnh4z2uXZUxCIIJbHBTcxUKEVAXb8jsA
keEnArVR2RaC9uZ46lPuKqOUXOC4LxSh4KO6tC7RTho+Bz6MaSJKRYPwV4ctA++dcpEm4XdXRdr0
BR+t2CKS+E2SMWR6UEycvb+xfFJaTl3ujCkC2wGlVQbXl54PNX3whb4IxW7dBpkn9clAVj6QX8hK
CBCr0ngCda8Z4Y0whlOaeuc/8g0XUiX54M2yiyGlW+J4CMxZS8cTreG4sK9xZWO1WcFAVWk5iHUj
OxTla4TLGRbY9nDWSLnkmwwSej9Hjlp8qaKpaStzLz0gFtsMNfHOx6bfxNikicL3kpxQBk6uVSkJ
S45uzXzqIZsbHSlObD9JbogKYf9FWcZ7jSAEECaPMG+5xNNjJp6lwaeV+JYjiVrcxU72SO6ZPlJX
XPB/bycvUrnCvanqQXb6B6wOZJ3Ywi1zQ5pjImKRDqoPgrwRvHwJyLEX5NWaNBQXokKQiaoMcazr
0XtNq+18mQAU6e95+XAXjPmT9YQLhK5H7q2JjwE8s3jBINNK7NHorhJinYRgUwXghhPAuxg4eIWE
flhs7vrPp8HoHiCdD07aKAiLh45GvrrTi0ag06XrE27Ygyg1hTYOstnEECJpC7pRmck8fSVaHRMT
tdhalFA9ww2Vk1NSOhZcAEs7zAEFVef1EczgHvWynHfzksDSsPUkEUBz3fZsiP+2jgvHc2/hvy0y
YGIOrF2QXf5Y1+L9kmz7lYxlhCHa6dmhQEmwAaikSr5zPlWVp1g+vKG4tfiLaifYrSJyC2TAGBpu
JnmcsIt+aph6TFHsM02+V5vsple79I5NOwDWlTyhnQQGCD2T8yVWMGoPRwWanQj4AWeTA+XGB/tR
G2qQecHSeXT46V7WPScHCuF+3SjQYMozCmpwBtE4UpHKm7mePLPV78Lh4ru7El8BKJqcTORQ/UbE
Yyu66TaJSX3OrIpf0Clj2kKrWQ26gr6JaLPrEgt17Mv5ymWA7+uGq/a+mSRtlUnNcWcu7o7F1Wq+
Y/9basyl7O70wnIMouHzin3cXdt7Ns0GhUBhVygDocuIE37CzCtu8vc9F68IHmROzjtVT9f151BW
p7CU/slRq8eU7PHmiZESu0DYJfS2bZSuxmBYOT5ngPfY1BZNrVrLuzzIlF9gEvn9XS0Sg50pEqFV
eBSzerkE4caxE2h0ZwKrs0rYTuqDnQCyGf9trNSMMldaguQ0TAWuP3VeUMkK9eJDzH/b/YDJFP8I
JMoBFhmopH5dBJhYX/EVC8jWogJYn+4EmzSQq/5eboa7WlYD7HorgwcDN5K2erZ6Uhdzcnq98V6j
5PcezTcyluj2K1KTkDRGrqXp1/lcMDzc3hRa6qShTdAnRAlObdoeK2kMKkupipWpPB53XsjHCp/F
PWgbF1DKcSn+8HuTwixgzT0j+r6Wd3gqlCWpTXcm4KMZxYM8cNKFqN5rt7qllpxYRACo90SuNCQ4
GXTTJw4zWhqNkODLUGFSDzNxEtqEWVlN/a6LfkAWC1kCMR3gbJaxzjGB0FjUyBPIltPKomixJXrv
DBl5hVDpU02rtIZGNeKIBgS9R4d1+PXLG+x3or3wlUoKSzO5o5vZfNOyPc4tXNUkHqKjzIAorOxP
xfPtw5l7SV2nf+q7venAH4G2nwy7ledVGfalO4e/Q8cdUWV4LQJ+6uSsRUIJHhUiliw9xbw7+nEu
mxi0w0bit5bIQHyg16QGHnMNdic6o1Eug8Pd0VMAvHe8gGswHh4A4usunCvWAHobmtWOJuEr4h8e
hrexgyMBEVhRTb6uEUko001swR9FH6axE97FO+8NatYTUK7zrIeOeufBxg+0WwUk/6LELj6jvc/x
Z5susySMPVXrNwZ03D7w+QPN339ZkSgxXpoWu7GUHvgqp6RLBNmG8KLk5Su62zV6Ybx4z2f7ML9V
5tW6ALlpuCktpPDnpPziLe3tgz2J9Wrt4PTXxtsnSe7PLgVXvHTR5ozOhK+6AsaYO7XlVIhnByXa
QlnUKDjhcuOns6pXZ8++7lZ/95UOwh0yieFcF0tTE8CIL+e4sZieY18TsmoHtHLfFKA+whiNC+dR
PhAORtY/ZZA9cKhbIZuFPDTq6lOmMeFEqZ/YA42p7D3GU8dnaBbE0gn2ATzzCXcYrd1067cJU7Qk
0Nfv0HrFHWwSmpbOsonBwdEtjXWUPi2+J5e73UqQkvE1Qnq9+zditmHTSoS6h+VTQezPZCoicqvP
EeXMIa+9czTeJZu13eReTu+XkEo2EFVdYCvl/D1nlJAf+MCo9vfX/yME6zTULv55Z4QTE2BPuidn
pk9innDQtfIxf4CnCuFkhixldJy1pq3GS2nu6AvxjWvLNClpRTlj7PJbY3XcCdSLA10K0RxmLm24
ncrHiPqIVb1FG5dc08svNrQneVB99zRlrjT+2Foj6NJeyxYMkBYzTMrVPFB3if35YshbSC5HbomD
SVF3k9xZYb+pdq8CbX5KeatygQ5UcUp/baon3QmUK2xp0H2cZCkuRK/YYrH2huFiSZj/Q7E5m4ug
VaaY89Ksd2UkxxKEGTlFyUIIBR1pGf+RgvOJGyeEuICm5Ti2nsrodD2qVsoKgeh1fd8pC4Y2wSUA
Mu2PadpxjD32yj82+wuOIId12BfrPyv8Ffj7EUcXDfaMztlFEJSYDRLQsaGQrR6FYvFip80YQFwN
F85xt5PHJ05dMd06HIvb2zg/4QYz/W4fx5lxpnSq+RUEfPyKUfM+TX+f0hUD99grSkSi9seQPL43
EJrhAu26TgwrEVsNFdXF7gltC92vem1wArE6CwVe4V38oe61ZNfrAALfueqnivVecyZ4Ni+ay/B/
qDf9oPeb2hw1V077bmQUViWI4ecwhXrKjJyAoaVzuj16p1WHpioqyyrFycS0H+OaclNi7h2fTnCH
1G5kHyxi4Z/JqsMvfJBKp8ZMzD7g+pYRhsD6PhTzkvM2x6pueH4cJ8tOr2uM8W77FBQv7VWTYPTf
rwZ1mfCvHZMZMgb3Ox/b4rEn5ru8InRD9f97MwyQBV9gSo0snImFlgaWYegNX/yojVq8jBE2pJnr
ohumlRcx7E1DWsOzh02Oqw7WdoevdfILn+66nGYAmjucNbKrXeNf4VwUoZuIrZ77LFCIzVdmMhUS
Bgopug5o4KDESbIgtq/9GdkgQ8M1colVNVHk81Zn/abAkx79CLv2GMagnYZutuT0O93+aVDu6BZi
3UEONaAeeMhQwlmfjGmvLoHckDlbSbZuY/3+2wTznHj1jqRbQaId4GQgFglD7dNIHXuBXETyYkH8
xUNTNsdwfCmEh+yv4SzqGujl9eHcTGG9c/O0h5hSr2OfAmjCqq0CeDOSi3vNxbIGAfyqDXuHeuuA
Z29Vtk2lceVs6C20xPfMEqQ+JWu4s+A/chlqfDvLCohswWlZJnHse5O+jUyg76G9DAvMIFG85cya
SN0H89zq4eNSS3gGDRt3kcD/advoIgwsjdCHzr+Wgvdu97CUEnMzxxggHtp+FsDjRa2eP8VY+HMg
ppEhr1zsIpPHhk5YBXrOw7xD1xOzRyHYoF9niICuvJeEZ1Y7lzG1VnucA115pfJt6zYnEVLGJw6e
TuMyV+ZklJrIkWsgehqVIfD/LaIudu0wLhXj+mkVO+r1JBiPpbefYu9WkytUG/Q35KprGDSy7/jM
n5JUTvaXmTH+CleJLR+caUNBZ3RaYGlCaUCFHFS/LbNTlZt0wOGnCIdeUJTFU7Y2yufNRxUIVDHE
wlO9BrXaRgunGSThOwPBKbPSZxzKEv5apAVly7wnG+wffOwi7d8ptvEniBC1MsP7Z9iS4CTrcFh1
IBLtCx2l/A7/qGn0TNacemnwRBUn/JnxixrvOtaOIcyB/Dd9ZjQRBaz/w41GoRWtgavZr23d83ei
BJQ151ga+SP+X1+xdGLfIc8e1tjjOdhhHvHkNtp3/YHcwAxgxu/fHdV2KnzYWPMHU8XHPVRGr7+U
LXJJqRc6xEd8T4RJgJk/WNTK+fhpXcGj1QE0tHlKT1M2+UBgAL19jNaUVfGFGgFx85ZSIdsLlr7U
raGNlNf6lunysAV29rVhn7cM5sVdp4MGkZgsqZvNmoGChg1i0ioeWDssFdMJ08Bm57LiB0FoTQgj
YznqiBIIr21/fROS8Qbbc7DLXQ+oRqXYUMhLwArWiQymUDVwyOV9XdSu0k+7UR0nMVYBxJiysvlR
6+1JkY4j19W+jScqj39FSmzHg5PPRIEb6ezacxFGdHZ4/cbXWa0xB2s3v+Z9c2i1VjBOzJQ41e24
jwfaxQoUAOr7CS6dqMjx4aB17L5WX1ltnDe+fYtoJeWWmVNexWFPRD3tyDBL1xS1HD0FBM05koTg
u5eOaGBxf5vvAlaBuL7fYokN1aq+cW1tpqjDAQfp7v4EOGl11k4VEmRhzYTvStvYhj8vGMQaGNLZ
fFBHa2Q2dD1kldwzAQ413SUQH4bDMdcniwjN7VDgOUcTxY3WdKgbfkJ4oa5FV8nbUiPizlMBn7Lc
rr1BJ/coAwBn2136w3qTgwjy02snsY/Mmwu91BBqxXzQLXb3pqZ/u0agl5l4PYV74qI64Y4CwNvd
d+51kTt8MyMUZ/h2AmhaFm2YvGsYmjEH7dP5lzuEjYNxlkkI30tjaX8adayivzqXx12Op5CB5L8/
TSvG8swdAP5wxZBssKYVb72k4jS1WBvHoari1VKpjKHwH7lj4By454hh3ue85UwZ/7t57KvS1I2/
m1tfpV8gx/6kKy+kvuAGUzHDb3mUobDGXRFFDl2XiuW/8hta7P9Dj2Rnb3ToL7eFJiKTilX8dudD
OlacCSRZFXUCs6fCOH398bZfkWF6Y3qdR56K1OZbHHfAVLFX+Pi24h0604BwkoD19KQ45ozq8sSc
XQHkN+UP/jBrt0gs5dZxXLLrkJKoAxaImoyfwUq+zBhCGgKfbkVxKnxd2jwOL/lAeWa7+xNs2A7u
hhMKLys9OK1mdPiuPb3LVoJ4jw5T1jh3LkCoYG7ymiLrCHcqjBYH7OcHkRXkDDGIldzuO02yW0xN
KZ/i6hSwx4Hx3hvyrOeZWhP3c3p0HLg5dkt3j0QlqVQnJpQkdhEFMgmfMBuTOd8oOzVHVMN+WeyZ
BowIcljy/o1ZLW0NpABtxq6lPH8UmtG2OljB2mLZ69Kb4AmmAF1sCkaK9Vi9DHDASnuYqBJIVu//
w0ohIv7jsfbz9HKE+MqLMyUaTCZhqzr/kzIK/4kqpB6ZpLso8wV9vQBV8J/je/g9Il0vbXa7hVOb
miWOlsX3JGV+b+XhnwDOfn9qHB9uD8Lz54IykHA1n3nBe7jA4FChe0QIuiGy4i34HM94IK3NO1v5
B3IVat7+GFYrPPDO6X+WN686rnJ6cIYDuajlJXY6FPz85NFYcZH5YO+va3AfitgBP6u9w5USaulr
excS/TZUGRy0W3J6sLbVfuUwSaIRH9FCPxPy+rv6cH2tpWnxZxsfZr8FpSFVv08IbSejdmtT4ZhZ
ig5qXEAxcJoqbtEgqMum3LNIBG4H9XbAyK+4Z8aVvZQ8uMyW51fKy+gcv5wu8FUn7bhVhBe9qIVf
+IP9dY8COjQdArgJJJr1TVSuwnbUGw+ALCwYWi3Qns5VYmBCHh/PK9m/0qlSaEHzxu0HKr90ZGlx
rJ5HFq6DmI3xgmorMWgAabM2BJADKDkz/F6q0c54cWh4lhas7jdk8wgd8EOQ88RVlnAkutssocmQ
9THnQdPDNJlSJGuKtFbbrMl3bOSWTVAIyySLO13PPkoVvAdsMa9fsVWnquhNLMG2uJxhWgsDaVqx
YZQSk4q5Qt2Pc5yy/TINpLTZ6CfIqo8vSUjThEYLJwxX8rN5hh/12ANen2btvhdDTr7ymZ18C+7G
iCt0uqS0XD9onz53HrLmJdJx3WzXrIniVl9PC5hBrfFGt9mjexx1Eemzhu3wye+C8Yub0dob/0pc
FilESHJYEe2sB8xx3wrqrnxkOx8aJB782nDZEcz74vyKy1FY1iPucJBOGFuaJUyN4KX08cjXjhrq
uTPvKQR7m9vXm+ojgnSq7T2Gn05SjF/HMXsyKUb2gqsXb7DXasndTWCXD2ZvZf5EDk3AQg2E6PMo
Z8U6wqQ6NY8RuFOXtDfulqhPN62mdRfXnlt/+eNPUcxbXTR9aul04VMC/oUTua+RTyQFYFmPE594
MUz+sa+X6hDsxRFUVNoN/vCf4f3wQCx5AzrkPkp2IfPcMNTMXPpNtXoMzFFn+/VyBmhxL6CF3I1/
/VyzF8jjvIx0VCW1rhS+vzxCrJ6tURLx5j/JdS5h/tfztRoPKVvmYD2HwWJLPPcUN9P9PC7mi8/6
R7f3616FQKhREwMKV+lXZbNXb7eoYm/VAD6Ax5wFltLqHUg2cKndvDbcSRH1kbHAymSZpjWVXFWO
15gCobTwgidPVpB0gmGLykB7nrY0Tk1K17ZmrBIuzpNw2kzaTSam/0aynR5DLk7+WX8j6OUEhBrK
/mqGTHRa5Dm16zrGiXVh9D8qFBLp+ii6CXIgH4ZYN4DfdgoWDxV6Zn2yDdJFWjnOfoR4up32qfZW
3uFzgk/1hTtfOTsKE9fiK7saGslxzERX6V+IxSgryLBYIWEIeYOEPHqF9tLWrwpdzdxG6YKLuXQX
VIASXJnJEdQd+UNxDbHyKfQHMSsuyoEzzxroO9whjdqZ2ue1tm02DSouIplyvnb59jPPwd6pxo8v
+l0gMBsNhNTTx7YzpOTcjWJm5U1bmWVmFK8pC6ET1+sUtG7X6tBZcVEtlBpCtTsuOVjFWgCsqDcS
giMVNGN/KYvlr/wEiVXQD+U/fpNWkU7oDyWMeJVHoUFzDesmcvTlPuAZYxb29xNpnQFRmjdbvSsJ
bhRCgLyHxHrq+IfzTZQXxG0egaYAsyLmK0MwOyIEIfiRvr9a1e+58dpjT7B16iqosWdGBYs1Hzyd
yIux1sOba++3hRo1A4M4FGocXnOOLWT+slI1GFQBT/szuvKgtjv/fDwzeTYV8+0tD+fDcXVwO4kI
PWREk0cB3uIgpxtSzjB8dgppwjkWpVdNLVH+pzh7ljXFxIDMwHWle96Q6YQ9ARVVj/Csj451KM7h
fXGNx/dW6w4jq//+AiDNLhp6sWJM0k60A4DoR89MXbeiEQQpUwH9E5zGNMK/4K5JDllH5ZMDeMZV
mGQdulJC/ogeqbSI7JAzHPR6dijHmSMOItGki8rA81aaSnJ3G82LMDKzbzZh+dqcdmV1wUPJZfuh
1Ydp6MRvb6l0TMemo8pAyBP8ZXX0lHiobT28uAAg+cIIyjpHrhrCDKi5RM02oEvMpEBkSe6Nu3ol
YWBrvH97BbBQ+VEehMzz30DSRkxpxN9Fbtx0Y+OZotGiIxauElb5dr9u7162iogQDGgeIKDUBSWh
bq7w82cd0bc0jxMAZkNO/Q5dAEiWekyzQ/XuFGxiMr8A8MpwNiZxtF4MrmIW3WgvqRb/Tf5RQv27
l6fUIpESqZ5aZ2+9ooQnPnEBN+eaaT6nJVhXW9SijAu/4djJ+Y8gWpDJpQldM3xsLVar5lrNYuVs
h+I/biFIBLgT/OhA5K9BloCoYC5RijBPXZ7cYWEQdQfJsV5Al6hsiM80UKcE+V49eajmQPAK9tMj
ClFMLsGm2fGbfdSmnzzt9YdrT89r9UBRQnX4nf0Ca6+m4pECCDfiioDrBgWVvpuLIkfdL4YLOHXM
+vjxW19oPGvNOSvRv0gwYZ98M+hqpo0zM2eVMKltVK24sLayuYAweuHBE02Lhhl3bS9VGFSXaNeM
mj33nR7UxWx9hFF8f3kSzCZvbC5Zr7BpQkMU3cXqKOyYdgPyOAnFia3NA2r3qJsGSdn1GuhU2LPV
9WJ04+/BPvcut36CAn8Zxl4TFnm45/ZPdH9it987MN25tEbDBJCDzNjt748jDR6mIbe4jDojAjSQ
td7DiyTYx9UTzG0DKCA10BbSxvBNWWh5ElNBV7sHyB9Gw27iSfVdq4QrS21x/wQ8NWp4cG7pK5dO
uQL9/MZ/8QfmidZOUTwD3FLY76d1UzJSoOgSoKSokrjV3/6oMNoocQeHyhb3diYvaY6s1ZBVaHZM
ca4UzWiImVZ70V50hr7IPMTiqzRZjiwFuRoGuTTy+DfpYZ/5uRrU+MdljnfzZ0VoqbYo9Ub04sDs
ye4Ipxdzrcz+H1HECNfrY+p1c+KD3/AGPBZKHqPB7DfHHhHu917qBhCeqF2kXRphrDKzfTkaCjsY
ybrk0vXVDmLXjhfLxoN/Sz19axPbyUAn431UfhfP9tjIQ3XZpXeL1evGwBlXYNuec3Z7qR7oO4PR
lCCxeIdDCg2WWaJ7WCvA3WZvszBk0xPSpmw7RBzA4nJwMjQ0mpwU9PL54UfTm1OML2mboirhxdVz
3I/Str8KAbdpC/Uu8aISarzS+P7rggq22grlhkwOuJi3iTF3czUDIyKJI/uYRdYC7GkR7IRsvubj
1+3ObAXgYBa4ul0hAVlI7s1JwyVcr5dxawJoajRIkulAl9mb8bVhvh9wjWU80mb6rVooEDVt4eI4
NB5AvzGnH8S6xB87fF8MQfhKHDYO11YJ5cfcFary5ll/zQVKdPf81r1LV9DOsKL5IwjDqhKOBKuh
IdquRcsUT10ux80BsJsFt8f3NhGxyIMTDOAB1oHXo61BqyE7MXh2i7nSblBHTRnFa8R9DZbi77Nd
6E07c+amJh7pnaeblRt+tqrRHjgr5aKm2y0t9N7m881FKXvg/p94igMB1AjIlZl6jhWAzRkYVj5E
quen08LlXbtHdA3zkQUiVH5hPtsNujevhB+7cdesKCuBphzdZMoVp5jbtUt1BpTSi9070RJWrIHp
ecL49GwP9BAcw6mmNqmk+pX+lbvnVvrIQxhEIV4fClbTQwVnXFhy4vxP04tysgJiPUIA7qsYHh3a
kTWw91LQrUGuflfAGwUkSUKifRQgaISoHcnsBZoXykgt8OU95ymAoDFzXwVbVyicZSYaupagOzBr
eJQwqchEekKeLOPwwR0staE2wFjqpGAhU+HsBaCR5UXcBHlnXKFXW8U6k4qid+8AeQhZGeRP5OTv
oFedJLFQsaaxLcejD4lzwNNLRdcmWxNLersU2WW9Xp1jQn4bqqUg27f5R4HYm4jKOfPdZ/9EsPUN
ladiLhEgPjFMEa3gVpJXvTmJqPFKdIVI1+rk9cPlemrtBRRPooxMEXXq+07DqtueC38HcjC2Lg92
bU55oPwZAwB0Im0d/1qrkkHPyCOCMmi1ZJppptbafb/cUxH7gu3cVOgiyemqqBTxry4f80v6OhCc
N11AReUaNwaDqRdTe1EWs5kSvDFb2dM4TGZihNY4s1o81alEDA++b4rIyl2zV9ZPQrlFB+/66LIt
LmUtl4sdchdPlN4aPbVkuwioeSu5hPQz28Sh5V4pfOtzYu1fmkhNJW4jvUIG+TPydRB28RkzJD9z
7vkMCkHjjExL9lgEoFF1TRdrmRu2nWdMnokxmAeuyXIlS/PcjvhzNepzYdoFn0Uaus56+YieRdYj
N2qacm35FLu6hHsZ1nDDsqRIG3AY90ry1nJk5fePAtE0I2dZ6Knyj8f3MvYiDJgUyRhiRusTgbUA
IboR8Bh/Dyc8jfUMBHB/3IjognpIUPfc6NDAXD69SR5NrfmBSkHlE7B2XzlpdeHiTP/KYoT6EUKp
lipx2V1/L21uaDBEacLxVsUr64G+DWI9aPEDK+5Uwk4RiWhEhgRT5RFH7XHLJicv0JyDdRe9NvVs
EnJGdDiNCMpptCZFOvv42j7PzhIIFTr3BcPerqN6UVytyPdC5oLq60RZwB9CEwVrRM230PyUr9GL
X0p/Painc+CyTAH+SRKLe/MinK/V5i/uCVc5uOe+G4fq/f/loylaM5fCA2XaTAboCdHXT2wcRBPv
tF7MPjHLw9XxuN6LoIpX2bEapSkHL5TrMO4kIRxB3jGVAGFMvIe3Wd0j+ngpTh6Ep9FJ/3l5xyVm
ptkxlf6V0rPPEvgsiFbU78avlH6JWMVJBeEtBTeoemPSxe2VQshO4oMwaUxtjLy5TZJ7vDYcOt4L
1CSbFaco6CFBTE3DIkOjM4poQYGxlJdatsiU1X7dyjPXE4fz1HNCTC9jjTfK8H5Zt4E1aC6A6v0+
oaqMQuewDDzjWkHUXt2a9Sgkktp2BiZ6X7DOfqsujfp1AZMOAhsdWkQ0r/9pBPVUanJnk9/4DQjq
oAR4UsgNtg+eO95og+CeqabivJzdE5HHMHfanC9xBxkryz8zvUtOb8TdZZWiH2ezCMmlonS86goQ
FK20bz2danWBjTotwxOicksR5CKa+6csXd5NP38plusrzphGMX/VEjWhLJ48zxRuAXiwC09E0+fB
VPAjqLLtqBKTrdA0kwE+8+hBt0dX1Ak6+KLqC5Lejx8xxF22ETEsZbhlJmiePuMO/TMBExXhqNlL
frMc/PYSVUGtLr/EiaX6L0rvewbiqYo0gV2tl/9nd/IgZ5vpahO09yC2v/GeZn0RG2KUKJ04Brb6
OE2EgzfKE31ETNTvPCE7gjTBWpOMSToL4MtPJQBJLaimYNRno/h+ByvcmcQrcvQeHQNhbmJBR71x
B8AB5sLPkzEKNG3OJmIGvUwnsBPLgPjbjLyZPqeqZA6VbRkC861iAfK8CUMJE/o5fKgXNkcRdoG7
ukfFhywELT7DTipHVIrN5uslnFPmnb/8uI2oPEbY03GRL9vq5eRtCKvKltqFO2D6luGZjHruNbR2
560TGAcFqLfrQfD0co4EuuS2qLLkR01lthIVX9tieGi8vLmT7P/ri6epfZCqFIB0pgczoL5pqg5j
tSXupsFvE2rxO8WiCvF0aD7nYPrE73qURD03j/4RGoPPiPxv06RtFptYkz87BVbnl/+2QRa+fuFC
M0VXVGSZ7diO0NErcjTAu3LcOfSNuUnHCoKPLCTBu2Ra2vNGRHvQYz2DRnZYdADjb4DahIdNbhMw
CzGCZujHGYyombNd5naHGiuoNbX9Mg+icS5KfRDOiVXr4HtsI4M6L8YLWPXJGsFqQdNENB3JA+kl
XVP8tV/+kG/coZucfE+qdOne5suCOjdk4FsdxS1dQuW1pvX4ySJow/IFZIEpgktoCCeGEXZwSliC
UY4RBIHpU7v9viWU0V3GJfD0J7DdV4hKgpSsxOtFM42Qgob6P9ypYGvzLoyi0/5C6WzqbZ3wBVFU
PuAFsH18dovXUP1AW8KU/ygUR+VX6z9S4ksI6M5ye4U3ee5XetpeMXnMcTOQbDdDfWj94xAmCbTp
lwmYFDLipsBMnW5z+4OZnBNvyY/bDaoxyKSx/W4eo8tlnJLNruaHbmzps1bWdQ6sE37oel1TN1w9
cQbJ7gOd0/50VhY0v2NpmUUPPM3TzGknt4SGAWggeKBgVIWW6LamMexYSow5YvyZL29gOwJ0VTSN
Gx4dfznqKDBCcFGeNLhvOdiBa7+QaYngRax1sHhEldYeGYUhTBya1Gs9PzlRLzBLVLF1Jpy3mMPZ
0xdK7k3lmffPXWAmrS7daKOH2YICmNr1aWTo3YAs+j4A+3rVFZLsDEkFsk7vhzZnDnX8+7VMgn+2
IhVMkfA/KLIHJDLcmessq2SGEcgiHoemEB6fnoQZCGHjquX9GVqvl1IQ++s6OZbNgN5RPIkPd+3q
iWoeW0Nf3Y2r0XwJRAfTm5qR4xWHks4M2LN4dYgDMZm2+vgfWVThUSB2sp0nz1263/c1aEvqWXjN
hU4pueF30EQv1jf50uqaeSkFk6FVd66qeTYn1tiHnui1wr8f1dHuBK953kW/JibRM0dmzsN3HELo
P3FT2eUPOPfHZMl6pZfuklsS98s/kKdJLXZjTonOTC+CJZ8XqYuL4iNY2ZT+rjoCqDJQ6FcfB6N2
mfqxVyn1jqm61lH8/tQFHNBVOyFtcCoRi7pF8zqQB2nJjVlySNurt/PzSAzWWcBFSGbT7fMj6lUY
bEtsLw2qaOUKgrtoyiTBbDJwAj6xdxVMgd1mmDelqk0pWpdN3v5xLDocXYSkjy86W1qUmu01Kuxq
fERr3yku+Kl0lLSR1wSEaqU0qoPxEnT7iRA/e4To6tfHQDI+aBSpAdtLB56WJ975FtDh3igXBA/n
3EUkZU5WHKmTA4Q9gjinaVD7JgnIJQjsKmcqE01w8VWZBeEyfcEiAhzT4L5qvY/TeVD7lEWrnKIp
sczCiOWbuSo8hNushqKbhUrcud58iAXvsug8Ih+sq40r8MHjDWnT7o7Y4ldv7Zvm44PI0FwG4+JN
7nV2kNbubH7USdod95XWdTrnGaZR+vT4uCGhr+Qlmf6KCiMJNnvTi0z8YafHGY5QQfCkcT/UKEKX
2ol5bbqru4rPzd4b4hsnURpBkieSxDdc2DeE1pPumNZF4v3oOqWLBmJ2idX59Tw1vw399DBPLJHV
+AhVrgRynZ8uitLHib2UY486OfOU1xvnfaYec4itfgRrHMgOSL4roYiISLzAAuWqAykqRt4TyOtK
sL8pCAsUh9lJU0SDCoeKZ8YVNNHz7ucvFo3jqiKuUyRBNdlA97e5SJITamfPL3TE6VfjwLQ/X0/I
5o6QTQdxZES6lxW0Zf4uqrlV2qo0rkDTusrk5heRr82pXgYGnFGmRo07upp/BtA1xI1eKtKGUiur
GBT0BfRh8GfoXTE0VY2nE12x4oySMBFAwTJ2fkqYOpKZ/KRj0OBNS7ZIYBUlQrFwcclKY8jIlfUw
OzTGnOZOX2oBbl32MkuJLNrbN/gOZqolIHb6s8GnAFwXL3Og3yNyvpXBwnM4Me1Hs40rFJ7CNY2j
UhCIvUtQY2ct7QlxVHq4fMT4r2Dip52xmgMhHTaXDhgFhIM7Fcw5PsQZTjkcSZZeOTDVUMo7sbK5
YS12M5+vO3eT2MBCqP0texgZo7ow5QGZEhlK8UiZGuNJ86MhUmg70PAb2JspHJcmBUSarsJPID6R
1Cj3ng5vpfpJjPz4hsS+MYUg5PIrLetr4ziiH/Yeu5HufJiRCWuXbQk0r4kp7ArxONMYFPkBfmO4
LcaONZcfNyk2PgGHxZCU5rTu3rjx9oC2hAB771mCWplkZ6Sk1x/GHXdyiTXf8zrMA/+2k55ZJJfK
rXk1c08OM2t7k2FgB8rAXJz8Das6Khlw/7BoIQ7AWbGtkMCiI66hnu2OjlC1NsiI1FspJyhfiF0X
L1nCAznbBMBZbb7htXaPUWwF04Kg0KYvNo1KSUFRGZROoVr5jPpM1pZL92DIG++pkzd/Ao9uCfJq
cU/HJuwfKfFgmBoweV+UsbhmD6KxSo8/3m3xv6DAReqmeqKZrFSsFlTKz/4h5eEPs9rZnmWjSNKK
So4vYEkkBgfHEaSuZNsETNfTtgEFA9mQeVJAdDmKp15WCtkC+KiRqKspyhU5SXBx83TuhTS7ASJI
bi1zzYPA2ARfvE5vFKpeXvjjLFNxXwyyHXCX+FM3Z62tWtVHaE2s1iHst4LyxPQ4YtB05qMK1cYV
I2QHS7ngoesMpXkXvEPzhw6aW2BWwsegA00r6AGUeXxSXn3ZoA6F+xoEhAkzwnQZPLvgHB2kO9it
m7c3RZS6yPlkArXPInbOI/3eKTerinh7suqBWs8yHP4/FCQM/HWo2J8nIaKLy88/vpKlU9jFcYC2
lStIMPQUhG3ftV2fONF0YtNCAi7nNV+QV2StOVNAO3gd+mWA6Aatv728SY/vE7huyLcHP87lm+pl
yJQgCfUoL7Qel2jWMI7EoUQ2HMEndpJ3Z1WjWPNaLxk1C0wqauy/qTkEldaN3y5H+WnCPPpg701v
h3r9IAExCIrwWssu5ZUDrYzODpKzQYeEkonCNPXCY5upg/2pg3CIMT8GIpEfWLvncYJfdtY576o6
q3riHkVjR7owaz8hWG3EwyJPloYZcRQonAQ1TDWRC2b0GxLX1pPfA8fpNF9q2zdOlbGc/lE6wjlF
VkwTMlbsyaHJYr+ezDd3y8i0HSOAhL8wpHRrZZQaTObGEdHYiLmn0XA/bcqicGaYsNBCyMJoBwcv
12DDOnwBIiS9Ocmmp3mExu4HS2kMFsg0fNU8/v2WXysjpIfmxfAvmLYcbTIojQK+DK95A+yf0YCE
7UWoSgaWnUUmzk0BCegULZkx3ELYGerI03dSySbaHrOK02R2GrQeEUZOWrR66/1STiuRGoLudfCW
0yeJCz4p6+uFApHyMdLGrViMoMIg3jBth6ZedXjNicNX+H89AUkbVfq3VMRXDYvStJAAqtYRZstc
lyDKpABWD2AFkMXBATVKCRz8mah6VPBPd5oqdb9gKr/r9IOYWt/GvY5Ma20eyplx9GYov40N2/bT
lT7wsjHqLMB7g69SoONQRitDSHzctE781tmiHbGi/JURne0gD8+HnP6lw8bBvgjAvCKrj4TF/KsJ
YvvwCBJNcEI3vBoJbUOivjx3mGTEYiB43aZH3PK7Eq32nqi+x8nag/sWdiQBSgbPjo16GWk2RqOH
rFBkS4OTJpy5P5ewPInZdl0qvs8cAyRS24j1ZPARaMB1mnR3CO1+i9FI4lBLU3JWmvTJ+SfTFuwp
UaB5qSXAfuYYLs9Pl/BD1KV1G1KLkDz8EzHZTAF45R0iMC1RN9AIcsQVFz/opi3kkyrIR16xFjeV
2G/Z1sYy3TM31IGY1/OBgAWWzqZO9BezqElLBETBFBaaniEtr6LUMOsrJ3+kmLYmdOI6Nlqh+hZ3
8qwt16Z/5iGojRN2SMH7vqMGeWjwINnO4GNt/jys6HNdnG7/P7l1O9/+wGlK6f/uwQkCsVsSUvS+
+TchxpqUg+5BupjhUw6gg8uCixhc/DgEGv5WaVRIuymQlUyYQrhAr1edm6iQPJCWsyvM/VurBQOz
GZOs5MLbNrAX9LrQx0s5TOoPdpzL2qgdP2jmWlAnZ6VcPIl5gQwCMyQ5O31s9gAWieM7uI/1NmfM
IW939kp3I7tY9saBDWgwWbs7mLjbREeMbpNTGEJgCmRszXwH/u/QWug8Ivlj7gdpEXi48bFX2sHD
dW+353mWKUoeo9k0kH+oaK5pmk/aPKDyvEJYhUeltCUZMJaQ+sQ5BkKCKm8PjxvnMeqv5BENgqfA
sY6RF4Sf7cqLFy15xLLYUFny2D1cLdjRrSDz/PqocMoppjIEIvt9BAFCjc1rDRBcCigXbiPzF9FH
M4yDPyagnGknqsJ9i7SXC3lGx0T4mrwwsuuqCS0hZj4SLLLnY5B5ZynImo+Pal0/xtLpjjUBXotC
WCMTdZCAFcCdefPwUvOkbint7Buxrs5d/wTU4PKM7Aq9RFEQwMIlGPKyJpmrDm/DvKvzxyawu0Il
LwqXVg749033XG4RN47voUhFaOJU2t4RCCsyeVRqdW2A1TKqUiX11NnXo48cS2iWVTxnzAp32+i2
HM7n7dXpvoF1OKC7viktj2AVtDX8K4PWQpgCo/Q773fRm0VWN+2hl4Rc7OaU7TMcuRSg3EyFGa+2
QkToX6lEz6CYm4SImOteZY9H0kkid0oU1XVdxJj1wWo5S6DYMChSZ24WT/vrKIyHXgm9xqFL11XV
k9mTkNY4vlOlBQAS+aOgqYRSylxxNb+bthh7l0b7o8TIYobrbs2IKalhXoANQTOT0wS+UjGQACHH
TIoNnDTU+Dt9XL3YA3z3fZUdjQM0RMVkZSJF1MrO/pVOcsVYC1+2ZdltsgotjvytuVofd+xeN03n
BEt1qvu/0zlicqPw62k09wKu+ZppoJ0ulM6WIzuXbtksHnl8BhtoXh5sB6jCG77iEAoqtlQ6S5/3
6DkQ9sPQCHczxCizsqPoXjstel0K47yMr6QVskF8rz7lYtKlCYOIL4cJ3vQrfpUitZAJpyWSmrLw
TsHZR733DpDN1Qn/5f9cxB86SqCxLDzOB7dC20odHsM5fBNLzhDj4VegQlvVOYdTvxKm5rE331Ic
1vxFsnpUsyYJRdF1QZ+Cp6CzHsmxJoB0t81WDe2t+R2HU9j0MJrJYZXqJOFvezoziooUIYcAhnWe
2lHsDCI2y8oGFhVOZF/73jBL1Qk8eg2mp6EXdUl6S4330aM8gMYL6URPyaPGuqzuUTlZPH8gB3L0
dnotO08gQnNSdV79hK0UnwnhdlH8jPRpnuvJgsmbdO+hPdac4611Y3ohXqT/o/ruOh+oqPNY/+H2
MsSKka9+WBqxt/14iAbWCsrpgAN3fY9T0yTwwTgijU30KoSn2XVOdE/ZZTxVessRISpxohTt53bn
Dvx3pFtHNYzr8M0mstvEu11NCppIuaniduAtgO6hnxMxKEFBvZFIsTzRg3MhM+xGpjc/wFcRPqlH
XZn6VHjUymxR8y2K5E4PCMXsuiGhatpJtV04oLWlqhjvPotHDPY8TPpg5LHaZIeqWQApKF1mdP+F
N3jaVJK8QrOfK4K+XNBB/p9HxlBNNVbaxCsVDUOguGOmZg8NNnAZ8ehNFgvS6eIuqWlO5XIpx4cV
iL0m/8TrstmYgpEAhW50PPyAS4dgjP8AJnj1GtuoaPH4huJ2zcjCYcZASJTgzeP+cBZqR3JT27Jv
8OjiS4pzR4h+hXkbPwEwioqzTuU8zEmjPIHLDwkNzoxzuwD4slZqKqFkx+8s0ErgsAPxQcwqyiq4
irPeSf7Rt+6FRqvsZ8r4gkpgaUopseSUOQk63ZLofb8z/4rzVAAmUwMd1EpB2jnzuBQEnHZky3wy
9YhYQgs7R6YKDVNMZ7YZo1F98los7SKFWXoSKwFiwYOm0NBK2Kx6LfKzaPfNjuRbXhdUgOPXyan5
kEA260CQuYueKn4jJF3gnb53IUIj57g50uM7B5SIq1bgM+DSEb5Nneh2hKQnTT08XpstgyOhIamc
AjHeaqQ91VZteTCmsRVtpjfw8Pxrem8BKLFRRgEF6mDHP+6h67mOVsQoPsJAGLj8juCA2QRnlHEv
z/x+gvJnglGCX/CckzBGNjoKwQnNDqW/Ngb/ulgAGjKgXPuU0E82ri43kOJ3jY5wNScgm539MVN7
AFqd9AT5tj4cUOlcWBnAeM7I4Q5srkvXo0tzE7mDqXejbk7JlpcFHt/mtevdPV5lak3KQVlPL2KN
PtCFt0I0zZGvQUSLLdiAO3oPZFt7wHoLATIbgswxp8fyxbLntDe15Jld2GOtR1wvN6zVOmryZjMS
88hPDY/Dg64OFoKDd4WQeoOg4cARF0Lno/5dhWHk5bNtTad9dApA90WFxuEQfZZ9Zzj7KEbRhxyp
X3HTkQhhG4SitijqoJRLYM8SSxlm2nQs1zyW/rER+w5wOor9AbvlGKpwYr+rtKcUwN1sUml/PGON
ZmajD7xruio0Tw8TbTBajPdc3IndF2LoIiXyXV6xH9EShGJreb9aAXMuU98G/6Rok6qZMEharbvs
WBvRR9ey6qErPYqbRCEOqu8O4hFQuanlYXbF60bRRuaEQcQSol/4V80A2SNwnCaX5AEX0vStETh6
KFkcdB+T4ZBE+Q8QPIUSx0CWYOlcBpzsuj83jMmXxUATTZild5cNpbjeqcC7u0aBks8DAw3YYGgO
Tpwcik4IkWMazxa5BJAEXeYY+wKpbIMmISYmBoNPWPA9H3Oejq6vtaMIwnaj5F0xj9t94ixTKEln
zXpRVfVLGS+G0iZPB/j4q+gAE//jx9/AHb+s5/UFTZLoI+P0TJpiNIGmeI66D8kUeRmETgrF//D0
PgAQRysbJiO00TR7QD0e5aOPTrfceZpZRidYiaW4RDE1QO5dDdCA4wTJD6kUlAlJHWJq/0cZknVy
HD4+j7DaioTvTWv9DGSoHEQs6C8BD6BMPjYb1qfoofmTM1vaNjaY//iKYtoXAZ0Gz/3pRYM3peVd
Hn++ZWR/azxOVra5WAyfy9FIWsPo3fd+2GH8rd3EZmMgb7ZbjC7Y6KtSagX3C7bdifUAyvMl61g5
q06pXVtBR9ltfDQd5BYcwg/LgyhKmuB9eRMehYq+qqhsk742nV1vE0sR4fS9nUiXZ9iDNBNVkDDn
2yAwLeoIoJAUH0PJbFUQfyFVgCGHGhQnwdhy/zl0QBSCDdcG3WGKqfonTAfYrAoAz/ZuJJQ9Ql+K
qWPJvDmzBASr/eTY1QZkBij6B7qOQ15EDXLbaN8sF3WIHNLC1v8y3CH3xlSRDxmQHa79cUXzJQYs
UTXbVdCdhu+NEl3znLUwjp7w2w0E0T357lMNaenRP5npJ1LiPNbxD4cdb6R76flQL7cGCARigmyN
tW+GjDmHX1jb0pupm6Awnri2asWOU3RvswD1CxNiA2NBYDZj6PDd9wNmBQ2SxltnBUaQAm+Pb9vA
mAWCqGxb/Ssl1ysARHOgxloAcc5OGyQum7f8mBmypWG4DBMBOARHyZE6kxrqDl3tPbYAdlmInXVW
olCnle4I4wXp3NmimbiEMgv6cgylUxZtpllqFH2yad8cDeUy4+d2dN09UGGd/ZeJVF+wLtwHOEX0
y9kzLi5WkjGGEW9xP6vyPlVWZgxvhEfec1N47T+dN0p4ZoUvHIbDbsDIgalfOxYduAbF++50IWvS
qgfnYdTbgW+MpX1zXtPcCphRf+q5cuSYEXmkUnAcj1/Rt64L2A+yvgLeQVFdTl92Y9IvQiDUUYdy
cZdP6gA7j3IvV5HQqHVLLW5aa40wncuXchYGsQZ7lvoQj/r5fFJLv8UuA/HEMM89TDvg8Ul/5ihd
paMvxw2IhV+JsuRLBAAlFGzsFmEeMszPHfbqoUhSPmdq0zNS3KbynfuQlrNuxpRv9NZctRVuMkrM
G66oSq+OKLPeVjjF2ps5a2y4BjyV2qj2F4fMVUFOtbIwDNgQkqoNIcafqzbzuhJZTQiTLmeZRoT+
+DXAsdfe7kvtg+tlotODBOUn8UKHmI/TnF8WoH9kAn4Bd7DFtBl2pfOnkYQqixH3UcQZIPrv8M81
MsBw8+bfbG/pEIRuqyFZ2SFTo1Cq/XFRU0o9T7LjmV1JaI2+fdcuVT4GYCe0YUhLnXqaW5bjB7SG
BYZ3M3bUpgj90pJibo4qQSHYwfy5v2XEc3exS2NcKX0DgHNoFJ8PrK5OtRxLyqzecQECXdXX3TgR
cPp0j5LM1gesvDkN5I6gntd8lhkhoEitXsipvKqQjsr01k79gJTTSftsnHUdgk0Nqw8VzIxxwAlW
PNIxrLVBOPV2KvTkv/0JJNjmi7Ir43+OXQhYJ/w3PHOixKnoBcHQiOnqlPX6k3rfCNKXqdi6ZrTz
2r2FdwEP4TGH39Sow41SZvxSRh3qIX0GSIUhGi2+Ot8k11u4C8Vccbw3FjEaqUN180KFa7sCZPgr
BuV0j2kuGPoJTs4RMDBPlGdY51iiPGYQ+8AsHoScK8f8SjzfUCKYs81JS2KShRcDtpaeVyoTOlYs
MgoMfyWWCUbO5aWJXsrRt6dimpJRr9aa0YHsacWmMRf6Wf2eDwvH83n+0obei10ElXBTr1gRzPBv
dKU9JwdELCDu414JArBGwGw9XyO5rpYcmbb/S/2BHCJbLq/3PuWboI2DkoRv3nKoZ78k3kEXLEtR
vdFhzOIw1KZQfstYm5i65wTnVqVE32lRcM3DqbBoMisFhL9PfLSs8Gdub9HufSIDpQ7qj42MMHS8
a4CKITrMQd/wxtGO1BdViW5OKCkm7bbii/mNFFAMiOxpS6kbmczHvp3ZUPBycjfgDTTjwA2YwQJw
77iTd6Rqw+6nSN19egTIGzwCNTwh1xcCH7XHq+VbaSKHNwntT0Mx9EWaiti868aQUoSqjhgV1lwm
cMoSQT6HaKNskMXrGkko0ut7n+K/rpaQSyyyytvortvHGdNmupHD1De7mxkVBxSfrg6rlVT1KMoD
rKHyHQ9wQh1BLmFquvRUU6r1XD28uov+lKty7RlocHlQF/FEwPbmzZr5O8MKyg7YePYMAS8jEpiI
H2vKtFw3wprH8theGWkUyVJ56nyCqQDsTPIjTakGPDcOwiiXeXjmN+awqDx7l9XPkcau9d2Urpq2
YdVCZQphgYIj32Hl2MsU6nkpVHM6STTqCermoCp2BSNw2J5kFvSnZ5Zd+CMNKfjrATUCCaz4kR7E
/chSvXpdlQNef3JjhmMuDyOGqGHMSWHHZ6bVC+w9l4V0C1yKg3V6/8yWqST4W88ZfagObjvp1cPX
CCOTdmRQNroFR1NR4+cBxm6jfD1OaAu7U+abx736S6eENlVNSS0D0qMwwDpLRQeaxHQsGfkxdvIG
90CO+DAW3xfcNUb1uMe2EuZkWxoVJp+MJYrSH2ew0WLGTFMVqQB6/EX30OjCJL4ylxdnXZCvhWUH
lFPfduYL6Xo90B9NhR4TV3SsSXddPTf5c+n0p+7IPiCheok7nIcGSl+82R37RCAC15IoNjwPXlUv
C9lH+BmosY1IVeGOjaPwJ6Tng9QJXW+Wl+t/oNu4jwP92sCyO/umTYuZ/igUCUpXBTiShxvS42XU
DaZvyJY/CK33i3386ZP520WAI6QJ7nK5/wGYGV0UwahwhyG9rqP2AFoz86iikpcLIsNnXM9fLZpI
hrEBLfEOkCrjmfJNQczOWHG/H0hYb4tjr6a6YNTAfpWn3oLd+khVL5L4BA3u8hjy+fNg8Rn37Wg7
CQnKzOKOO1tmnlr/iqpvgYacVRD4g5q+MoTiY07VWyBjhIlP0KbSz0DDtk9ZGVNYkY/JZTJDjXyU
2mk1MRkFJIDLrZA9kT6wz4YHtWQ1G6/viq/SplD2pfLEKvFajUXBE3XEnM2Ehi8nyznRKjVvbbGX
aYVABCVhXyOjdwf3hsJ3zEYiqbG6HdatiQ+IC8GaGt0bPGoKUEtSrpWYXZg9RlBJHKByUYnaYzXc
h1f+0W6lZXKeHl+9EAt6LS1NSM027Kkh6pxO+9MLyxvnKRDlgbVzfTgTyoHShR8swkGFWUvqoM/N
HyGd167CFxPtQfgfGBQ/YjlYh5D7PHYkx7lTsZyrV/nVxNZwAvwrZjV8jr1E+mhBcysBmHwHmc5s
DjCnwT+YTycIJ23YNkkaqD3pQ3QPu7KRxHJVqxEClosfCIq3o7FoT4IDC813Bcz0zFSDWoYCn1YA
A8I7tR1pEX2VVjSjygATeWhImSM/96JaJowX0oDyRx+4+5dvZvLe4kHxdiCVhvUWdjZvGyGlThqS
yN4O7BuIVe5hFieSY2nhI7gPcP6bW3TQjPCScUWXXMYG01uNp88T36LqNENep+iq8vJJsnWu3V+T
IIg1kEUkQP84RUWRnM2zG67bpJr0KYQ8TyPhF/YjIWFKTI8y+lVQ7/BZURn4PcsG5sqQ6rbx9VLC
qdneZatuWIJ5B4GJnirDBVkEXrI+hO1pT9AU98/np9lovqoF3cfXAEqF2nw1pIsO7w8GzAzc3WBI
ZjQ7whWx+nU8bljQVoIf9FkWek+AcVBnfCtf3+Wg5I8k+BTjkqzKVs0F5bE8s/2fAkF1CzNOmiuD
oh5lS3G6ijZscKfNvmhgop84+s4p/rVkV3+GLAnjsKCT/SUEfpghclXEVBeOlj43jieZdUfdYGxR
pIJrsCsRc6mweucsAxGpT/OQym/xxhgqYqAqNtTTr7BxGU6Ep+Jr8qHljgUpMZtxetPC27IrG+4o
12tBXVcABhnn/k3T1BVBpVqtf8D0HxsyDuH1uuzMzCJ6oC6iz8Sg35HBoT/wuxqA69My5aVw0COt
v2LbVdcR+hR6OuDqkbwEuwdIa5247CTZa8RX/yhwvux59HJga18nvKYwBC9KUVsdaFPUcqPsfWpZ
NQnfdarl6ZB/3ErVuEZz0RwLWdeP4SSmvxZ4Of4DyTh/T1cC0NUkZRivb8mzz46IymBeshnKgQzR
gT/zWB7Zo2ytxOSm8RooHjcPX+uLZQYSotEP9zE82h8g47W9VKfEDOpw7Vdcc0xw+GkZ5Pd1Dw99
Oo5Zs/uoZDnasfSaXFHnd2rnU8ax3xceqddluCHl6z+jT4Qzwvh5H9/TM/97wgnBwMZV7F/nC53Z
eWVVfvEJtp5KgtndWshIcnXUS16AGUmBnuyCN96rF+eDNfshwjovVTiQi7CVPl0XDtK3TYcD8+dN
FYcACIiU4blVZpFzsJrS0UKoQ96uf4JZjm+/Mv7KlurvindA5pu3+i0hRBX9xFGtRcwCwiA3pDVr
r+z0OushQwS/IPk4UwNMEGNraPyL+ezVeQwUjA3WJWA37WqXjjorIuHtl+PhBy71JHXFzrrLX0ZB
tUfqCLjF3GcVFO/Omk33s7uusktbpUarx42wZPztDC277Abzar/KG5sOC8O32Xw8ypKAvaBu8bxl
ZLwlyyjR1jeXCls6MdovkXMKGzH9d5V8af9D2QXzbJOMX3dyGWCxzT5u6pmXdTfmUz0bj2wjutxP
9fsbtNxb9U81BCz3sHorw1zwBm7kmx+qqxs0v3zzWxCFEqLx9GIyrmTcEEuS7FhZNIeaurT7gKC5
3o3Zi/0tDVqcpX8TyNT0eeQok7fs0bQswn1LfyKveIXlqzM9B/JLEBIOknEUySSRdS8YbvkUzXIc
kzIVd8P302CVGxy8owEs3tBL7AZ74ouAyiHgIQyZZSpvbyyHcPRDBScmey/MUJWz4nKzN78vbsP1
DV4XPYRdjAm6XDLey8a2Saz6rMdjidLSJdfq+h7fhZAbjo+iAqXyJGyV3zcyF43wnkaFR3+XjfIS
Qo6cQtRSSxKlbohn78zPdO0c7Pxa25MaUa/tCPK2zrGqf5hTpjX7G7Mlq2r7g353xf3ghWWspHd0
OP30vXTEZHli7tTlbks9OigMX7PHthXyXw7IFUhtmH3taGQzjvylZ4JsXBvr7/3pLZck8Gmcip1W
7Jw4P/zOP1clcs7aEvNYfmzFOZc6+rYNT9ikZ7oEELO0Y1K2KpF3nCiXSCKuJpZwC2ATXfZZ7NL1
fe3h0fgzEUswMkSVEWVvF8G5cLbZOje8IUxLjULYE9jbMS7ohKu0cvb8heUMlTW84Zt8s7HsWHh8
042NEcxaUrMklx/zKp2TJqk6R+oXf2u/Bw5bY/6MwzwrNvLmEKYMSE3OPL6zQCl2RnxrqZLTQbPK
Jc1wcQ9g8cZPdi8nHyxxac+KecRuBV7mw24wyU7R1BcX2r9X6KMLQOP1CJt41NiFrsLjVkqc1IU1
Fe4GkxgNjPe/9PKy10kTmo/QWx6KAcxjswsEJE9rdXbLGMpFPWqz/ZCdkM7SYzTqHx4SxEyDWk5t
eV3gOwPelMhvFTG2tc9D4GhTs+bIGDXpB7OWrQ2nPb3ieWc6xeYIJastXGRuWZe+hWw+F3qaY/kf
iRYNnqghZu9sLjTaTap7U1Pt39mhC743uldf1sidkoDQV21tiI9ozqWEmKIe64vHb0DUwV84H/Mj
/oD5POJhv+zVdxg/5wMpsRxJIUTI3TZ3O4KLgDTIAf74ZN/JPMO8rSdRPIsEqN6RyC7PC9z8I6VB
b1ymw13RIOHf22RBJH7OYlR+ud4bdPv8HNCe98RKcE26MYGEIjic99y9pbVM8cZXvwKz+Peqq/a9
kObrpGFfMCe1lmU1Y8A5YesJW+Vkb2E/XTJquoC1W0RYpl3A73a/R4oMVyrijhN3AeD/vO5RkzqM
34GEduuRwymRUxWhF1Aphh5sl7/n27s2o8NqpgqqIAi52q+ZQ0PwkrvDj/iAp0mtzlQN2tiMxEOj
EuDMRa/iPUx174soXF156XJvXtnWBRi2bW/Ey4IQ6I5QQMs3biU5Jp82S4MkrL+XiUm8dxkeR+ZP
J866e+FUICudGwmPOTd1WocCRLZQyvEG28EkSOnTeQN++L3oiwxpo6ZzQQ1D+cPhLVGiNGAMdizY
0ImjuWx3ZEILacoAriX2O0peGYjcY3B7VGvvH61erRauEanMXl5oQO1cT98NErJGfqSecOMBgo3g
0D8H8jQXUeCHuJF1XvCvOxj58utAPr1bikXXwkajUstJ8l7ta51fZgVzfTmHwv5Uezlr2QSfzncK
18oUiG9u7JV53h7qFFEd/q3p/XKu0pXyak+Xr9hV2GZGhrBtEIkqqQUAVvDleRTvM9Q0T1mWuSv1
sPtkIWrTKrbkHmG8UGdWFgwcfQ9m/dZR/o9iDZzXFEqCl6tTopJmM020D48xlfOPnqb81ZHlvhZi
N7nRp7qt5UrhcfNCtHdh8RHrmjiWXfO94IW0Q9CF2oEQsz2armkol5IG+cvPHbf9kdKSwYq8fHZX
/v9ct6xgmHOtTb0uiHVbhfuXIU9U/W9LXigM7XapVYhE7S4CwuPXRko+7zjrdsTui37MCd7LGTcP
4rUSlnM4AAgTtWoxJc7Z0Pj+/fSvKx+iZDYNtrBPneC7Pp0JkrhC+gzqa5lkaAzImDyPwNRE7Pwc
Hu3PwU0nc9vaB2DaBRL1twUd1pUWd/hvZexZxcXHdmF7TFCi7c0oWYbqs9AjUjFuOp7mpv5+TQ6v
bfvg9CLZZV++asryKMjXat964CrcFXHAHoERi1G2dzrQNB1zAUNAa+ujewgP7uQTUHrmiKQ4c22K
LyNpmAfAHGaXJpslh+Fygvw171RsSja43btCugZnooOEabpEOL+uy5dVeqHAwpQkE8F5uspngZ++
X0Xgo0tHcy0ByDpy2fmRwqh+RbLqmpUF+NDcOvF1u6cinfy5c/TAdCZPENxfnXsgIxH4XECSgMJQ
26CZEzxbhC4xR/0jaO1hzZ9ITx3TCYt8D/cdtVsVjye+I4MhY9NEBASOowkDzagRMFbIYqdVlo4s
S31fJsYjuqdRZ/tHatE/E2zyYwkSVm55Nb931/JoWeDfrJwhw4OK7RcmV3pXv1fG99T9xzALOEoB
wgHwywyvlofdNkCGLug1Tdt3WeFXSAcg3Vkjc4kvQBhiibbgo+sxEcUHCz8zkH7bfzKmaYnHBoxi
m3ER4bGHvmWuQ4FdFzm7JsuZIT/IFPkHdaVoxzxc0m/MKKCjS0deDW9Uugl8hFWbqxY3WOC7z/Uh
PnHHDVQRTWu4PBItes8tAHxTbQ6tfsOx/J4ZD81QuCfnQH4SfPfPUo0eiJdICuBHrJtT2S00T3uQ
GYX5UrKOqY0g05jPzTB3BElDY5wYQEBovghDCkPyiXdlGLVzpH7D9CwFFnN3L9tuUbQcDBMvlWwB
hUsqTLsPGxsbBh0bePaj3B90nGEA/ATJ50faVTW6yNMi1jXP8vIzBe9xsFPlw+rRw+ILPljxBuKm
hFb2bqzNSeZaJ0Jmg11vj5YzspdAuI4j2OLU912KibxuUaZBLkhEWqclYJv2dlzPls+a/B/RBXut
zQYqoqYqXVa1Qj4FovnKsX33vv0r/PG+PNhYfSW8VNn3KGXz4EOw3diG9h8K3+zj3rCgCFO3LqMs
afS2UzC7bTyrf6hggXc47lwouYtgKEfy7ZHOwIXlcFLUYpPN6vc1JAngAGU6x3aU6m6Pi4n/sthG
iNme7Z4zPsi+T1rVPJtdJUixfQCWrZHg0zK2Sy92JRAagQKTpIDn81LVwKi8jCnkqje6gP4RRd6n
fgSZbFhqiFHvqnMwyajWsBR9fWAbTIr4rLnHUYf7/ZwhcOBSLoKGbBaahreh9Ewiov1+Mmmdph4m
K8WrtcuLGTsSHQoJwXPcaRPEOdPETEjPtF9TQyeDIO5Ob0Fv7gft8nYIZ+WoOROwtAlyDEa6TzHp
4R+i7QcaXYMQW9ykn8ZECNTu1IMmwyQ5Cs2PzromZIDqVkaOtAOIV6wvxy1ABPuHaiL82vPZxHc5
KIWtnGAzj7vkP6Zn8CD2W1iJj9NHsENYJEoisQhmS8rnc9l4eckTb3/0SOXnVsbEMeaG9osQwihA
YlOZbYoT0a5/DomNwldkBbboGQtq75q+DTnb9Uo5Xym2zwEiw0gaGy5a/a+0stcgkVQIX1UuBYFA
R4MhdUpkq09EX+p2CnkUvOUUNfQRDO5SlQ5syaC3z/UtLEMzSGrDiOhXJQNYCzSJUzeig3evt+lQ
q+P6gz3us3Pv2k6FW8ys9xUbFx7j3bR6bMZNMFuQFW7ozrt2XWReDZ36csxRU4FpQAzrmyUlt8x+
R0Y0+rDp1lJGq3hcIColge752exQzFD0CC/gLlkPhjD5iufBXaooRBMm4QWRdZyBDuDVcW/0g1EW
l420HgJNECT0kgmOeCRYR7ne5ZBoeJxsDVeigj8Hamr3ikg5/+d6UW2WOaPoZTiNuiIX6uMYyCqt
Ywi7Ye4+YItrcdA25ifJ0/lA8yQvJXAUrZVUjbEwUmlkBvGSYCTJ6eep2e7pgzBth0zRIxBqPszI
WrIPlY3fSKItxbM3RmTqkueP/+uYqgr0xp2eD3QXFXZ2+aU1wORDs9te4LxvrJXXhPrRvoh+dQZ4
ysMHEJaSuxtX/q7ojuBSN1ZQIj3bYqOPyijcerBW30dnQjaLQmfbIJ+3rjqKS2kzal/ZIty2mCVa
2Fltn/GAqWWA/Ud/k5qM9LdlqL5xNOtixXI244y/UkOABimcD2KDM1b9cKjWx8xOgkKOXAL5oECk
I/w9/9mT3anV9KVe6lWk3ASmgo5k3c81mW5pfiEBeCkjNmqzNtJ4NA3uGQXfut+qxUqa5VUjucSN
TkxKUXmQ7YapiMwwyUJEirpdr6n3c/cC4Xdp04Udyxz3GxzQIithY4nyZ+aeSm1ZlYc3uvbRjcCm
4JHCutokLL6TNayUajUfz0qURa5dKXJb7Tms6UVOa5Ah7CMBW+pNcpiY28e//uRVEJFJR67kApD7
BHfMl61p/W6bT6uMUlgMUZNm7vbjxc1gjwxdj9dWRs3A6w0FKVyiDrSnZn1KxNzMnOl3MnZM3u7q
SwseSl5rBsezRPTF//d2rbaG+Z5zg94GSl9DbmJZUC0DLTT6YDUoN3kxTvdQHnL2vf4GV7VQc5jK
JaixSzdo0p9q01TfXuNTrFt78s4t7MH511wgp8OQp16V6hGX9AE1eyA1s/wvvB7KKuvP66b6oisW
m9ts8HkKHONONb4gdo/k8Wi7jSAwKWf+9mUUi7yruRwfaYE2XcO3CWgSvea6R7Cw1dssMGtFKwNY
/81DcFifO8aTwPFOzLs+WLDGCMzAQSMNDmyilLpK5P+ydynBopFgKFAXBkAJTbBQg3PYEjwhc59y
1SSD2nUdzVVpBO8pyEANH8ZjEYL1lUNWM76tgSFCxv6QGOfJuoBWN8BBXMQ8hDJOMjGJiZRS5Hay
1+z+jTcqhoDd6bhtAWwaZL+T066JC1jp2Zhz+kUHFYRKjt2rcVGg6+Sh2FUa+lZQzDXohpPNx97V
wgqpFnSx37Zr0ZNQ+TvNn2Ub3dy/KzH2r39jKi68zeHKoTjbOtWQSoMXsuRSM6iIxmxjkq05/+mE
3Csm+EsxlJIVByoMzwHCGbBu4lJsEcw+9nVZB9wlEr054KYxNhC+ZgF747sewl7dIs+U6796IgLd
2TNeDRArpklEIsbTF3qNnwrrQ5An0DN0lPyepU9hlKUC9KBazxm9iIUS+2dzNqSk2R+UiMXqiiev
xTZS1rHB9CVS09vfvBJJLA5L0eSOtdr46pDKRK5JSAwDJAG3PvghkaAQ51RD7LOiWUZkCBAKV0Hv
h5/yvHagKfnGsWPame9EHIdMVaD71OijC3aqMBr6W9DdU+wWI77NtzZ2EltOeJ7tQoPkC5oj2fdx
2oWHsp80tfTzn0CX45LjV97bhclFth2bYyqQegZn5Ispm7Hbbg2+zEBtto1rZbhM2fObI8lUFC1k
GSf8f63FfcTwoy5qJ1+kAHR7Oklr9sQtLMswpIc46mM1atE1dLlEYZJ4WJ0jvd8HoNbFxDW+oSWN
i7aav/E+D7J0i+UWehiuGmXA5nb/xsWQpJHcDr0+DlJbNvSlqnURMyH5Pgz7S+DiuZreJFdhQjcV
DxPnIdqHZPLVybESA3HKsbauWdENpUrIZrqhwZudkUtQsiXCWA+0QmuZPXud5OFvBcnQh1SgxUVc
vtjL9yYTs+axqp0nIwvVJctBw/2lng/4gY/e+IlxWfdGVPvAYGgzfmwOpFwlV52ro8FhDxfG9vT8
ftX2uIZOaVxDE0OILJ6ZzBHj+FYQTRhuAerQyvxJNFcU3V4Q7NdA1qXAMa5B/p9NNa6YmjSa2PFr
voGJ6g153bFRCO3EW1he23pemwS4qI/Qf1DjvdYoZYCL40nkCeod7i3ZRngv+G0Aa2IZ78J/mGOU
08o/5/gG3pXSWIxHIyj8ZvBrR8Nr7iAnzXB7BT063HbjR7VIbgbxNzkPcDRQuEDejXVUeUOqAQoK
BaiUxwkBTI2kHz980038D9z13I4avRycM35GlcpmP9zsHqLd089kz20wmJw2PRRNAashk4CQMoaN
VQGI/BQJwraEZ0lQo5Py+y16R/+dJksqSecuOFDKyEW/4t708eImb1EmKBJxIC/eTLplWlb01GIW
fSX3iLijV1aZo6C+pQdxpnqzH+PfhxVkv0zI52qm4nDc47Viu6nsj/es1zg9Duh1IbyxWg0+kh7O
hPQxt9yRlQmi8/DKMzSA89rZ6eKevXgqDbGoFmdpq/669cQ2PhS7jGiJG+viN8R8GLphBwyQmyi9
gWEBpJaL5fqvBTOQ2Vt9AE4wgc3c3nGgAdJTk8b9Uf9JNkG04NUb89RtlRAQFtjTmZqBBNdqt4IW
Ui5YmkWP1Aez4CzxpPE1j62uty3a5sPtFKOSMhgRPww1FhyXxdsPxcMIWothblDn79/tf0z418aF
qU+pbDf8HXTNJC+loug7Ug56Xmd7M4yJOKVuzAnLgj5I2icJXjlt4J8LTk5tNngHukMSMcQLpQrw
/5LGmtH+FM53S8s//p4mtfAP/+T5ibrUrEiGh4xD10pLMCbAq3hqrOIE+3Od8lpULDcNZY1Sx/cw
nXcfLBCYsw9T/HIpcFcN1vsqSzzGC7rQT7pS6kq8lMjhsajaRv4NX3iHG0PPMj21j2TMIlFhW1AP
PXsiixacxz8RdOK/CJZ8H2ARw5IS7mwae9+QxNWu3SEIJuNnvD2fPnjFplhX1xKWvFwq+HHwrnF1
WM7HUAkgs04wleHZIZyOnAm9QkiIUgFa3rFqxDhfY6C5s1w0Rx4Piq90drLIuFoKl28+eq7LDi+3
ZAtINvy9BwZASoVb27DbyIEMtBom9xzSamHagkyof/ymDLt1wOF4SOtbDPy7RPiRA2Juf85WBkzf
wRvXoKptlhRx3gXFfcuqSpZL91HtM460WLp6REdYhAg7wtlTxVc00KwYMsmAVN5wx6LtMXaB1gB2
4JBhGFPMKoZdUTY8U56spBAoOvywkwIsdmB7TNIZqscrgy7dooKUnU7iwLv7CLCK3LR5nZrl7jp3
AkdwiP2sqOEWUZ+fQv3HbU6lJZnKnYF5qpVeDeoIOlK5tSZUiLdrbHqAqp9vEM8TgZcWj/eUA0e4
uVtvuE+VumTK5H3TBaAUPGDDD8vltartFHQl3yeWtbRnxviP4cm36LkObgYDthnQIgB/j6PSBq5A
gCSH3KQZCuujx1APSyLI3r36261Qp2srbSTXPfVOxMlcm5vNkEQ9qE39sYwRX2Khc4w94Z7ctXsI
vQLNCeXw+rmv3wTpWEyBCUgjA83cR1HQ5//dpHHpTRG3Gf6uyoF+Iki13I0jl0rLhY82+FWrWyp0
Vh50ysFmlxed48/yDGYYSLYVM4iwmxWWkdUHfnmAdbOWqfxrvwEpv+EN9sx/VKQM7iXlr3hHHEO2
vOCVp1TFmLSO20WeToeMqg44AK9msseN1kRQke5li/67TdKd1I+nUijsTBLSpZwVdW3BttXZxVWJ
W/O3iHLTt6VuElUX+MVhtBIXw8hM2+7l5oyyxq6c8Jqb4MKGAPnZsFPQfaWL00OTvcqqMrKjKX6F
zE232iUrXmdATlTzGqp92EAQiAEVl+n8kpSlQfqKE03+IHNQoJD+gbfkZkaCLsWvwyTGAf5v//Xt
Ip8OheOi4LuOtQgTd1Q4ygIOV+TiUxarCLx5DgaEQNcCkwLMhcMQMy6xGL01Nt1IKlD8LsabICaS
eXI51J/bz3OTThDxd2Xi1dey5zIanbDrJrFoiQOsLtMYpE0Rk5NJ0DPQ9vX2h1McJYvflhdV6LL2
+RdE+gQtyBQnPuFcnwYYhsJCAdgVg82UB0Z9BQodUJrtZJv3nDfvSah3DyOazmrRsWv+5U7b0dZa
7t/fo+RLRCNdFQ75D0YWITSYd451TxTBMrPQ+Qgp9EH4Q2YkTBDq3sWBmt01p9Rv25NG8UcsX9x7
w6upBM4TSAADN5ikLKx5LtvGpx/tZHe9Ysl0Vs9hApr8KgCrO8kJ/U5jcYMV2mowgWG/SE2YE7Mz
sJnZjxDN/dMFrRUC0X6+iu7bTwvkLT5dkE/BhxS2KVg7BCu4LULOdX+lKiYekgiWPOMXkJHJW1We
v+QWpAIcph+koAY0RZZ36cSd4XsbGPOf9+OJN6r3DohJ5WRaGUSIYkU/CYs58jiEckwGG1pvIfyn
ahAYirVChFuqRcYj5x0OUsb2I3yQFpb0uBUKTfbc7Vax8lnTyZ1clF7/QpxFPMybJpi7JwZqw52v
zbKC0LSPCKhJvIw2Ad20xTz92YAjF7j533fxWlWlvVLyaLRRGFeSNzuDEhpP7D/eD+y7MqS6i+EE
0jLizD3YOhHTG1OnFScr7B5ONXern32fvbmaSfUin1EiHrC1kkg2FSLW0aRXVA5eJ0WkzChZ+ocH
FTgUdXj4NVUuzTRPTiwIxXB5lbrpcH1vP/iKiSS6G74B7zBSlpl2rrqc/ogDkmuJQvqWDlL/X7RD
IdRYjV/6O4ulX4zhmR2LtvVpmLXDXRf1ezBt3G2wyXcZ1o7BVeiB8CdsDBKvpjj8d3r6lDbQPWDF
fJRk/hMWgYyrMkLmaGHyD7dKBgBKwl9PzO+xoH4sIUHIw9btWObgxWCu63P1B9kXY0fX3JpR4kxL
cxOTy9kH76mJZBlmIurWMgowQJjiW/z43bL/z405tYdBNgxEOINRACw8p96POcji5/01FIRJLAHY
sCUT9S+k7iwKigWTmUDJxBQ9h/yO9vmg/5mgKgA5uXhUTmLYlHU5TRShSGQdMhMGBNsB+MspvURJ
t6/QUfk9IjGpwCaGh4QlZGmMDnsQZjmE4oAS7ffTYlK9wtQb59BnI56rxdVPvvW80KuotXGstWYw
X/yE5zB1bddl27JwqKHvAxfyyujKWiUJTsEg33vrqWe4qNe05FgKg4+ycJchYyqfI2DhCMR/Cz86
S6t2TFx8bjcLIyegkF+89TFEijcRDnvUZ52E3mevAWJdAs9Z5Wkt3QKqhKSVMaJuK3Jpw+oRlDZ2
Xmee7I+abWiTzqV6N2Dr4UOHoube7Amrt+tsQNbhx6YYA4Ft1AU96/DXxr+C8dTVEW6DmgbU26nM
biZWSp6Hic6RmNIjw7JjqWHSIg5ZH0wVBEkancOMw8fL5Q8oGli5LhK90/zASNHjvPVBg+yZp1f3
ikIRawy9qmndWJyhoCDY6f0QR+xtkIdONLxbkJhnYNVgAJVYcgmjZ4l1LmT9Ojb/3MzMQPMpepGO
rM56yIBOkEuGuVjSEI66cG+kNkV+461Z+ZrwAKb82EJspztRP1sDyzBgmP6PGQGN4ZLmibX7sLbz
kqqL9cYyUj80yrA8iLvzChDYyPS0w8kpGO5PSL5acbIeZ31JPjPrBXuDM/S7vq71q4MsEaFaMzpK
G2v1DKeOgnoe7BKAEfMa5UA3BqqKStYw321u6W5abae4YgQmSLmbHitLkjwVmXxuFOvfHvHQd+0R
+7XxYmb/sKfnHGwAv7AtKh0aJn+wPr+EH9BXmT7d/a3fkfgX3BAY0Xv3lKdZ1QOWQw5k3irct9eL
o2/UKiSFbNV6Hl7fStWw+eMQAfLhJTyoDA7J68sYTZy7BJzluFzP59sd1jtS8pCSOVMN5qP8aJLy
GNnOwDFLMpRxXoskLLGGsWxJwFaqdad7tL8A6FD4Bkuqz4HSdz7vc7rARpK0eGxHompLiuVHxPrF
LTapfHANutmorx1C4ClIolsFiZ0D+xqHHdHBeH+pWgszbh9QCD2NuGUZ6LOKAreF5YJLZqXzeA4j
7xOyiQRFSuB25FpZMI1sIfhvZbstu+XBNo8Ag+cIxIpGgaCSqT2F9wdUwXoVAAjPALl8mDmgqOgv
5XsMoQS6Kgf6TKxQj0rbI7nxWrQrfYRD/T/sz7G4ztojpf3ZJ3oBSEWSilbtTjbT3EpHlEIEH91K
TFM5PUL5JcGEnTm14GooeyuLRC6YLbnG/Q7HH7HnW1jU8MVf7uV3AFu3E3uU7f8eUik9pkH9Bc/G
jd63gVotV+Y0jWhMjwUiIGhQ+XrU4dGrmR3qw0we6eyrYNPRIZKeOoWKofdIvmVntlnGA7CLbP1G
s5SzQ3t5TbpgQ398RpZJeDBj5TOj35zgChIMhrJqOwLD1xA/YvmigmJJPFwcT8iYS4h9VZ2hiRuW
srlxpHuwZvJXo1Yhzch7EzjjZlcky2eyJJtQb2+eMppjs5lotBtyx6mqAVKC6RKJoLEXWClXhbcW
kG8IxsmTnRtm7uqnvq2NswDltx4+mS5dFPKbFTiTPVGuzcTDq25VFX/vVIs0zYITizkSuwZmy3X6
KdUVPcpm/oaUpkttFSZrqNZLffN5oRzOsNzDMFNBJcd7yUa0Yg3hhvEYDo7KxFvls/OCzh1Hg+NJ
b7TPDpLllzOWY4Lc/oP193E1salY+OZqzX1wlAjrDxbxCsPJz5voTXPYvgJQjXE1qN8st6t0H4uP
ptOdDbRHPfF+j1lXzE1H3rChGcvgtzGsdUDoT4CrSDi+QmXZT0BR/iG6EgYaxAiC/JekiDTQHeEw
qG/yNPYsBgU10wqiBy/oKSimfgvd/iIToe4RxxuKu8SGUd6Ao9yg1IXKhvKJsuD7GSPlUDoULEbY
+972tSIUdMHXFzrjqYsng4cWXkfGFtemMlPnpDKr0xFEJOU9cVN51KUnTDUiCybN4KqY4G0OhfMc
eMW8auTuK5aZsuDY5mOsHf0wpvPTbo2g2pUGTVgcjxfjTuuSDR58YN0gSK/wrX1Wt74a7imOudiv
KWbdtRSWQquSnvNmua6/iwR8IfPE2cG6GxQrqAXAqi5voJPid4Ve73hlFdcdAQiTan+Q67+GiQEx
Ev/vZTg2g4sRBM8o+kqg+AJ8xt68U8y3m3/yqmfJ6H4H1aO+FdMK3KPCSzTi9CYZyyhhqHlecp+a
cDZoxey6nG8RrmIBKAVQ3e4NJm4rKGPpGrbnAFaZUCDeHsNYCEpJzKw6Xw/h7UGWjFGn7C/GddgJ
SAq4QIgcYtlnlGhDBOcZnGMFwDmrZRWdAAqZCaxNLTCZkOPJVvVRs0GnM6JPcP31wmt1svHq0lBr
zsv10AWELM5P9fJxlIBGktqRAhXJi9cEOEKbG+CxK0tFIFjYrybnhlJZld+2K64HgXZnZKzEARan
ds4M0PUFzd6Zygtr3Pb+dG5St/PGwk9RHj3ejKJb1RszvB1h2QXInmYokszkdg6CbWhmgfRNmjF0
eyvubi47IyUvWrXGiv9EkXJFzDYNDZP49rI4Zk+hewHNRMN71ekM1cCw0OIdsqUt7eStWDBv25a2
tD9Nc39bP12g30CJxa9WBvcbeEUWRO4DDrVeq4s6TUcQpCvyJNL4JR83OOhPFM4oqBjIO9WrIeve
o66VPUdEvdvy2z+cRqXsKgEGkSbnlT7aKKzqLElP8MMIErn6+8D1qFPfD12bd97sZPxfLP0xhMk9
a6PGjpSz/OAl/i1tpYXThdDxjD2GC3cjztNwga5pUYC48RI0TomyDM2hcJYMeryGmUnqUMzag2uu
kIUqme8iogWNjjum/Q4+/qzwh7rjXuAevzYpTVWQE2bGWcGQ937HAxDPyV82k4hGtXa4BpE49TiX
nXpt2CfdsT1oFr3g4pg1FK0lHhHr1/6iyW0X4NJljeaJNPgbGAqdCqSkw9lVstH/KOEec+Savq75
F51v4jBNTSdPDLhntTj0vJt8OBBjpH2l2UAgkiavBiGlpZA9YPX/pJ+ujS89VaeFbQytGmvV9sS2
8+tcE3kKcVTbj2d+IaGRtKPT5ZWhcGe3xgHYeZGzOR/6cTW3BKPOf/ZRmXcjy6pQ0FoA/OnY9+cg
Ams9/k1JOf/71kNmO7x94glt02JxgaR0OoUWqKsIrhFl6q2zw/KoRrQ8BrNsDES19JdOveCxaNBE
jHJ+juzbQtG+PFWI6aSVs2b5M6twEXXVwu/wYZfUDp6o+Wi2WDL5PnScYfTnHFzZlwQeWqkib67m
x3VtyM/UyExnYwrNapecyT+5W0Z6WB3aXG8/q2D138VaZRIOgrpdmMHBKObdk6g9Yx7ILSq9/oR7
J9DMugNsjY7joTEnAPd8PzuPr0SelwLDJiC8J8iNJDvjJpGsRnv2RlQTHbFuzPKcAW3OVtaAvNCi
2hDPMm0MeS4hxDnme+f7dANr8f1H3K4ub6PKa2x9gmHK4icw4U/EA6TBOEhau5XsVEGPNfTbaXrm
6j18GTHnGcKAK54+la3WVgnPrpt/bqdxMYtnr7umpl4I4TyR9iwoLJRH/vGeEHWx8eNB/E4bvRDU
RcEjoeGBvlU3LCJFXIqKc3jnebNwm9Hc13QMCIHJTeIBuTRl8lpqxoo3hNZTcomaEOhiuOYo5nSb
NSMD/po6SM/8UsBfcVplOkUVf/KIjHHJk/b/X33BgcVVt1rBEGdZDraeG0ZGwr9qN7OY/lmXI1s1
Dh/N1JPO1VWfSj+6uppwRMEGpuVcNNsdzhxr8wob0Gvm8KG9A/pNM8/mi0E9KlNbiBBcam2UNWT3
o/6RrNv4DJdFEuey3MGwM/AJ5GiXFk1ianNjBh13LI6bXcEhj3K3rLpaG1UP1gmEJ1vy8GMrEi1g
UxWWAvXB6kxhxz4csnar9UyQl2YZieXwcUEyvkdzqoMvj8+UW9UY/wVBpa/DPLkc0dYsX0MMUSTJ
UQT0DkzJ26rJG+WbXLDKFB1znJYUZgi/4s+FKuBK8C0l9Gd4+sOuB5g3LgATSQ+o0jqCz+JwbWWU
uExRC/xqrCKuxiXikE0knjAjPJMv1DWUOoxV9439OMGXSB1tZ0FNcFxvEL6PMEnAAJnZyZim0ZJi
H5zI12yWjK1k13zr3geXSf+4Yi/91cX8E+2L9ddDeIP7IzLYDUAMUPo3UTqIo9aAKhUFEIfdArj1
aUFDbVMKa74DVsVZBolhhy7/NvNYjS6MA4ZBfE6347fLyLgUmjrlQ0QzTFp53FDo/r2pmOIKPFeE
mS2XZc3Ca/MnV0QgjwKU6zK0pqzCdipL6kG4B0S4Pcm5FeW5+bdbWU0Re9dW6Yymeaz+NQUVD4gn
V80uUXCTjQBwK6j45+/cjUeyVD6r+Th/3hsBVgZW4+YWcBKda1gtev5+a3mR9mkHTcIiNiAcbaPT
+xAi4UlvNepIyv5akv8qFyC1lBrbQ1vLl3dTXzBRe0rU41Ffh26APvxiDP65uWGqRTt4xjARL/z/
W/Fc+7g8M/F+Sq0D5iX2fjO4hxaN2cJasz6w8wSJPlwtVCT+3KPQwQl79nTewrHMUoJIPPdrGHBk
TqRNuPnkZAx4tbtFqh5ZllJF7aXm0MeN51S9OEW5+VXr9S3oxyzai9VQtaoVkjDEQTyu5JBE+hHg
025CRuJ0gkl6P5FyvJ1drqLX99ckc5ErWQurx2nSaKeUmoTTp26sM5eS9GOQb3hjo/0dVukjK9Lh
qrbBFyEVUi/X021/if6ybpWMIXcR9OJh1WmPzGCGTcLEf560EbDCyIkjNk7jvPVVHbh5UJGeZdUB
qNgOhXjejyfJlu/49xxAHnjoLGkA3bXF+56HXJ9L0R1ZrvtEizdWC7BRjpLKkUDVJMgH6A8umBWZ
Hh4n5Qcai/V99hU/rSAdp62KE4lsymG5OSiydJZXBYudYfa5idKwoQ2zwIm2DIwQUqN/1Nuqw+c7
TSTICzDFAgSxLYADn/CU4a2zYQU0pVKfHXAOMofuu42Jg/feX0IFkMl1v2+vhIpGlS2wKhAWM+RJ
pc7AgZxYzX3zheVUueuQam31E1YqbVeUrvNHPwzYkJJ0tSAK3brGg39XIyAqg/T4lS0igWtjShGn
pxyGbTZ6ycddZoX6t01b8xBNI/8e7f0UlSG6TO6Y2tq71KwQxCFE6exCquziu9/FKaPWELWNDqpJ
i220dpPGx+gnb+Xhx43Bdk+o+vvzIa2dHUrzB/RBsh5Vspcu4vDUSS9jrJgFlLm4QiQU4nNjObgX
uktkcDqKIRrOMLZ1JnYBvSMd29AghX8eyBBZWuvi90Ma3hUANqANrwNn4Lt1LQ2OtcV0n7YuV8oi
XDhFImz8xal2i2VNiwDVg2ySaldqZ76gwk9ag+ear0fN26UMMyxEjpD9hQcwcY2E8TfHrcCKBBME
nU30euV+XHC8m0uQT9t/BX5pob4yIPBSAidQ9fBT7YIpMBLK+mMPZQLqMXOrWRrKhVBcIvshgVWG
DUoob4U0i9KI6zPLMgnIzK6C2w22T00BvlUrUYKT6v6ad6f8cyL41KIqpJUPgJ2sAqESC0xdyLVT
M8PeC092ae8BqxFFdsOyKmGJHYXFfNiabz97NIZ2aD3rsOIDMIvie8TNw9dtbwiiG0ZTG/sAnvsq
hfkH6q5jr+n1S/iqLqPxOAp0CsEysCIrN9MWcD/z/3z9BFtq+Dx/RlWIO1xcoPdCeL/UT1QdiUFX
+DrKvO31y6Ao/T7mFNGMN8XjVk0N2N1/fZdx7cjfTgFE/LaBDN2lTwB4RItRDO6vTYG2Rn8u8Dex
6dRY8ofCMCiH796VbzDiiEHHFLETgknUR384/qvCex6Bn4CWJzcUX/Hq7vcW5b6YJZw3mZnA88G0
4PRnXglo5cRCDi2Rl1Sq373D0qzM9MGnMLJo5/CEwUCNYMO913qiTDHNgBc0MweJi1MzK+uttuXR
TSimv9uprAR71qkmNB5YQhp16I5SHj8/v584tBvWTmH4qy2v+Esr7fof3dstZ8PbuUJLD8ELWElG
YDhQIjpDIw+lMC4VRlT6D+SAq/lJM6BbkPoEyt19gk+tWG21IcqUjnGqefiiX+AZauQ/RJ1//UGl
0vBc0dZDp26PBvqrmYWGCf5VbGJl10r8+Aqwk1/IakN+R3ozLwhhPmjTahHljXAlTghod2CITNY0
yNkgSlEqjVRjGGI20qm+BMe7zRuJLuHItG4I2DXDq/US9QVTAdd9OJh8HXoVhouetM0DQ/3EZ5ws
F82yTu3bbJY1f/+FPMPJnSn6fRFcHORXFsBYKdY027e7TWU2jnM1pcsXW2FjLDh8LTzRQWfCTZ7o
/+4lMpmJB6pIjVaqbFhellKbcmZfx73DVpD9KEhQ1kJ5WNU+fg7LejO7oRgbhnhLZdBXZk4dX0jV
N3J9f1icJEyKDf5RV+6vC3UuTScVvT4ois2XhlfKnqdx5kxqZjDWPQPmbYXTqUGRcBwD3iHHmBqb
nYqBnh9HCaeOMv1lnM26B3BQ25asDidzHg5JqNnjxpDTM/XdDtGSIF3Q2S5ZGF0eQn5gbv96v5BK
phvunCl5d6nTjIv1mYDoK6VjOWq9PJdXrwspny913y3lwWwuXPI31tPHwaQxg58yLpreyj18c0DN
jUUC0dVK0qBfRRcUrItG9V0bRu5KGPSR9sEzVuryBl7MEWdbLSfHa78ZWtaf4VJ4LNdWUjch/6J9
CXwmaHxAUo5E6gP35N+2Loi1+4dpLVkdyku8K8RyjcL2ob8zVfyrzok/lKUosn+++n7xBZbD6ids
sBzg0Ia/nQu3ytbKwI3dfmMa/DqhyH6JTDu+I3xIWBNo62UX+tMjSps70NJOZkvbGeca035JMKQR
MOi3Xo1NLhrGuPaloEGpqcUXDcJTtjfHW99OBipSEr+Yg83/pWYHJQnig6s5R9IwVH3LE0RXTzjF
O2QKDFykShNpuVHX57ZamcY/fo4PpGriYU1WKlsTqO00hMEheOBrW+qvRjHR8egS92dkvfzWG0bu
srqzIn0Pt3MVq83fzfIwl3wnYowG/EnMpkAYP8C8Ui6WOZlSv27vlWOTVN1oTNYLZqHtQxVERfmN
16xXt0lr/0QU4O4Xc0ofG7/gELVWVyoXaPx2R07XLK8RwbOnNNUxcXF7X+QKGWd7E1uO94jC8khf
lxIATqnssEuDu3JR2d97N9/16FsnpgCqSXtxPhzfvZo/JXrGGzLR5Te+WFiJjsfY9Vxs4rXvipfu
Ge4WGf1oCCtvm8qS1JSyGdjsEUhFfjuYPny7VaWnuVvCEc7IKDS/OFq4xf8ma1bNvOSzegl4TAzJ
L53WsoaUNx7loJ0cxL7F50/eRus+7BK6Qxs4A/NzlFt+PrNPtjFDdQhRt6EkELAbOs2yK+b+d0T5
KG0ErsYzM/289A3p5eyyIMKcX1tHbkgZmVRnRIAFOnoIdCrxBXlS+JPJ5chNXqX1w518+9Hxk8oa
5JDHg7hAtscDhD1h4+c43RVO1sbPYg4Vogx08kHib97+6t51NZXu7qPweVL1bzdSri/5rZoQTF7d
hT/ysxj8p0XT7IZ/o97rG5bAQsHB4oYbd/YlETqpWRQda/rJHgPsC0+bIHihx8dkVOx7J/0ODQ9O
UNyXFDgR+7tqMMJ3XKy2ZrOflfMAT7uuhrdFHYP1flfgQRgMaN8Gy4Yzhf0D2LXdQuaQnd9QdeK0
2gL8hMKzBBSTDzja40ejMprOxCZLbWQaILqYU15k/TW+hhkK8US4hLMnn00WY2LBuQ8llvltKCBt
dA0kL006JO1q8MzSoO37OhKzDUL6xxrjlZ9Kd+EBugPWUcSKiXS6np9Mev2NLWsAoDAj+wyUEN4g
rchtL26WpLUQ5oXCRp6n1AtoknxKoFuyRV6MtT+elcUYr2yZyVtW7PyUlPvMZwVLpeR5ohmQiKPu
J99IWQfvqdeRPR/5GHgVUyaYD5yOSTuu1q1sUv12ukfgxmbFKxn9d5oD/Kb8pnCJLMNcnlXcZEon
odvlfEywQC+zTOf7mFJYNv+0f9Zah73/Y+Xo0Vci6wtp+nEjjIKice98P/rewFK1u3Adxr9Cf7dD
itSfv8a0NMKKM6EbKpYfSUhPhkNvLXADA2K5EavW2oso/+UA4rAeA9D4ABrgLwQHP4G5PtyMSOme
z0fL+E1sDK0L5AXcD4AE8ODHEXZ3NSqH7l2AuBRnShyVVBfeVksV/41nMlMGuX25T63V3GKoheg2
m/5HuoeAcnIc9wTaxSKE1KXtHCKaMhir0cYa077ZXONekEk9T9g+TVNgWYI2QyEFLeBDNs4oXpQN
Q73GSOvRl7JfWitjE5Zk/OlLap+rRz2ybNnoIt2o8hWksAaZilQF+gqR+bJhSXZp5JX05ehXhXo6
RQuTwTVrcDRv4prbHspPXUNgBoPfneq+MJ0HFvDtJPc6gyUZBQ0wHogECTge8vHzRkYxHYpfxtzP
l+Zj/91Gf89KWNoowxf8y0+8CmIJ5YJADp3nr8+y1Db4GLxT2TEAdL1XbruFijkCa+y6GaslGmT1
+wKHtqtaEgr0N7gSd6joHmZZj/YodYvqeqaDmuaJbip2Pcw7Uqdp3ITj+JkC5xKssibcnvb9/eef
168K0f+53mEERbqGRV+lwVcXX6fJY5SlfBP3X1q4bQTMZM/B+dAVotfnk7FX0X6Gs4U6c3ux0xQf
7wWaJZ/UU5NA4knNK0mteJPRoqQGqLgGjYfl8/UhtNdPJ9OM6p3h/oej3ahIw9ELuKTvgBlkf9W0
Xy/jGg+sy/GnNA7EIv5TzkKpPNLN06PbENPeR4MKG+aoKAw18IqnURJBjJMCWWwg92d4od1/T4GK
8+RRvBZqbJW6UukxH1YIKeXIHlSecyE7NyjFctYIssAstervxe+DSHZNhCcEx0xJGN45lrR8rMT8
XL8xP0YeD6ABwam5J1tO3xSSZgxX81KNqeTsJE7y2YrpXHIiXUfCsxqk9Ma4xBcx/KSHxv5whvcJ
mA+bDG9jkCGJTuPRWuHLVuELbaGxJrUo/7k7IIiUONYFUZIyG0c2MUscgbxML/MODceA3d7vzL2F
0JkJSKKy0Hadpny55EwLINDdEIInVA6Bi1LENPAyyxE1mHilmrYtXs9OS1RzL4gwXtqGUMvFOK5i
71IE5kL18azMuwupco/rKRGc9flUbwbmexoZq1az2Ncozkssr3LTBcXL8fNqWVwBz4NZN0cuSdgB
CPUknriF6ERLRoxq1pGFXdyrih6q7YaSyfbsHPptubPHwhO5xe/cuLal6+M8dB9t0FpaBsB37dgI
d4Yj1aWt5eIzdTJjbykh1M1OKELhBeEzc9MadmYjQ6FtJtDsO36+ZdEUzA9GRflb3xKBo0WSWkot
uaxX3CrEWXdd4Sd1eXWXOx2hhJtDZD1ol/qrla1F2stPBaWQGscm9kgRh6TkPiwHEf7j8+OHNVEo
+cujiKL8F77gyujfdErKZMYhiFlJGxdrWBcqZcZVVzA3lx4ozn41F6DbdIUY5ZvUBsnjIV+1nVkH
CYHWiEeOYh2yYfqpaASESd5GzuYi9wfeuoXDVMO8G4fjg2EfF0dyGO+SvayRg7l1eHPLWHti6OGB
H/olINmnPuGYZWm1bK0GAY5BFQ36lh4CT8JOo6l1kiq1+tDfE8cir+mz6vAmKezoY4lIdVe1WzcM
0a3mjm+90TgwsZAKnSmsG1PYAy0/m/48XFnB9I4RSLXT7vyYptOgS1j4IDKeKigNTsrL4ujtDHwc
fYl7G/mi09CqDjX+yNj+1K/+yauATWYPGPe7+LUESmIhUXaf/sWEWrInitPVy+3Binii18dOoX/0
UIkXlxxRzYUuFIhZ3TzgJaZgMIxYvbeocBem5C+6gOdFZyvhyWOEHDUN0OJj+ITzMr8W5hZJwRlg
lQNAAK0U2UXof42ZSP6DrJClT7lsMaNWClPheFS9ik5Y70LCr4/Ma203h+l+XaPTjW0LG2emCZDI
xR6rDxCcipLgzExQvNqvB5WDR/xXr0OsVHpqi19COM6I+zlEKPTSdY7nZjnyoD5dsk3bA6O1bi+4
Q7R8YAVRWboZ5kf6UoOwGW6A5/v6GcD0zshDt8dPFw7ts/Rd8ZgHA9giS6858CeCgFrqzX4jc00g
rfIc66xN4C8YXuo58JMoybVOyYVIHLnmZSrbtAObYslRV20WcBhZbr46uGWd1Pi9rQyiDJ9J81fN
q1+nMCxyvlmNg8fJB7/SHCgqUoMAgAOc+gMHXuxwNBfyJGN5L/1/UOqBFn1tWkK9io0wO7gvsXgp
MltnWTsU+1n+VrlfBIDRT+bOUf3CQSJPZOSCMMnWQKnbMjVlLSdUYQi18uchmYvSdA/Q3I74KOQn
DWWlsDuZJ5cfXdXWUpCMm5GSWxrTlwDZfLqbsg4Cwqdq7ZW+WxUOKKmNgL/+jNDVhWnWVthpJ8UI
e9+Glhsr0F16VOBy9/VvYd2u5I2WScKGJpKZ7lVxhik5VV9M8dn+fKjPYyfzfCCQRgWxW5EtY/uy
Zz22wupXrjCnGUU5/4K21/HvzzrFHoRfxs3jJXceE3F0ei5zCyWKq98eDFEQm+6Lq1U+hmVem/xA
6voGiRiEe7Go45IIu6ZZlP+UuWHLvCvH/dmQQOBtMuwWJNvHJRnCy6mWpr7bPzD+lkrejxrE/Rk6
geHWeU00Hq0Ey3aXQuEc8dxMESQC/qqRz7aJbHp2yZm0mJd8y1jIeOD0SagAN3O5CE3DMV38/Lg5
3FRkbpge9pEJZPnzlaw3Dj9SV2NKM4N3135Ly7d9jlungLPWycCSoLwZ5F9TamQXe5sVb7Ql96QB
Vh6oHhqJ+aTue/0Uu075+iOPKPJJ8rJBMXeo7H2tHfK3dSswdXOAgP92y70u9TetbXG/3EKpl1Aj
J1hYc7isnH60l+SRh26rkI/R3rmG3plQg+EypXVTS3iMN0dMjex70EZlGd+rzBEtr+HPp7VGGcyN
LJHXpt5Um9b6msSJCF3McHQLupaeFHWvDgW7lbxG1s7jkglsoz78qUTD/WWD9icw5lnNRO1QSOd/
PvBJB2U/an8hRBVF4Ct5T8jvZnq3FjQCTI+m8Ax8x1xDReeeNpHVLGQkSwWgQ3YTyKsVIw+Tid1M
xD9tysJ+HomnyiaMVtr2a+tvSiZSwU0GM+GVyCgmQilDiGDA7LfWI/h3U7U9o/TY0HSPLbSVA7Dz
fndT3Ye4/b27SiHViPCqWkopWNpzWKMkRLLmGb/E6VcfdDNyJnEB2G3GDTjRAgq/hbGy6kOD7c+J
KjmwffTWHDXpvafXqr5CkCz703U2wcwJ9+CRV/ZQg/HSblYu4XhPRqqY9PIQw0PkiwLOVF4njMIQ
MRN9szcRqSBiNDCH2WtIH1UewYbTUBdDTeShp+7s/5Yf8QI+te0dbRk2MhJE6/lmH47NcS61zB/g
ocCDvA17Tvr0qsYnC0D91vnaMw7G+3zmLeou1JxQEErlTTOYdO/4qm3OAfjL5RazlX8Pj7J4tPD+
RwUCQRtldhxu3T6U/G+itHOCN18t/3UjSsDpyqsBYTD0tHzk/uomn1SNZAHFIHpCEJSSS7BC9NQS
Z6UMCdn5FQB3u2P9fBBmG348ywf9dvCy1WXs69jBOHk0feBEITEykIg1eR6lCVh4IvotqXLvRAhH
NQDH17Jh9rDi4pFTRdAVUictiTzfwpm5GdusAmUR7nzsolgawZHYp18LlvtJuG9g/hdG+t+Sx1tL
K6r6ZOBWNwH7/i/t9wFMKT61/mkMYuzDYmlldj16oeiZanzSmFLxnMnGUkFpYBJQZ/MgcChCv7/F
5+dCx9DoIrDyadi8ICe0STD/WyIeDSUPZ+mXxMnKGGNwKf2BKUdz9HtuFU/8WjKySOfGEuu4xrKj
6hiszMN7ZTzLZd13BSkRLOFmKqLPPkIXvC7pXCfdxndhG8ocB8loVzoBjDrdaU5RXQn4LtfgSqXs
jWQsnE27KCcJP1UFbOxz6Nwbs2z8cgG6uVJBtLfQuQoJal4Uw7JMZjC7yaV0tT28wPxPsJ43waWJ
6Gl89mc2LWdEw774XOS24Uu8Iv4yEr723B3xiN3DFpOHO0Kkt+qveZHT4VwbYo9NoUJpgojWMRTy
MN+VhtYt5F70zpf7UD6xD0yldSkPT4a0A64d29af8kxLhY9Y0mHv6OJRgt4bio+70cffFnw07vA0
yekeCc2c58dthFZgwXUzfXemad0AAcAY5uWGpZLJXgBQejKNbDQqgoN4051UPyoChi5WmN7yzL2N
59hlOl1Pl89pKDquOogjhqKW0xGT7M4P2dV4ZUF7cCRH+Vobp9UM5Byt0ZdmjxG4dOTfEqyFn0gi
9/9Qspw9tLb4qGmzCuYRA7wepktTs/GyQipKPKwhocxVAv0JheWqKWnhlHDxsOSBRbTO603ITSPe
A5cvd2R1KmgRJxi90LpWdlb7z6lFmwWmb4VvEjEizrFF6bGrto8O5WLcC0hk2h/d5R9MguG8vjIP
ci2haB+OZ+djYUSU5NkzIN/4sscYoegbzonga0JiBzgz5BpA39LOmAI/IbW5glfX91cajYyU/vmm
QZ2WBwDRO7YqOGSOJKfFSFm4l1kBj25ZkOznLU0K7zSHY3LvS5UMzbGWqyJh2BRuRHcAMMAzR8aY
bEPFJ/8Zxk4la7qtWBZdwZ12vRb1mkSfLNgJdDA8i2NuHr94kEKocKOZ40S+Me8tjInkEORQRZQe
/LWxxFiPai6mVpEoWfnJTtdnA+ZZzf3JDBQMr5C2RhXeItKQ8mt1JEQvDxERYBikPWvZT8NjoBpM
E5DC/EStL2IEIPlR9gngYWn/pXYZVwuSSok71gjLeI80cJdj9JxqkpQ2+nCI8m+FPkbVdgpedijA
UBoL0UPW6wV8TfzoSvEQkLe6kd0qjU/ID59n50i3dhEKtgfvYkRFC3XTfCbjM63iu2KsPVZ0bcvN
/biIcS8Br92qiSKEASAQo4l0qGRuHWdhlZh5RgkFb6yGzc/apmRxS0jQhTC/G2Ar7DzoUaTdY1U5
kcaSJWJm1LckgTN1cv4SNKqL4l8/M8RvtJl8p0ul1FNxKx91rnLYe3YGPEGms3PMUJsNWj7ZCA7u
yglFLx5Hpujul8+xRKVnz0+nU0Fw3cezXq0seN0O+t8zIjEBbqY3aUF6/kFdwirbWANEpJYVbt28
gjn40ctX06oUAae6jM69jkkChvqzzFP2z7RDNPQ4Gu2m4FBd1FjqNLiZNB6vekR5vkEqNsqkktLa
4HQPPFEoWzHHEZvzaPQE7J6K6fWQ7rhTvc2mHVmCWrLr8/trstdaTVBbXTK5eunSy49/y+jXxP1Z
gbbXJSjt0uHasGB+KP4cvIaF1fVuHFhtL/w8Dynzw+bxYFLfbfeNIAZ7Yfg8/4ZTuT9GxwHzMBUw
YIv+sNRaWyaSckchIItC/edtzIgF0wlfBOUrlHn4x2AcWevUTMpH/3KARuaOWQtNd5kjSmXEkBB+
almNBlaV3rUhHeKV/8IFbTJqUmAnaz/i8uH6sXryxYmOyjak33FilFchNpgKmpOhFw5JvSFbDaFF
ch95kK6kniu3rSKpIpMMPvP8QnNuXm/MGsS4sixWCtoU1zLR3UKooqcXAVGn1aFFBWABPK/u6/3L
3TVMEEnr0tTgUOdyK4AHybaRfSmfpgJLOWsogA0SAJGlXAZOvcmHjF19dA6jOtLjr5YZ4QbFeiP3
wvUTnh6xNy1ojIMGDOgnkt0R/x3g0D2Zm1WlvoZBBtRSYIUc18X6vHTm++avQFlU39bLO/wQaQ4U
nIDoNXZZKaOIlvmBYdh1N1MmIPuNcgqq9jdr/y3VjhCMsRWCo5oxx7VawiwPaAXty81JDGOPvsce
bvkrkaJz4QDhA/QV2RgO8qDJbhsJFenZz+oprtSD7Y80nvsXocBlEbr51o8ETGS3liKCqT8/VIMh
eSrBXAMrJ2iGUN1F7Smr3XiF1yEx4LANI1GdDJxc6bna/rV63sIjhPGSaiSABlmdII9Qu2i34WuI
lEPDAvpJ/AN8K4/qFo0evfBk9KPxI0aozca7tslD3owPa4FRJKPMccTeQmt2qewpQwvidN6S+NZj
XxFV6f6x37LRtUK9/YDM+591sJvT8txRi0z4/8wEzB0DBQx4dQS2YXaP+AL33PB7mQxhgQscV6Bx
ocRgwTHAAOqxSoFzPOnc5osUSf74pXbXxEswsTJ4mmalOgm3EfYZgVB5Z7+/wr+yimjU+pw42w8U
zGqkYrqzLLXSD6HUHGZCdiBZXfnE5gcs8vz/A6EShXWhre8sI6Q/OiwbWG+ZwE2rlfFhscUez20Z
54N5GhU2pYOu0X3PYbQC24cJKZ8+zoIzLG8TeG87SHJhxE993nruJN7MOyB0lOziVVvx+U7N2XVd
p1S7kcE4uEockLSmeAqyQ+B911U0qpQAyOvPCOFI+9WM8qJoaLZRoxFIZcUxLrpYvAw6UDJGOdAZ
ttYpb894cn7FmDdsh9kTG79eXYmCemUHT9zXR+dUIVN67G09WsmIcJW4yaJkg2R6BNIgGWOZ3HCo
81YIzcz1uiI4BgpzhJe1P3i+1q1e3eD79fkaP5g27GnN0V3409AzJDJ2zLkbUb8WxnwEvjQ6gzIl
2Hm9OhHRlpOYwLwNj8MNdzZN8VbOAgHz32uAfxnvm0mQtxXE59HSRPnU3c1n4ieHh/OXRWdPOo9N
bYEK2fQACXTNcAvmBA1+sHPNJDqzE84K5LxPxXtDnfg5dtac5hxSQ3wfRjMgQqDoEBMqayinJ2Hr
8MAtiHNPxS/AVXz3mL/QtJ2HgBVg70cBDbVgHTjmfRgyDVMdSgZyZtXArdwfgSt36q6m645Opd4N
Wk+26MREx+kRZoF5BPa/a1Xe7NS5tpc3j9lUpfEqgTJVDqtJdNs/MoPyWs26ELvJR3FyFrAIxlUi
in51eqdZVEyIAFOuYX+T1Uk7eserKJPQeS6ZGl4Vl9d2H3HMafRfkhXIWVyz0HYQGraezlncZbjk
oEJ+SdiGzdpo48sjre4pDsI53kC3ElMnZE196fYnC+2cuIGXaEx+B2NKa2fjusjShzxrhL9gHldv
gk25JWhY/1pN4V7YPCNsjVXwho3C64UnHMHy/Ufk/RF4paqurY2TYiTiAlWmpLzG9bZ1e7GAbZb2
JoK5+HUTCX1DrUnpTOmvp4WVjMdydja4/Fuz6nw9WdvgapzQkbe5JWkRvJR0BxcnHex1e5KEFPJh
tuD3pXlyLrZQbKGSdYXZG4+7u8hVpKBoH8f64WtbnSD/V0Z9rDST3XQS7FMguDPoQSO0aH8e4tgj
lkeCiLw10OzDrfgWKpUaSVw02H65lKE6iYvqIGfjFdDrz60aqj8KkZM7AizaEUddmGf5NINzMcgB
wTh0cBKIfum4Tg3jfljmxS8FQSBBNMVoHm4ucW8gO9LXnHoIrTch8R3TE++Xqr7X4wKn6grtTMvV
ZcyA5phjVXt0IkFPPUwMvgciHzaIKaIpW4PYl0EfwXossI4+Li2++U9zftHHWLGg2nbrniGwpDRB
dB9bXzoce86/JXpGP6rczIt6mIkZEkKhT+O99/Eah8hAYUQgI4Qi0b3gJTCKfz/509vM9qbAbxg5
VeagXy+BT2X7jHyWzhTWFMi0gFC9jgyd8h0aHQ8GEcObd8tXGweoRGHacxtO5+s2u0NDLY6GN9rd
Q/f1pIdFcXZ25yBDB/GYRNHKN8e5w3THVt1BiMSZpm/KLAbYVDJcAhddlSzfN2yY6RHcG1he22uc
aW1y6wHopXfmv4fb+18hfxhluTwANYbVNfDvqDrkzyAceDcPaCMfwAoEgthEehHSEU2c/UHNqJX5
74UAmOF7OQw0dgWV/y6reb3IC/9R/9/1qG74Z1f+TFR8BYrItn33VXrg4JstD1Pdus4A9JUxiUjd
0F1Z8+8uSypb36Eo4QdZ1TATNLwKAnmJ+0W8ZgOgZajHQp821SfraJfvHabpAHpzUTZLZrlqeSgP
w8sAjXrp23XHJxQInBgtiPMMFRWhSji+pETsqb1g9CuB9ZulWvj54mi8zNtYWV9XV5zklqcGZrHG
gv96mZvBn5t4e3Tg0IKuO3g98/0XFVlGnaInhxYmKBfMMMQ4ZrSsFoDcvInestxZOLkQMmNM9nn/
YHkQYIT3W5Dlj8tzNFYeqpkS51T4Vghtqq/NdqbMyG1pS3uyCDgzstUN+csKy+zzZzuhdmMmu5So
+joVJjt3MBTIvNodSYeGTjaOtJFEw3Vy5RAO3aBE1CUp1klweu1goGD1chZMBOlS1+apsc+VYSUO
3Bt61O1AoM7wjYKsn/QJjwLLiZF+6WTbv99tG/e5BZ63JBeYtGLuXPyO2yszYzU91BcNh+AObJfi
fKYw8v/J6JWyjc7XPBBQ/Sx5rNBDgQnZq30pzxzYJVwDFbA1NH5oV9XX1HUA+3IhLkfz8huRxhvl
bcmmokKi4TqPK0/wW5kXWAWsyeyB019E9mcEvQuhEP+xDfEv6yq0H/rFVDPh8DbiCe1EJBzc7AzI
qK+2z3fafzZC6VucZfbdNFGQfLpvpi9tK76pyTXoYIobfaVlLrthDWbmwwVwBP/Ecd26zTbjMKQA
MlPG7Sjp3NI7AZ296CzF8uJ8Yn/6I0fybFcoFkpyD5+7XqDHcf/uBLJYtYllfs8kfGJpx6K2MFn1
bPH3B/EndKUMQtMKu6S+ZXz8JB10Fglky8N+yoQi296eYd/nO7hK14fLLg1sgOi9I01sAU0OBMTa
TMmCOnyYeQ3q2194830IhRhFgYh6TSEDacsSS5mYd7n6wdy+YK37CS91gfUaNio+SiHseFIEIlkj
20xHXW0UIgU/WfLVVyKNDXrwsa/Y8MlC5Xj89NXeWBZ1mETVcmt9R/QDeTEMdYWdTutuYlMytYvX
cuWrwPrM7PzymWlVlWgILvGRGOIrPaIDMbtKl17BRYccR7gYLnBqZIhr6w+Z1dMewkmpCDbNEhUE
nyZac8qJqsZ5kYvEsen8lyUb5oiWWpc5ayLNvNw9RpU/M0kuhzb0rVN5nGOUMzOd6Ugo6neaUDSD
Hi6Wy+oZhUfm4JdWx3Qp+k6cjW0vmeArA35xf81yDhMg+Pn+RtEKOW68VcsWW2Jy/fmMt7qHXKRW
uJQBx3UZQeusQTleDS4Rj2xAwFDxBs5F1kov5ZsfTvyCMJ1+dB5OZyerSYug0pRNK5fZR+sNN7pv
yrqvcjfsjsAQRKzID6ypOuyzbBfyA0rPpRF89go0MmAZ8AtntP4qb0xz8bF1gxCE0SpwuNrv59l6
PBGXrS6m2P7qiTlQqYkeYZdHPHQ7Z/xhBTeipEt8WQbfQaf8SmcRPGT2n0HsIZ0hjhPgCfdT39wH
g+nKCgMIhNB117h7eNqQf/rwQ2YIbQhGHyiYWRRAdVkxkhHmkfl4LlRK6QX3/C1x/zTUIAYvmuUd
Ouekn9zMPVyw1KRRHAc4XTHHZRb++ZOLzwRzSpPk1zBF6W6ShDFPiAy5LxKQhHPKoZzN+0PNwYgZ
5IRzEc+UqO5JDI2/tUXKcMUehvf4UFQsQxHPBE8nWtwErHlp80Lfamt6VIPw1fSyndgqFUjCJ484
3P+iTzatLAZ5XJny3CVKtguokBYaFxSKDnF9asnWsim/HhS0zvWdU5KnAP47R8kFLczIiXXAQPZp
xDxkewnIEpXuhjBhiBH2U3mEZ8HFOwAIHBnbSaH3V/KmR6mDRCHB0AltW+V53TI/bn6NU0udr2jA
DLyvxAq9FX45eYJqXEcyd8w5eGDYoJD2QF5Boh8YszGcROK9IoBn/T7lp5Lngu+s4pLjJ7Uw1+ds
J0AX8YxTCmaZ7vJZo6Cq39bDwPcgnJxSTVpzHpgcLE7IW8I6OyRhi5WD5KIsnHmo/PnDke7Ov2dC
MyDEp0LATwZPoZxjrwo8DPCyDi6IuLDqTaCT9vhp7+kiOm+ELiJlS8Mrij2GsHgZKtSHfaDeN/rE
oiJ0Lk/V7V3+K1lsdbNGbhJuLzr3trAGQ1N7iGsu7KSKo6IU4G4PLwJeZ3vM+xLJAe3vaEHV5lcw
aNWXOAHQ0kcSNhhwJLGjPnxD8x4an7bmpcVSnKfDYpEJ6fSaoZqA/hSebqNVZiD9mXOLUEKqjgdF
OoZyWCUOXSCTglQgyyxGwy/8AjagvC5SbWoWsAWEvjdmr7DFEs6wzWE+uEh1RbPqSCuRe/ftVRSB
8dPNXIxEY8zm7+lPBGjROf6EMVeBq26oUpNqvHoMxplmDPJ5w/ztn9i6EOu8kSD5zVWj7ZsDh00w
KLT7Z3pHFm+uO20bC6z5DfR0RHj+n0umtuIxKLbc/Lsg9Pp6X3TmVYO1lOp+4XmgFjqTHz10wy0K
boANWCFbMizXcEbaToJy1qWcofOPcje6ciUeLff5PBezsUG96lPd4XpKkw/LMFfYZ8XEx8tKhqX5
7Z0kYeSwkGUE0xyaiuLvShj9MQYPOQFse9nbrIf352DGeUEXAlcYtVvro5yO41CLwOnJwgHCvAPE
OA9CxamuiA4TwqJzVAhQz68s0HPhX90vJ7Uew1xcMulAVBEi0suvUlis59t8OZ+icjQ5T4z+WOfZ
EnKzBVqGsE6KQc8KTCTKXPTkTQA7Fq+j/TJBerQx+fsY+ASfFTJoiSuVRdIv0PproLuTtW7eYBms
HMLRtAVnNFGyxB4sW4031dlPw3k/ae2a2KljaTQbkzfggVbheJTlq3EX0HmsUqzvItEOXZ15vrdn
HJHFQSjc4gPTXLsEULQRKCShJW6jAP4zaZd2jx7K/SVKAejSzdPuI9WIaojtAM/qNpH4QV3Of6ug
Hd34PfamoUt3lyEAePITwUDSnhTibiAwZlb4IoV6jBC7IYIQyHINmm2yjAsnsORLojFE/mH3WMfE
C940YrmEOkcvgmmXB1CoZJwtOP6Fd0svEpad2pDj85V3ibrh6j8iDCo/3R/cQa6q+oGRkFC1xKf1
CuY+o4GkZ0G6b0pENWkSrCuo8ft0dIYB3lthou1Lt8NC1vP0J5YH2A3WX0NVlcMd+3MA4KYJdwpP
Uyrknh3WfXJlVt9E8LNsYQnGtsn3vnUvQ+bo5ci6rr4cfwc3TVaDR2ectx1u2jwAPgSbLhHdRp0d
6tuH1EMc+YQbFym7AlLDHfJC5A5ffbCsYBglcKXr/Tif9KEvVUGk7YLN0ZsywyhdEbyvrBSLt8vh
SLgybSnsW7niQXZk35af/5K9yenErgD8rQ9zDBU/iIcNtP9mkPgLQeWp9Wp/N6LAeIfJVgcvsJwi
D0kxB4svw0rj9Zg6+49DBkBoMlinL7OhkODUH9W3tlpvdRJ7x1UjRg12U4xgN3NS4hwDTtskwxxB
/Iv2MVm+S6VYoxNlmLeIkgYchHfyicqUOliJBalU+EdgDY6Mpn1TWLnljYGRWtoQ3f5ySLJMhzTA
7edJ2pdjsfghqUetnyFJkfkvHIGLZXO+1zcHaNS198FEjiU96BJ5OFVeSwbr3BkDq5NKec/A/d2+
UPcRewY7ozQ2H+BPj0csGkSjPatyaIeNXibLc9wyZY5IqieKshe+nw1J8UJz4KplBvT6TVS8Bmnh
XTj/8Q/P3iRMqLI8li+sjJgF5sJNonuDURZS5Z4p15a7XIVcuN562dOzMpbDYPlOl/vUi35njAjj
lQj2/ZnvQ6KrDL9dVFqWcRmoz+/Uhc7C/V1juBcEwDbtZDImj8KhmfD/u6lm8nHu+Shm94ZSItNH
PWducKXA2DxmBQlgCYzwieEFBZnbmmLo5MeUYbFt8AMxh1t3yT/QTRbdmgC4q4nZPrLHyHqi/yaD
YxxLuYmOoMz7asnER86QE+g6UrifQ9Xk7sHOlF17pIyGkVB9ZU9iwvlduqNTstxOnqROd7vUn/oS
5SV+8bn8Sm/XDWzHovkrYKRaFbvPbjap2eaoMv5H62zvcGoXLTDEoOw5TNkwmilfmlbTIqNRxLgr
rm+VqLRNugNO007ARNwIDa4MKfuGvnDudJLCYEok9ZPmgK3jtcR2uT/Yb3BLtn+9AF+5USyw0ekD
50fiMjU+kTjIaKCSr9S/3AsLKgfebUp5GiWSovf0mydvAaAl/suMVl8XYk8NWsgzHGG72KaWboNc
ELTnG3HyCowV8Pct+PW6wjpJQpyfrQgsL7qoeu+DLMer19uynX7/Ud82v0MSQ1dGl3bIfDSV2nys
aXCdpA0LhU14Zz+t/XrnR7OumIqXLPGYZmPTa2uL0CTXqyUG7JRF++uPfDjKN35NO5rlF0N/ZWA1
19zU3Cj/8bKt8YPSNz4QWA2jSBshZ3HclTm+W7aejMHIqaDl7ZrqlQmX+TINWYsd011c899UasHn
nmVowX99Fk71jRtNXg5OGwX1EiOr2GgwBIqxhuO6V1MpoH2IdAssp2pgIFswk/yLJIH/Hgjja5KG
9N7opsWT89GhyQj5Q5nAklWAsHV0Qst6wbHZuO1kbODchIkOj5bOiZeQUDsQZD5CVXuOzAZHG/z+
9XavjbG8b6usqbDjhPreqvXgkDh72ZA8dfAedJBaqbXZDcskbLgWTG743dy79Gv6/NF1H7TkndOn
W7CG9CvdSo3M/tsiIWkRWkFoUHAjo3Bz5H6XtZ0C0fx6YLfFbHZrozbsxrIsmaaGgymUAe9/LnJx
q8YdjFNlcmIZuL9+FIRE7Cnf17ipxnZYMW5/fvV/ln2CkGkNf2gAGTfMmjLeAWCVjQXinhwjHFcV
5EdFWwu760gRyOyzLKRzWx86Iop47H7ipjbqVkjMiroQJSO0q+jn7rsdq4OLtb/wsICLLQ6DENrF
PHLcGTdUnzNehmzKSw/8qz7LFaf7r1KdkbGzBVGwSPIQRWcqPhcw1rEkmEUO7liI9ulA2qr9lOr2
myOJqhGgN8b7rDUVACeMpEpsVGrDckiQ/TZtqGi9xg2PbliP78KW/V50wkEGmTmhRkrvLXuyDlTg
+LkK2LwX9LwnFgYfrxu5PLhP16v4UA0e//gill8WyavhBZle3PCavBM146Epi4pBw1vClHzZB09F
ELXr0VixNwh7q4zEdTRPrZg5Y1/x/oUvuLyHpMgH2eXZuewMeLov6YKc0x5rZiFWPysCTOdoJhmy
z7g7XFfo0+vOc/oGFOaoghPI4Q91MspE1Vpgip4yxNXLfJqbHetuGXOg9y3eOeqX1tGAWQ2bLaHh
T3IVcykWO09SXtkIEdaHzn+59YfQiaJqRuHBiK/iDXM/YZxnQbY8LSI6dJU+ypzsaxCwFc5YlKF8
nkrOVbV4daDLaRga6v/hV228bDatzbZ43oN6d6pGSnHK2VSYiJVHaA4Wv6t13YawOIlQWd6meTzE
MSyT3i8+CT+bXqi8e8IMYdILjSs6bEgcza25TL7f6epwCH79cSxBG3DfoCxPsWIFWotxyg4OVUFZ
cUs68dtw2ZH9wnhxwfFWhimxuHXUXCqSAbVgNKYMgQXR+Bxl2u+JRbTcBFUCiZCfue3w3Vd6M8Dt
nPi8mLY+ZfCA0M2QUXsM9WZYIAYA0KZ0QeetQMSQDuhf9iLWFMBvTvcHgbu6rHBVrveXwenmSdwA
xQau9ZfmHGyWtdu61MoJqFwsnqSWNs4+rXFMR+Mb+42Pn4kKRkbzAqpcPBNyzOnaJ5eZPPa8voPv
qF0eKd/2LKunC6rt0HOsgSNT52iRix1xhrmjJ+2TPWympXT0ECQlYpwrXFxc2G0UWHm3mpnUf3Sv
g5ZUAgyw/lf0DHHyoNmb6e9R039w3EYLLWjqwv+KIg2ixeC0JOLHJPlTetBPt+NYrcfk5uHWN1ok
+5DxqpKQ9da879uXSKPsBY5ANfEB228UvY85qOCK6mvAUE7Nuse04oyjHVNOsNtOWu5sMgHNr8OY
A8jN+awup/QLZSotHEHRL7I4d9FsEiv3yhi6THn3LKxxomTYZKm2WYMp7izG5cmmcn5JUmU0aYvp
0frliJF2l7L2vGzyikKWBEwBdvnCgW/NNIfa1aP5/+uvyGfugoJPa+ujapPZ52rxlTsFS2TXpeaq
sw6D118evjATzBTb46rC1RwdzSeqfbxtdHs/gr1wwjM8ls6srw8xxRfuDix0OT/Oa0j62V72OOJs
pKQXz6MHkXWxwEepC9XnN1WGYNPVIz6SWCVNxE7gcVdc8OZcx1V0oEk5PPh+KCe2Ho1cevwnhAxD
H+VH/AAT2DxmGlZ/hiuFnjEa1v2Q8dWRp/u4rsSo9RHa/m7z9nI66yKyWbekIzL+DhLOANDv6QIe
2NwAxH50dWuE3RJ03tdU23RFE5aXYXkpF+y9LqYoSeokbq1CqrGEj0FHMnnKgYS7G74fPiIIMYOZ
D4Bz+QWhTgIk9tALSueOrbWhGhe07NVe8TCwwOoKsJu1Hjikz83LnBtY/FfVeNX8mhhm5CDgPFxa
zaT1ejptj9t0qrYjyvy/9FccTEc5k7AFJ4rZD3Dua3Fm+0wsa4iUEiwx9O85f7TsRbQbYwcJ6esm
SnWpCmVJvWbRdtmQ01qWyzsEm9twQkjEwGaK6BcNoQSxlJZK0yU51KC1kv6GNd/hjQjnPEHPMAZH
lM49yH7rWoWeNyfZOzfkTV26XHL9tjP26icBVfnxG29cOWI9YGqWeGHnew+zzu3kkckU5rgh/lGp
Who8PNNjJ1Cgw/ll31FBv1RtGqJXFVQQwDKIkqo12GwBxCIfD1IL7VeJLBUONEJ6l9XP1cdohBrN
jAeOJxwZC3PnuwA5svbgFGomZPZ05SHTTz9So9mTBG5NAcoeTiFQl7AiSyE9bGtvJA+d5ehJeFRf
K/kM25tjgLW0ooJAIfWW5z39tOdMZigun9TMVGAtMIcSGCP3/b4tX1/fjqJGjyyYvgkgACKe0sgJ
7zug2G+ieOgaTFObv4Z+nSe+Pil16dfq01Z/TDGguOEp/judu3T/BVl3VZCmeh2r8llzfczAid2O
YFUVpIqb6C4K0hlqJ9oGL/92DPnxUNAMwQvxr2uUbDmP0TU6nDbiKXLA1TDnSJn5bx9zQTKMTdrx
WQeDRVi+R0vWH2TpQJp4TifZCGaHHSkXlCBIdztOaPeNVa4dViRKVCAVxfZgmNphltbAexQMzZVh
Mq8HvkDQIZ1TJBdm65+3rmb9tsaTPYYlwC8EU1x8SjXHWltE9Ad5vpRXfogxuRhZaq6T+fbPuteQ
qQjTDO0VSwValgsadv+LyW1eYv0cckxmfYpHo69tpZP+/MgioF5QtMRnWE4XPZ3L26URFnqkTEsX
x4NR1Ly7yu+3gGTZdV9MX+Al51REir9DmoSz022YtmBbcbAl26hC70KN5mYpZAruIWIpy2V1Z+yO
uVhfMMcfJIQXOn1+HeaPqm1TG2q/D6HkivY5jo14fdALjKmYvAp5xCJjXcPqpf2HkCgZtADVbry7
VCSxjoCwlr3WdzI6CjpcHMlkRnaKfUAS1UqZCxKghgEpjIVwFQvIgEg4f1VDLUHy14gBgRmK8dd0
6Q6qk3jytCi2Y5CBHB974ThzC5BsV0PEmUbq5lvZ/Dnst53CD+xBRXw/MjQi1lExdkICzvexdfub
3WrWHogwAaL9r6XhAu45qEODrD8vMtI47pzGjsm+0KjtM/6HYn9f5P3LORysDR7uRg7Lj2NWjJL3
jfDw+ErggRsDiPKPU+BBV+rnaKg4Mwqexi1RGD61Ov7ikRLLROUKg+r0FEjNrow8BBR1pQGb49Ny
yLzfolfjyzf9evmKFgbMM/dbpxezyiSnWZdYnuWNlMZbRs481oKGw/LnCYQnm7VdjhZ8tzpAXYdU
6VIJnD2UpsawWW8olX+Ej9Nid8Yh8MWfcWnqS3bBCadg5RK60cDNZP79XE+XhwzS1qFcmthBWI0I
ykSxdKjRoF66p1b4lq77ZnKadm4HZ3IH+GDmVzl4KTBifeLrx6UkphZWGujnA7kSn0Po5Ox2Jbuf
iyjn7sCk2MvvJVxoTR9x6k4Xwp6SSORTaOOmPN05TOnvqdwDvJZYVI8M+El8bPeCsN9fpOJaIaH8
+fx8jUfyE4mjYfezkruuPfvi3AXCJ5fE05/5sr9bs/Zy45e85cco0bZ6kEJ29hqq7vsEDcGwQAVB
HrgTBGSpxMCFlg3agV4L1ALhSC23X8ces7b+r9MNjsBdhi2T1ioBHje9LMZdUiplU4cp/6+7tegY
c4I9Io6vJZB+W9yOo+mlkFNiZQQ6El5s7v8AJI/WcITZne7UgnquQhcg1+QYPfDpfwIVPlER2PgN
5sensi2coGCehW2bYbw0JTrjKxL7KW3OLdgh5EusyUqiRUvKcBI6bBLP8HZKPcOOZ6k/fMZLdU79
hbRFKE4xfwpuIdgkOrqrO6gnEBCNmJZ32ipsYpSA1gJ2WmsZKkxCRR+0gfQjA8oVSxtKjZCs8vOt
VWwhV29fviJ1COOT6C5XXjoIdptJMBghVrxjGW3pyiwUwS2+6FvCAUlUu0tQUSc0dJb8OSXgHJtz
ifsFgDH/7iopl40K+YdsuwGLWaFyPCEXeEIO3qQl1Qs+nu/W0Oz7A/wJS4GdAmVyAbCzbTHAffYn
fAtzjpmIsm0K/e8EbT1uNxIHHo/d378xoSSBmHhXCyfTjd6SLgA3vVIzcn4KqKr+BNxdk+TOCR9a
17ZFxCr+mqZo4hhaoXbYifE89Sq0q+hwP2c4SNnlMUyJVWAr1pnh0C/bTPNDBfUCeA1APQ2zXpQs
v3P/rcyb/lMOU8E9z4lC4d9lGuEgERhTqRgURri+bBfsO5OOjIXmEmEYK8NnsgenOvCRSsiylQxV
YoysFn84DMHQNX8p+DQmP+PTSn8AYt0g0Sc78BxGfvsibbSyWqBsNmPJxd9NjUFz9QrF69q6q8lX
E91Bg7XcYvJmJqsqm7qAThJev/nuvLz23wBLtr3+EFbkPTEE4WEi4Ue51o+k1/BbsgKYoQkcYynu
ueDIqtA0S1w+KalS7Q02Ha0IWJOH2UH5albPL5KiXMhHi0309ezeUb0D+oBjHb3if8n4eogQOHXf
OP+Mz2kjt0slztNG4lwW9SmqzRoKdJaAZxMRCF0taqh4yCBxuXIXAaLsp4gIXQTV/Q04Zy89TR94
i23kpTwzvoKCirlFxZXd2wrFVAmaoLwKiZwxnPwie+lgWXm15M/LxwNXE/7CxBX7ygM8btnLmSw+
HxhtYM+FvyMl5r+99KyrZz+oryBXAaIq8KMObjPPkQsAlqsV2bRxVjyx7tZudzj8RMmK73gKKGgo
ElJ8pdo7KtdIE3t1sJZEWRW8tH5RoV0VMBoP7tiP6Au7VUv7Q8jumP+/3mhvVlpxjzs0/SiVdfct
Hq54jia09MrCLCNtTPTPUiqjVJ9VPTuFYQWh3C4qzcn6dPcp3C+lkdERhw8qzIwgyT0edDugRFJy
yB+5DcdvrD8bN4QaeXzZVHAS/xulBSQ1/OTW3CGj3dIxoe9KqnccpwTjPtZAWHjWN3d9b3G6VAV0
Jr50L5n9crv/DTx3vum3N1nxs6EVc+WQZWnqA87ddMSl0Gw2QSW5UexWqip67H0MDD0mXM6fuT9u
MDGvSmcG3IRcTW/ftYijI5nB6gaso6fqd4HkFP7nQgMIpAgM5yolw1lubMeYfu9IjYefdD9g0Zw1
EnU3vOoLjKbZyEDYoZu328c4CMVT5TsZOEMyOuZ6LptqIIkyIqXC+TxrARMOxaxJJ+hV7UwWlACv
ujCjOhW6zYCoz17gA6fi6FdhcMu2pbETwmArI88YoH2tnlo3SZlO+rIz273QuX7d+DF/NtBuvakz
F6x1Anklt/L+hcOhmIfVJV7AUvrfWSWuJgjWC0qToWXwkH3mp6dBYR3EU7ev+WbVL/tTE+v5J2zF
aCCI5gy6VHMLNkqRdWTKwrISTgZT13UP/xpV0Q9tI82aY0E3zV/j0T2kzSSiwcWAYkmSB87/vZTo
0NAjowQwH+37hCfNBWbNpPrjEuagdtwT9WeSZdQRa+7lWgoBTUAjuwi8L4i+whUb3pPlGaqzkXyX
GnheQ/lMYDAHBuw1kja87r2+whNQ3Jddk/IOt8gQtzuBRaTqL5JhRvkwZn/t9C/llExI0ZKd+SeL
ZjiIWW3ZthW7f84VAatVPPXGjiwqX3V7BD1ZfK2ZGenrPw52lG6FEioezDddLF/59mJ/VRhj6Bb2
vSHwfW2XHunkd8OVtYn1zaq0qV6XWpMdChpborjnbAL2pNLm0IFYyTN5H2tT+5gsDWdv/xWDPoml
sGsa2yEUReASmp4e/mSl1sOd2Xslfz12Pj9SwfpY5+MPnuOCWe2B6QizdTM+mvPIP57bQgXD7yqW
bvnf1/p+YRGPw9V7ae+YHRAKLp5GrWvEKnUIOxomqVEqZPhnnc66fLLDTPxtVf9p82K8A3Tte48s
p4SE5lFRXVIkdBYgfSLG5nWsBP6BcXOw3rAYedvIoitavaemw2/VoLu0d6flyl1y5ihy/lP36q/X
PvpD7XW8AZqP3tmBfp35cZSamQ8csPeWjERewGDpQUR9Mm0QKlP9I/eh1Pn3Z7SZPEpr5OEHvKjJ
9IOZPA1b7nObbPTQy1KuTqiT3OSV6ccqzHlXwxV2PCMFLm0d1RY2ZEZ2l6oUVrEesQZBMA0uuIPO
e7UDWdoKsGgzMuU2Rrl/2TXFpojh5NBedaYlUtGRZ6LOzIme9ajyWUBN0hgCZPhQCI14PieEY+e4
mEM+farOrDhwY/zIe88eFdgO7TOB/UOsx8kyjY3tGWIq18or/gkA6P0oAqBLCl+DC+zqDjLHs+5W
Dksietf3TkXghlsavT+gP7CthQezoLG2lma+mBF7I3h9KZGDMHLzTK4j0WqBdDnp1B4xnyBx09sX
HgHacMifkdo81yYvR4BQlX8lU9wvcaxrH1Cq5lRn0n49o7lC9QbQ831KInNQQMk5/Wq4oaeCPpG4
HEcGHlIoEuN+VfFgQCmwu7eC0JMxyyAd86Z+3Ld594PT/imr7foVYh7nV3lmxOJyd4okJag/lBuX
g7ZxMDu6U0REMaN+nNwlxE4jemzyTeYgTWj8J2w3E5bYjxel+pZ8KZaFRIB2udFRu8U2j6hjzJRk
5vPCcUi5DcZZw056Kq+yJ7RqKFi/qnpXTMoAgGvAZcXVlnwx52Z9RCCJo2vFZnY/LyotQIFr+yku
AwoJQtGaNgWTAVavVm8jiVbsMU+9x7BCsRirTOXmrho/g3mbS+f2UK/cOFXxm7JVfaFD2hQsFKC2
Hues0cgcKc1OcIo8tClbU+J6SRB7lhcYBvcNxhtNdiVXcpXHptSNgc42Jj0xtlhfuYSQmV/NO3Nu
ncXhmcNXSZ8uNNlV5mqAkHoL8fD2Mdno8AA1dct9OvGL9op4RwX40Hjc14GDp7OcS9DUoPFZk0lK
mOZ6TLHwZbSQd9Y3ZzITlfrtZJH+RRWhSq3tU/5dyeCwCqvaBf/L0CR4pO/VY3aRHn+HKx18KJoo
KuTLpw61RS4d68uoJFGan9dHsw//Is1sryv4uMp8w+IYPNkIQcAgR+jnB3NryOfQi+XVoGvFR5Zj
MpMkxUaUxFVdSdrDUSpVwqV32ugB8Bb2FyJ7XvygkAoIJBkFi0B+Hdv1fLr+AskDklh7F4j9bYfv
SRyDeKg58EY/2qIV945V4t3UKeODvqAgyhLtZyb86dBIRw8LoJo64cYXnATUXBD7QciqDr5P84T9
/DQZ2G7k6TxFaUcnPTq9qV56Pb63auQl/YiCXovGvqXCaoeL8ubKg737SuBCrKE6E1BqvLXyS3Kc
pVkccvJQKOWdT8Ohed3nuRgzXQPC5Htvhk2LsuVLoGHd67Pe8kZkfEUfQg08aw0Pq+Hm3eKsHVri
Mm1AadZH5nKKkydM4kIu2T9XVsv2uXNTw1aYwZzzrXb1dz3zQQh5MxshpFux01LAVJHzN4Pg/qYI
I+QwIS8VRd7B2BXvD4Hm4OuWtXn8sR8EBoUwmHoTYZbiwiT0Hzzd8xq75m4mc/4omM4P3pjyXMsU
ZpK8i+ZaumppC7X3CEjWk7NNtkelKZalzH9EPKs7FzLeBctgff/W1vqjw3g6l4sLIbtIvsLgy6yw
apDljqw1w14Z9rvv+YSJvciPc3nfWecHmCTZU+UFRKyvJUzAEs1RlA4ZJtdoCX21j3yk7J4gsCSZ
CIRQLSpqB5VtMxT5o34Zq1IytAVHW4jzH50vSh2mCdhKVLEKPtBBuF59aQBydeBsye5eKqgULQYZ
BXNa5XEYZKlh9avbTVj3ukSweUGJpIzh8RtuY3dem5tB4V4mPRrpMj5FfFoNe1QHCV5eKXls53fL
d8266BQc1/WeipddpqevS4SgINTFv7iB3oNLBW5C2tDiyYK82vq9ySGJDGMfTve4w65+ZuvItN3t
ip0QIOIA19ou72U3ScrGwLyFv2cqehTJoK0oLEGcYFoWTWxlmCxrMZFHxPqxCp9o7zPuZUFqgvuR
UXc11MxZLIIIBmnq2wofi2K2mPcmPQjbJDPey1WV3jGx8qTcAoKDHcPCf0QPpt+0bVBxc0dzjLHb
g5OwO/H0PsPVqBDQR1TDUymcGwZswQpyTZD6i8RXcfeUKS0JOj7d6c14S7uXiNpSn1A3BBPjtEeV
h/YcWZJKjBP8hico/38W9XJYkk8qCYqsNwdcASFJG26lkcslSN5rbf8pyNG5P8nKQFtumUtSP2jl
GsRhEz2W+9m4X3auPgekUoHv94h7flquCGTvV74GHYSpsSy4X13wnzeOn/Yb3hNxlrSEGVYZmSE8
Ags0EG79rMmx9NkJYukJPs7Q8wqTvk47kOuPLsuAD+1s2mh+DkBcuqoCaoW1IOqPMqsw7YHymOjl
ssN4Vmot+cnjGuA2ffOHjxswR8XSkqvbmWntiTxmTl5VDl3wWA3ZlUz/XvsSv1aW1fZ1d4cWWpRu
ZVrv2xCMcU3kEAibqx4lpFPN3BP/c1ciYXXbKaxfhzHDhLKXXOKvFIQ5USseWyA0d6ga6RmRjoYR
xZtu1RUbwGRxs/z216+ThyJvPiCbTCZivAMCI2Jg1FKiy5tZuIGTVNXxv0hEAuxuo+dG2hkFciUW
77zBaVUk67pFRbr3albgzU64LD+pCjN541TbV14uD2v70ZFfx446PqyFUhkb7dS1rBQmC2efcUOY
yulYJiZiiMKq07OCdG4ubdHEcFVKHHnXzVbIu9T8hkQ9ajz6ucN92z9Z/rskgXs+JqpcE2A222cE
HBNjdxrKhK0WUrhpwbxj7V/JkL954th+QSUycSRSnr1O5TicxYHiigaK5ps2dvjP2RA53vNcSOA6
LMtb/uL0efCFXNmwBfGHP1fgI9zUOv4PQlmN+n5d1ksl9BzhYU7xrxU6nHVj/u8oKy+Uni890VVf
+826PYzDRgyAuwwV+qWHPAUaMD2q4bPfJyFJm3BgczRevzaaq+ffRTLzqRnsmnjYBysmC+Wqit/f
siIJSRLeOI9LobgEKS8ul5VuLgEoFHV9dS33R4ai693G2NHszZsn41DLdRvZ/9/4SC4X1TWML3zh
Ozy7Mb3eMvui6fe5Tg7TXqDzVpmlETyOfwI34ZV8ZviUqSxjEVs5sqY/6xUkEfLLvQy993VH4KO6
4ZRTn7N3TnwZK4cQXvrrzWz18BRKmlrEKIEVw3Kqrnk9NmszMFIx26OAHJGG/debNbBQVRL3BFFJ
JH6Lg79mdlw4550QyKihKTAXBoq6XrmnsmDqfwANBGy8EH9sZ0m2h/wMQ7/uQWQHr7gAHgSgouNq
27Xnh/GOGBXGlFxtux4HZC3LBGMegDZUf/Nm5uQR/SPyBJP4SITq6apEH9Zl9uKQF4ar6yC83RGS
nTO8w36Dyg6lW8gd4YR8U9gWgoM7iUH5krJFhjJaw2QKdyBayd+cbfN4tLCP8qkPVmMUiFbSq3Xh
E74xVhSlR4wldIlZ9qxddcryOLcWu9KjXSj7+xqNJn0oGxfFw1VAc0ExB4lAodHOct96GWGTOwjO
kGqBQndNdX9eknQdOIN7E89lBhGrb9eMcDP+zFi7KiSs8P/Nlz4oiqCmFKk4n7N42QLflotnBTgF
RfbSBSJScrHMU+lgfaRcv9E9V0DB/uwcUpSi/Wp0exymPKgz4IqvH40eDOZ/yiSL9oVnFRJ1CyYd
IEltpbIqw2cvhYpkw7+HdJmNwnGdzV7zKgoFkSr/PRL/9RDd1XNKDdftjla2OhhpbLNFArmTYDwp
45piYlsZRZuuNCZ5uWaCnV9/FZL5rNZrzJ5v9NnHNACvLkaQUILphCUIvYTG6gQlJFgbWvGqsXBk
/voiQuWy+ZOvjKJzpW1hbIlfHz+/reH1j3qm80rJH7LysgnMD/ptJ6Op/e0D3DFyuJkVBJ4+TeRW
GccHO5kEoqkOYvOYics682v55MQFZLNgefOYMWLB3pJmW2ttw/fVp0m/ZGIwLEz1rMzhYXtAU2w8
Kk3gu7Sgf3j9eDEdnNbVQ98rhfa/1ePM9h82bxSP0yhvQ+GB9w0SFXHg4EJB3ncnEhC6O4pgOjkQ
HfThnPG4AB5GQRKQqrR9am+UTSfCCmINtPNSZvssihIOdLuhyakLeWyt+ET/12QtEBJYAnDlffGE
uI8XnJl4MGCRW92OHqnbfZyvTDiBEaeS8PwoIgQ1VlGxzgoARTmn2QQHsuiu50UP/kh/1+pdVU1Z
8j9kf3SMh4D4FMPRlFfZuI+YpUHfrCMPDgB3OS+m9T0hxh/amL3DVL7BozJIs3I3Y5Coh627mzeu
1tpjCTVS4G1rxmFlyG1daCYXhWTWTrxN7vDdz+jUfDgh6zD9/745kxnaW3Xfer0aYusc/D3BAaNE
fv+jtpo9Ib58PJLlOop/IfvQwcnA5X1wW5w6EvUE9FUTU+vIPeQfUn6mEa+/UOC4KzLvNdKUDhnc
IfbvNfZwZ0M+VeGFnVXXsnAkHXncN9wUpTdEuH9HbdAnnAC/dpYKlk62E5HNAzJH2ze0DuEamgwh
ceizS3MOrrP8k7nmdxr9Z/mOXf5zxdHcC3/7xDwI6PnYNJRQzXMfI0M6SVZZK/DBL6M/V7LOIXdL
XRqFzgdJlZ5hUv9kE/kwmKk82EZNx3PEUzt5Lcgt/FewadfeTyzr5gAp5wkLj2PUh/CW94PgiKr3
eg/Q3BEzC5iKVKQyO18J8Hi/89f3A4cndK2utLltkSmSHM7/GRQbDL5bUavW29ydzljqTEx1BNp5
Cz9gMsabuum+SGxv5BLEX1ltCn3ACCJdr281A4vUez11wx3GGB23AyaBL1joPRuOo1t9mvgmIKfc
CUFyq6An9MD0XCZ/jEFWeZLGZ06GvUO0iZyAMBSTV2+RMm+f46JJAcWcBUb0Q1g/1a6lOWaUIKRG
lZldH4QFdpEpuekxRLoXD7J0/+ByW0xjxO3xeAf7YLfmnQl02nZAIWEXTVNVbH+oyc886+4u24Yy
v9FCYTFH3lhmDopMAn8Wxo2CPsbOFOKB3plTSfKufVsWg52WpS8llPbIkqScFz/Ay0Gfc4hZPIpU
83QRI8xJF1lcfg+nsA2QgmMGfoNp0RTRXXSpwr86TSYYUbbEJ1K+GFmu2feJ8vuj/YOi9QNmv2cR
Bhj9IWtYBOnNmUcvQHX97oKhRKXUOfN77h9CIjP8KSdr5iPqgNgqZuwjE+E0XTCEad4svNXLKG2m
muUA12B6wVvoqGWleXQINCeLxzZwOxVc8NCLSoT+BX3aXS6oBGVWvR8tkkOozv94ObDWICib2Ei3
8V3Al9RrP5TCFsQSqt8whfNi+g2qYuVU61kEfJqgR8oaYMQhskDwpSzGX1s+wSF0MoSmHp97Ql8S
PUTdqSR+tMtVeGv0GuF25AVTQ0Z882xwlowTaZNuyzA3YEAKnAvwNMF4OehdUp+Fly2f9w9q4DTY
ok3cye/PQiYNVReswu/RJm2kyKCX2icqjhE4r1G9f/VycMOjK/clkNwIlaoJ2m39ztyyX0pYtTyX
vVubh+oouM+sdBkSuwLwESEIiLmjPK0jTTPNVT1mhfgltwngVITxsJHz91taAvXldc88SU6qFeOZ
cabOsf7k0ElR4vXQTPzaQFUN0p9eWzsZIPuCvaSL0zvVGhJtBm5TJyVzf0luvowh5G7IaBE72cdK
k4muMGrPWxUHh3dXtOZt2nYM2tmxTuqRwJhWzlE0pBm46O7Vo+E9hwfua163g4sPiigQMtkNeASs
++7UFNdxwCEL13nx4PAV8nCLhKUbcKIY/o388KUPRWXpUp/8tbTwz7okqONmP0eKn6zJzdxhKrjl
506clom87IDS8zzYb0EUVN7wyaBiVcaV2gikyVXDRSpO6D6/10C3Q+DQBCk+eo2yvfI1F2a2rybc
FCuRZNOahP6MQEUbxK0QiYaZ/lmqe9sHeaLS/MX+kKSlkBAkyGDegAqbt+36U1wE1EDu2KDkRKrq
rE55kyGaM3aDYXtyXn7o9QmwtjAivp7P1cy4p0edNHGWZy4EaC65J9K98I5RrpCygoAN2phtKmsy
j6IO0en4oe1TaHMIALrVHBhdWI/MMBHak0lu5AjdKsDrQZbHlgYWoNjP8MPqat5dlAmAPZZoc+TH
QbhbnvpKJcED+vVT+6RbhySUxjqAMIKdwDBBbyYLfFo1OaOC5Mg0WoDsnfCaU5MD7LAW5LysgXS4
YjPjm86agVhpHvKhRcaaVO/AYsC4NuCbZaBfmPFU6PWZqrKkRe6ECN7mJ1Bh1qgrDrjcsTvYt5cB
GS5RsEr37ar0CIg4sqKkFrK3nzau5CcZBYnmCCYGs5S54woBp/4c66RgWIpdHWhitlMeYaZP72Kv
j3u7PFYN2M7EqviIoR1/7Tn7y5Em9F9lKKZciOdVWo/WF6wvM9totWNJpR7T7auAbOWDdxqMPWWy
P3tswYal+z+73Zrkky7RLjgemx+YFih4lIIAFkaTfV08whVpejm0rCx61UqHsiVSn/NhWMSo8YqO
xJaBFBYNYzKvlS6XsYCFJiodT4oWnlPl9oaj2skPcxzbVZTc/fAQZlBcnIQQsiKqJrDy4+gKnjA/
2gM5szZw9nZg/W1RHWO2qXbxCvdTm3oQzrTYOn+1cGMs/mICbIG8ehSbDJ8DJRZlBfnAGeBjWZLj
mo1Vdal8hKgQaJtBvpIFGcGmUGzkZtEJqkIGSIeBgfO6OzCGLrNrdyphqQ3tBjbWN1lrhex2H89y
fB9oJtqhpAuwsYKB6vfZ5qh+HPnk3/hU8/y1HGNkt8goM0+2rvAUYPZEBqVUXbJv2piFi3mUD/mp
TVM2ljW49MyFEVtjCaIEliWhIgVsnkkivxlRynR19V2vfpL4PUuVRQH5u+FTNcJwKSWpnUdNlO3t
lqVMmxr1FmPd8DNGl86636ZMfzYAzzcSfvwOhZa/t+jhoG/kLZIGJHJsVkX91u/74UkZmefohLkB
TxlMt+w+MV6ZGc64kWEHFlH7hDE8BAOX8kmRB2rADtIr5zCZJUDMlnQF2EzkLLOfuUs3fQuU9049
UYhzN4GztlBt2pWS7MHLKV6Ki+X3dFPHQzQ3asZTEZiIHXaDV+8bJaqxTn1VP2OAAYicK78wvEW2
hCwNPS067TD64T8JIdcyFjdQe3T6Ct14QeSmQjnUXYY0dlhcyUZOihYU2FcfpO8wx3H5gEMb7huk
t++iGCcyUiirLpdtLg4nrkELxzlmSP6AUnAjW0Dh3UZ3liEZfpJqLhWPsk2y+CEuiFmh3ijA/tLp
llt69GbzFnBaLhppVwRcBHK2ZX9j5CeVpPhrOl8MqGmbkICG7y3cx0ZLNnFcPsf3d9s9w23H++eQ
hr+vhtsahvw2KALBue+aouxevsuc86N0ttr8++N+IQ2E35y6Qqs7fUQyggh5h5Qs+2CtqVHzZJ8+
R2rEuGPoG5TQYM1JeiCmg14XiPJdJG7AXWxkCYlbXYZYyQWcPmurYLmUULyINwUZd9s7v3/1GAbO
hnH7DrdAe2LUF3i+zdAzqk/0IR9jo0EDX5tjskyyK3AVSvfxWkk+eJuM1jQyImEOoJhYPxx9wNU9
n1sNAm1rO7jAY72LZ4BlUFfcasZkRoxz1a736UCTkF/OYN3HB8Jc8tjWbnnCRVsnV5ukPrCcdw+J
oy/yDQCdW1XDeH+p+vcT+rphYHVOUusTBf9+YyxFYKdmVgn4Ma8HKT9ATVHBpDTJfqdJ4kZW1Vav
/jaeN5s9Cmf+wubYmZPXt8TNnnTn5hj/4R6Foq6LT62yvF8RTd7lDeR3Qx7RK3BzPcvN71MQBaC9
2Ke7OrYR8Jj0QymAZDmKu+/lmy3vvTEi9+SpTXsBQUTh6MrobAnVe6LGp1D46rwPMrgDbNjHMAjA
Jd/fui2x+q+hhjxU5pf6xD4bKceS6B6yZqKVQmWQrJdQmi5msTvADIyP1W+zTpJBsxH1mSu/AFHn
0DDrJCZ/eweTUXxsrUHnppS4gnmO0Hioew65UDqDZBU8TwnOQxbbrcSAtA53bfQ12vjYNJYz5ECi
sfNcrU0H0xu9S8OsabWl4p05qTWydkKbVyWmGftGYheLKuRP9ZdCuRCTAj46ZaMgeIc3u/2Ss1AJ
CqKXXT2Eqqg021/K3USfxEsvc1GfknkE+aPioqnlal/A0n7MBZuEKoK3xKqftq5ZJ+HMRI8H9+r+
ILy6plj0DdE60SfWQ3vas9UB9f7DmdXI9RiA5LZWPZ+o7PNeAiTsgk6GfzmYgpYYMrsTS2bP2EWK
0madYVT4bxXHAg6/5aKRFqghxRzIfgJ8LkoeMEAkKK75Eg6NfdUfNvycHVDJMs3D5X43v/77WtN5
PthcX9x6o7EcsR4Y5P438ce1RLMgoKtPUCYI3mGBUKYm6XZb5lNB1ltE8YPxo/cWJwW0EgsKjFXm
QBBe/C+Jyoyn+orWPtDD2/PKbbNxZm7NJYrehej7/8g2GTmn6lniMTyr1BzT9h3uZAZYVd8BpyaI
6ROZGnpEE4RTxF70hGY/8aXqm/E3h8li+wk6buA3eJZrTGymxn4zQY/wjAeWZnPt9rCbCwicAU+o
8+ioW6v8T4LIOEF8znSoO9nIZkWFQ3+l6L9rNsp7ZzUTma6dmKseuRFDMKhCFJ1gWkjShfuKEgX2
N7I30Kjplbw55pBwvclyt9QUbMlcRyLu+orTYHzQPkZ20eCqXiHz3m7U60kXgsHp02fiqhh4F+Kx
ljGhxYjPC/smVPjp6YzhP4E5thGST1q+uMh0sFCYfyDSbC5qQ1EttQwQxozggS4ZaRgWpy0yDvHH
i8kf5BkpsmBjdZUL3TOWz8AUjX391U2gBhPMV++ospCWuIiV40ytngOWIC9A1g/95/ofOybCooLm
yK3FJDxfC+z+aIRtg9i+BOuGU2UXhKST0CYClPtRkxkDzV0+3bvjRHQfMX8j1sZqaGxe7e0xmhvP
QBlD3HzSgV/9tk+mo22f6YzvaqrpWq6hD7jcZoacPhHfNbPj+SRX09sZ7mx/jj2rZpdCYdsirSPF
mu1jJZl+z8SWZ96eiQctDjBCdiY09FQRthj5l5Wy3iOxYC96Ce3tm3QPBSB4thuHhDMMsO29jojS
LcVm0M+2kQ/S4grYaDcWzZwt6VJ0hAnLRvla94ON0oRRxmBXKkYl+3+7CESOLEMBt417FtKsUNE+
nsR893oKq9FPnhYtpUYDmmoGk1VV2oEbFONHzdzEKO0mCTvgy6RLqGiYO+2edDg5372qkIcrOnds
bEH/iI2+Lxw749Bi0FswsEyyezFVxaNFiJgPIovFCNLOLg9rigt2e3l11sySY3jC5pQNYAbORi24
+ztvlU1pylZ6M8ZJRisvqvQV1K28DVh+urNLV+rakUmVwkMOc0CGaH1mR3Z+9wV8fvOrgvi5oyhQ
rB5YDHQTQEES1ctjG+R4kYe/OELQVWTm+GOWbrsDAJxTyG1wPLiZ77iKAg4gip7i4Z1g0+QMREUu
12Mdvq4yo6ywsIIvVAd44CZpvb1D9pRNOj0nKkfez4SCetFgQs/Zlwi4m7syQlfftGHVEw9nY3yG
jMQhRnotQlfZFfLK3Fqq14ciHJysZ0wZa/bnC8HH7HMEvK4EBUJyG/QhgzcBPV8LhM+00C0mwOO9
606RtUSiDrRlj8xUbqpsn57pA1F3fUev6kyRjTdLfZQiHZaFhv7+fvOkd8rQArlwuYNOAxh2ggZC
hetSxgoUPG2D247KbIqmHQQ01NQOb7qMKftOHh2ojcdtJ4xTuI3M1Jkc1JjyTjvcJIP+5mxZrV/Y
PH9ig8PSg6KEjy9vpozj23Fy8IYtlFvO4uGTAFZIDP5VU4O5BHfAAo0qitqXOV+dFLDGgMAkMtoA
lLiY7Ddv9x/SlumE5wccOhgQ44kb8T2NJOgVSi5iYE2NYmawdAyRRfP+40owRrAYXbNtX1/Hc6kh
eFxwMSZUPEdATzleYlq4+mSDQ56y0LI27rMKck6czfYVmindIZq4F9NDULP10QfRbk2EpvNpL5c5
HrP2pNO/mJ5FGqUkyLQsqa66gSSQ63cMixS35AZTGIP3p6KeMV8xQ+jQ7UKLKkUoxWNQ3/Pp11Js
foTGSL4BY2Xtff7iQgN/ogWj32YYUruQZp0o0PA3scOLSEHa1rwEiF85M218EHYAWv1ciWv5c0Ge
u2pwqMIm4Ga17JvQxTCUV3eCs/INsvkxzvJ4UgxJBYUCQ3vuCijGlzU5fkRLpqJwBiIBX4y8f0pc
WFi4mB0XkUA4Fp5qg3SvlyTdC+WSHNMvpdlKAa+jOPxvaQepL7IEklaPc6OVN8up+KVNxeTw3/Vx
1LZFKKk5kG8/88TQH00i9fSdNE9t4IY1jh9kwUiqPXLorw7CBdAh7y1iMJxWHefqK/E075Vl/LLt
h4xyOJnBIfbalZEzgacHCrI7VARiIUvD0+sdzaexhlAN2iffeLIQO3MLLpd2gYqEOaySVwqxMPNv
xX1aM0Ih72SMSeg+c3G/4ozn51/Hv6En6aqV3A2C09nr0e0yFUaKDxlYeUl5lVLlcUr8QSkfpAjb
a4mCUliRtJ90vJrOJY3oR7yFnSlYAAOyM45S0J2Vf3x1ncAxsFlTaLnkMUmp0n5QkPWEqP/eJWgA
zEqDC1ROA6+KCHiA1jecLH5w/JpkF+/O8goODzfa0fl5bzobalRjTLeFIdXkWH1byTJ8RLsvPTKl
X/Id2NQOnMTKkNz/j20TIzQ0eK3Hr7ExgV9obzdUChgUPllDMba0NRKF7Xvz3KVBZchcw1VKJGzx
iDuvRcID9ql8j8lbs6Vl29c3FiF22+BQw8ZvkbnoXVjAtwG/r+UA5Qvm2GuBbFCo5WH9Xz6KgDu6
NzGef9tUEdh55uJFOweCJCWVe18/tkkLMCGhS57NaMhcmmGAnY/bv3xk0fuqjI7doTUamP1pRzQU
Z6fJTdx6BdW12YVJZeD+vvbKKr8XoPZyH1htWU0qP4PJ68Q9FXRS+70Rlx7o5E8jdiG7jFQAPKH2
8qkTXdNgO/7TyF6ngrpmLuUOQ6CmF7s2+QqkIEFn8S09TBXvf1ZmidZKZdYt5KSWDF1pSiTXLu/9
jg958yE+Kl0IVBvFPu+oyAcHn/VvtvlmDDQ7MZezqEnJkyFKaT8d8MSnflVn8c/ZgqfFUqxCT/gy
F1ab2tP7Zzg1CRfl22fVoUvC2D5FTIQdHATou+DgRGxLtCDBRcnX34FjrdskgGgVSEYdiGvE4DAf
ngBzd9u/ZcYbKoMXTFt2vbVwl/n2O0/O0g6V0TcFl8RitSiRs42OwQM1UAtVH6eTfc8g4NqFGxho
CP8Zznf7NCSbjQEy8YEW+Ebom8OTbl4oB6H/xfd1anCadNv4ZGGbfEuWx1gnN+PGqbkXA4GgsoEp
wTVZUfg4O0ljE2iIU1DeZa4yvW0P8bQuuCkdf5Jaac7xlYypMBTeYHtDLVIFc0PUzwqWyeFiu2tV
cg6Xxc2FUMcOVLcL0nP0C+umOUIUYpILtu+C0gjPX7dMwXovYZAm9WSwYl/XGsEctLvj4mJQhC9R
ygeFpnurDIlTEpdtpQ33yRerKoH5djIhEPFKBMmiUeRVejTEbiJ/i0W3NvGsJ/FaLwsf4gfmGKRg
T+0vKwzhDje2prm3HPKl448AEYklB2yufTaXNBOSkQ0fH67wXXteB1aS3/sK6EvVA4RK5+Ln/tQv
+SjsRD+AyCNJXzAGqZueYxEJDaxvJccSvBNeJVqsQsGaa5tCGX49dd2WVZnV0HsKW5J/ECZw9HD9
/hpwF+/o1olhD4J8aeMTBwLT55Bb9uDzwQgby7xz0yU35B8ZDOJ+3iQr+7IsISqq9mzjgLqrqBDQ
B/Q0qSJ6R+W/NQ6j339bjmOoGfdqNJ+mj/JuFrEP89FKmAtPEoTL6T76ny9zSxSkStSWv/s9pUfp
9m/LsEWI2zs/OM4dRBhCJJWHZgG/LsaCiZHr/9nyx0IdEo8tYtSPH4dcH4tmsP6vtg653TJ5UhKo
NngCwzxGORgODqfaw4o60q3o4ipO55pv49qe+WHDWD9kcMyr8cgj+8zdf18eclkPWHL6OQC/1qtr
GoDdzL+g7TYMoqDLGnXgI0syFmT5pfpT9ausa1z0Gq2NH0EH34RVDsnio3X0cM1PR2BXIg2A+75O
2FntbLbu/A50OC6d1vvogu7YXt1wmHaFsjJh/YV0MupEjXL97QPcV6lNnKPQJBzyagtLH439hpMU
3gsl/eYYcWtjXyuzaA9O5DkS8DB0u8Ob6fmufF5dPkZA2QW+fDaosEeS2ueMZdfnmV64TDqu+PDW
oeRRS5Si+eRa1xrupthjCl8INdA6javXibjgXBv0LLRbIgXkutwKlCFE+GvOlkTJnW91ZdrPJHXn
Va0S129+h0Ow0ZB07dQnQdQm0ZB14iLUUVLUX47aD+0gN7fv9eUXREdPcI7LGwQ+3s4/WsMnjmhu
snlQkQ7IfV4NCZf6OqQbMZyVyu2Z9ywApKKFNnRh2h8+CGxAMpMm4rygW1EQuxa+CY4PRb3gcwBg
B7p6CBdaJUnAYBATacjjKHbeh2oj9pmps0gZJPXkVQf/SsHhB/mDqAXTHyzjeMIIudvVmdpDwPCb
541lc2pnGlqdicpySrejiXfeaMpiwRD/dLBskjp0dEhl1Nv+loZWo8ojQeRH4Dc+LQsWKzy3sfm6
58VsRuwK9FY5rk3QuxdLnDvV5UQB49DD9MBdF7CAQ6anSUd9TOmyjXTjA8xvDHtrDZp/8yof2Ol2
V7mkU8IQqa422M7+skMQGW5hsxL822vrmFv3NogbRyeZMbgql97ALhrS1/nbPFgRaQepiFmZ3N0n
DuaZaMEypqtYnw2G6bjCvcRny+QZVku0jKsCM9J/t1tQ7bnpCTzDBid2+K9nAYzaNXLhba8NLwB4
irGanxxG4s93BYEUvhuH3z9EQSOLP7TnNPUDwzpDximPFX+CQguxdZYyWALAY7aFQtZ5b/9gSkYX
iqJ5E6njJ1N6ORK8DougV2CP1XS8QsDX84hu6nqqb40Es3D6NvJXL2807F3TCJwaU4lMWidebHMF
cCbTwYFeMaTyX2tcYBdwqSsxlNGpBFq1ZACUOJhFpm27KEJBOWHlh9DvjOXmQVjT+Lxw7XldhUd9
R1QCTJEFf91lCKBbAltAe65bYfxfh+nyNvgykOFc3sHNktimoo67tIDIsmDnhLouqmc2FM/f/8Pj
e4EVd5ja5dbDJbNOj7Qh7+IyEXFNi2PGE27Uw2ZEG/lflEyLRVSuckZOV538xFlbKBNy3xvsjjRu
+EQfnuy/rHP8XQOg9H/dvlVuog1m7CcJfiXTyFVLyRjZabO95Z0bshMqM3YZ+xvODsNlbD9Ly0mY
t2gUsGqihfx9IIfMEvkchhU7xGZ3J7mrJmL7Ef7cyHo4DITOVeJTFavzvntow2lLQmCSSOH3NjBT
GnqgPUrVi9UdA2c1ExveA9UU8muFoo8jvAmBgiybYD/WaJSSNh3cOaajzFNzQsPHeO28iDRuJqxV
5oyOIa1FWnM45Xl5m5AbE8wdsrQPM9Jj8rMzIS8wrp29cL8K768W7dB5JIBlSCa7VnkyJWaG2kEc
ERWYVpAW60VVu5LOqFoetccqNFEIQ80cxJPn7aOADt6wie9rANWvnwknFBLolaWmt6El4P4wnDaM
8AoDUwayqksrFBs73UrdCmruhW2VsGHR4YcQKsDRW511ynh4fJ1JJBROVr1K6aMTVrjyd1YAViTf
BHOTTUlSdiV0tS9rptjtvUnC0F8z1pKsQobm92JvWvMuH17dJWr3qQWarDZAbgrhxReUYul5Dzgy
79KcG29vIjsv7HAWFUyC8Oq5rkRnPyVGuG43RoZV+i+Q/SP7KHDK2KY6ZD2U5f60HnyR10l8vC6K
zHdYFx/HAapHxTJc9bwOKvsfxd9k1ybi87Pd8wEUT6j4xJTc1+2kA1JsqNmH0TEa9sBreOByBzhM
8YdhsCyxj6FAzoE/4Havwy1tsvJWzTLhXwwMQwRYETUPYd/wYsmoMMf7IC2nP8l4IHchT9bre+dw
8jYsbKIqP7fkfz31USOZwSrtVkhgpyVSXgk+qemT8uF7/SrigMQzwlGp1OPamFqKnV/LI+69v+dX
ULKUzsmT3tc+tQ3xmcv4cOSG628YlmtnIBr+TqCGNOO4jcd1IlTm2YfFmuRAL70vQdEVR9WvnF28
pUWIZ72JI4KYJ/DiJuzj4logojzE2uwlyZ9GyGIQq+mVWe/zPG/jloVD6SsieuBDdnhDeBwkA3xG
E7cq271x5AOJu+xrgGQn+DO/xV38BlHHRJCirbr5BauSPcWwpkPxYVeZ4Xo+Zz3ztwHoQaoTt1DJ
lSWlU9SgV1rywRll3VTRk/RoqMjJF5hO4GuTlKkWH6U9u6vXUjnuDs993puPwM0S2js1zmvkFRxA
WVw0jS8OXaUAEmuEJ2MaeAfMFWQqmA1vyzrgFgi0RrzD4E5DdcQWXYBo8CW8XNSl5FNpOs4iSC2X
s/pm2WRcrUbRO2w8eqLrjWCN0t79uzKIlSxz+/LZ9xNCBQlcj39+PYFj4CWUlpHPLF3PiYCv0vVd
1y/POlBvDIAbxWuZI5K2dRxirAw8TnFa+Rx67ynsDdnisfhTwRu6DURJ7cwbB/CAnlDK/tVC47bM
3UtLnGq/FlJJILtQDrE3vBGh4q23XshTs1YaSBRwyTejQlDK7rOPPanihV4B9K/tQUrMbZiTBkn9
b3eQTnAa+KoKqXywWmZv4KroMZXmQCarbh3QjcTJQu+vjOZfhZf9hfeK3NE0veteGahLpg9q87QY
NQ4GLoffY37RMVCQaVfc1moXyKRP2pkIcsygktl1JolOKP08pbZQPW/aIAjSKbmvVgGy92Cf5H2V
kEl0WrxZ/sE/tPiU40a6nUE0gv3q67ThF6dclW3GUZU4tSowMg69HnQmYbJjXRqXMDD+7DSRJIwb
raAvtfPTcdge+jL/bY1c2s/pT+fk2Rto9RwtYymG1LB34LnewUUt/DoXakaAgrRziBWfaUY/99I3
ekYPhkDm0U7RaBQJsnzAUQff0xJxslGKMQcXshaz5+j6Voz07V6azANprfOkNCrisbb/CeuzSFyh
3hLNGMbzz/lK5VA8y60MjGI2rwiEaOByOHl1+Nissz3xWVgvjTqwpcmINNsUq/5uXTJZv/g2VCyM
6Dfys2GIeKIU8Ip+evDkbMj/YBLjv4U3Yik+yiCgpIWbuhLRrgfxzd0P0PFMcLYnHT6cdl6Lpf82
VEczWBbIsHz217YOewyw4vDb6dWlTDOVXelMHQOCgqWaRV9tj7oJ/R8Uij+/LBk0e682O1CydKcP
Qr8lhk1z9xSZ7uIpDBRZZ/drM/4WufwtFxxL+rmfwKCTiskLUrRj4we46034HD9NzmLecdmscvq1
X/gbnAY4+LE5NQC4BebKfG6Prna1vPcuVc9NFoRjgHsD4l1fGzeYs30j6Ba/6ddsCLWmVMa2adzv
xSSNeMrCxWnEbH9kFFPwspAuI22zZU7u5gpiS0SMcVsnBXowVZmOm3ij/yKVYn2AoT3409gFHfow
VlOGztlJFwOYZKJSiFUO+SOsBcXvK+zo6pj0689yEussBRPnRAsQQvL1HVH4jPHSTxI0ZTTbcjBd
iytX6PSZg/Rw4+o/0QtNyQOPZ6zLILcT2Af9i+9R3b1CgpWtzkUPbYrCw750sUfvzOqizLCm5Rpn
OKZoUxF/mzfxMwLapcHFfARaix0eTdlP8zWgAHxS2MsEUBl/3VqBCIQpbZZ1sT6jhnGwiho3wgzT
1Wp+bubVQla6eGt2Ij2F6PtLJnY2hWcKOIczJ5sjKbop4UYDERpZhDnM283SqIogFM6eibruqWAq
VY+s0VQzl7ICk0bMvcho9n4V9walUegcyRY62u/t63vBRNRDauXWJDFnc/REnEMKDGlilrXpCBoL
N60eYl56ko5RlYebD/08PUL8Q6AHPukLwqJUgG+q3Zgpe2zdHGWyVBn1tR4MxMY2dIeMQjJLgEfT
L9AHTScp0evgMhkfmRjGrkhbkQKk/QESU/O3b0O5YF0357knAnh5WnOiBwqM2rpCTmRdjDqra99u
XTLhoVmaIa4A/m7fF8VruKBIk+y5XL//X+uduqBRnfc5zIL6/nFM7RZlEC9ZvKoj9I1tfr8PnKzk
TXUkpGmx0AAajWlAerRnfMr4Hc/hiO3abaSPk170ahee8CapLatep4r9MjxebBdYeN3pzU6jjPbb
SKKPcEyMjGJuyPcfeK6SSwvamY0ZWgVPrqdqtGcF+H+kGUHVs4ODaBZ0zKElMp6fuYl4mexKdjYJ
qGVyexaG3yd+w1dPqjIAVoEVcrfcnNuw4zQPdpt97iAx2nprCZEwChrcpwzP1uG2jHFwMYRxa/tt
glQGd3n4QOTpVT/0ChgAhv3I6XG9VQbMvMI3ISd9tNLme5Ki//u8RK+CiiOfbVZkvZbtqiMnlJdx
Ly7X9wYM4x0Jsl3T0TrkjLZvUIhKPGmTB3rVuPuS/HIDNpX/LefuoNmFPNbhAsWbmtvskCPZQeNb
XCY2l9b3Z0JHQCF4dK9EzDykJb7W+AffmtLGJ/Es/Xr+0skbsvdgGYdztrpfYkuqs/3nOtyFvL0M
iWI1B5qK+gf6ihnbKFqIuFV/GUSnNl57chUcXVn+prwpvwGk940NlwWrXy70TRl31Sx9nyKoQ8bx
OWC9Pc0Ik2o72/XUdiIDPe7L2TcJC3PzzdkbjYp9asD+cm3cXxWKQrNNzwLXylTVbvg3NClUs3ti
/UtnY3iOxvWSp+RgF3c5AdSXi0J371GxZ0cPhJsdWsKI4La/vHyEQxMMc8tbC8G2eIhIjyjlChjs
lolDe8fLj6fRMPsFQSZGk4qYqC2EZ4sUTgyJuaTxXYOrJ4VBx96U74gYWtSVk9loKN90kSwVLOOP
Nvo+5V6n5tBRrOX3CVsdzvxGZ6vYTReS6sp+HUAXZolR1NVsi+NxmsFWrjjSV4imo82jK9aRrAlG
E7GwM8Fck2M2SsGK6hmjTkTPpuqYKcCvk92+YMdl8zlwG8DCPqhvYBfPfMBJr1KnL29P+5RUOGO6
0v15OLwtuQCiqCfPSXAD8NYUyaL8k3I+Mem6WfW/jStTOM88Imvi+WvG/+8nEAsJ1Bu7pnVRqLDK
c5HtHFTzI0G6FL1pmAVSG9sdvN9rfszYrh/VXnawad9L1T2vo0dGfKzHlfCUBnbyZEmWxnbOc5/I
bnNPa//vaHYelAtnE+SSXnDNkR6DV1KGBYJQdPOvXnF6qiCz+wy0qwI0rECnur4S9CMi051vc9OZ
PDeO5GVfn+Crd80i7RQpTq2cUWws4hEqFE2+f45zEN/NPCvu1AJy8S+TTUGV4e5HN7VB37SMe6ZU
FvqYGGXJOxdUkBsTDHqYKbeuKxnijWyvW7SXc/lVwtgRRP9uUEvvpOXMfa1+pVbHh50nIWOWvUA7
Ute0/eDg3wxcFFkTH0xmJr79+Z0Km1H6eoRw34VNFH75SUKsQtndp3Jgn2jC0ZGmgWp2WhLvNvde
OgWB4ZDjKB/9jnpa4G04WSzkXg3iBXWqJkYESy5XaADtK/MV8Vos/ebRyGlwPAtq+ma7jmkA/l7e
QFOBbQX1Y2Ru6g4HYUCBaMjnsIt/r5zEsSgd3+xC3JtKMcDL8+rn0aSDHxFT8tHb0AV5h27LJ2Ir
pHYPnfYlsTu2tugDY25Y6iIzrYK2kHexBR46Ls9r3SAQm2zuLC814SlU3Gj+HdmoC9xL0nNXfwRX
ifM/wG24x7bugGT7NmzmP8Uml9qPsfo8Um/iiFgyDmNy7yE5V9Nl7voHtCyAi6hYqTB9kGqfp5Kb
4AglDlenIh7H3XiKI7V/QN8tBAl0beSwxOb8UYmNQOmTuNWq1OA2Q3mFkUSN63UJTgfXpQ10zM5K
wYlT4jVm/Lv5f/a+sSVV6Ypea8vg6vDLToWAi6MDulDLOnHLWIK4qoiI+ra8NeAYo1nCDVAbUtKk
lzw6A8QOQRy1lzw7uDQqZ9kRwZkMb8MF7n6guK1IELn8FSZvsFKO71LBd78c/uTxb/EcsxljyW2m
MzRi1vCS9QU7GKzR2lwpP6GbNKrJ6RwsEw6NdbJe+I2oaaIcI4D0A36M+rTvDELvl08NSuRvaDJd
0QfzP3ux/RLyrljIgSMwdsOfPKin1mWJTnMPVOmKIMn1l39i7gBRjGORBGfp8Sr009AOP1EldE89
4Yw4pjHFIHibT0zQfrIkjRczNGBMreDtSsyRb5G6Tn2et/6LMfSW2BcOx7hirKQdzT+JMerq44V9
cn8oqcvzIGy0SxAmOkHXQPV2tbh2L+c/qT83RsFJri+vvtKmrXvFCjJ3YdoYSF/9GXIyQ5G4mEr1
9o1Mi9GIrELYER1ID82Iadk1WwSVwgiN9Xd2BcbuovHBlcLqKgYaNYj74bcI5ao54Gq/PkGDJiM9
ZtyVLXHOUQj9HC2tLQ+tJwMQbomTihyrhEpWPXnnnsG6qeQbTcHD6V2UslSw0294bYWvME5gk8hd
Ftdam1qCy7tYv0naFqRmJt8sI03g2JdnobwgBxea/G2gJ1tZpMzb1cB2nDICMjAKaOENawvE8RZ1
WBgLLxp6Ed+w61i0FGNNjyEQ5MX03urWFeZcbbjQDBnAj6J//slwrzUjS92XFoSaVdgcQ2FdwLjo
yLXE40600XMsopjfbnQtvVDSicumPDht8AcsiETcaQ3ozuAm7ghHxFCuQ+qPt1dMX6YDahUeQek3
YXgNt+VMOhl4LD4NYqZGxL5/F/liYCUHJYq98RmnS1tRdCt3WGPesMXRB1M1N/shaK182YCnDg68
ggvSB7lZgYmMvgkFJbsUgs3vjN3/kGmhdtxr5gWI9GfkjgCnfGAcrKl7K+fgYXdZ9vOW3PdfhCb2
SfPOFHH7zGVdT9O2yns4f9z9yuuH3UrhTCoF5XRzXJ1Ut87hMiKlEahLC0eRcX1xrsO62U0VO8YT
fRVDlFhFOUYyAnLc7EbIjXNn1t1pFXgwwoC6Bk2qrj36hKzADJt05a0BWG17in9gxzEh/l8rGcmJ
unddOHwCn/8qXj5Lfo/Ol0b0r2W/ey6rle7tSOcGZGgFxkx2DcMdF1vjWAj2cRgIu6SSHKvoPSlj
0mM2m3zbMiRb7OXz3qD3ypjS972dZF/t/IPXwJqu8FRlFTCe7iG3vaf+jB6Q6yoGlb3XIQ0DwxnE
vJ8nkjv++ysgWhKOPrDE3gqqIVX6nwwebEbaGkfh0qqmMK4+OeO5hsZ/7Wy5Ax5IuEQgXhN19wy4
zmOtxtDimBqpKwTR6icUmFm2ZZQLEPdHG4f5g9vwEUW6An+cxXWyCXOauAvVL4NASUj+1x4DyfuL
HiVKFTD8fQctSGUKLErXM+GgMoxw6UeCoRRWr/x2C3p7ImA35MGNUjFY/TsNPDqS5f90sv9Wbige
eQtdsirz31v+yK3U/ZeY5wAxM2S5IQl6SMPIY94rdGf+i7WgN0xNYTH0fcGokFrmbQQ9VqVgsXUG
lxDBGJL8kzhD4gcGOvAO9nvRo0bv5+f4W2Z/Uem5xWqOVaKJh9O7LXDXsJrOo7iPaAQIaG1LikVC
IRSknI/nu7h87aWA9Hm76AJ79TTUCh852YqsFJmMD+YAD1gwKcAG9QxB9t9gzvEKnY2ywtKOUeW9
QDbzYThRtNlKOo510WKut3mDPfDtCKMHyGiCzzECvw91wfx/qALH/qqIedKxxxnFgvVGOVUYuGlr
fNAXDC3BuBapruFPfDMcEpY+eJc6ZksdspL10PyAQcH7BFf0Iec4XZT/mwulvxPhIRY0RF8ptEkE
wFZQR4hLzhOhOKvk7DXPTmNkeifBOKSnemfpdcG/+npYg39MkJ9VOGol5Z51+FLb49WrXQQ0SfsS
9/iQi7mof8PhM6Ogd32cRBFs0dkHObJqJUmiP1vPgH6PB/N/yxZGma+O8p8nEN2Dx9DYKr3e88cl
bRp8V5mLQaz6iRNyckvReheC07vOG1YRS6a0XQWa7ziwHXUb3uom3QcVtt7Tqy0sH40v4RRQLH9b
J6v+4DZaP+LIVgt2q4UVtbyVnfQe5DRbYZlYg43mPPRykuF1mfAb7nBeyKZI7QOfNVAdmwF8HTdp
nywMtr5YJUfGMIju/frCygZ0Ql00pBVgOMovZq2vgB3k3+Za9pcYhMqas1z2GEwCSruNQ0nhU8pf
rK89yhwphNSUSnRItml3WC/EK0+ANrPKR9KTY6WQtFXiUvzRdmlpmGREQiQFvfMwQWd2Zecz53LY
6otiEvkYdQqfWhplnRyN9MO55fse18auTPuoaECTBOyGjxw2JnpAVAqQNl9Usn4y6iFaaFF5VCN+
wB/XAvwkOgrq6YdiHzVuLpDJQ/nQgDkx4cWMXjQSEXVOb9XIDrtDL1ZcYp57iAZJdK6OpaJTUMHF
m5Mo8/lxBTElYY94b4aBjAr+jpzINs0nzNTjzy8R8r90vY3/rK2i1y6cpCjVa1l4egmVX1GHoY1m
FeV0sTxwGiYZ6ji/90q3z5o8J6nXEMdx8fUVxd1EFJN0uWkggQTzDAC9uNe0jMxQ72BlB5dyQp/r
xrfKgO9nNpK32hvxyOL1mMbhdyfd0KlvKAYt5FA7sqCYtkNnTruOwcfRaaPfJbIHOfbQQ5nDXNXb
Tz+ZyuCvCj6ZsNFIfyFMvQu8oUa5WKgslKEg24rPlsLnnoWVx192m9s5gEm2UqIQZg/XhG/RKT19
XmxFm1yH0SpifUyGL1MU7VXj0KdyAVcUGuIT0zIXW6a6mkLS6iTYDbJkbubG8hrHJj8Z+yIRaY8Q
bPOD/AgdyJPsGrrX0NaL/QXg7Dt1/r1+luArG73Ls2Ltmd5KcPQ5HVTZdXnmeHBDsZq5DfN1mBpz
ol+nd9UUqPvF09pgDSnplJA5gTKXE26fxrZgGTq+Tndjd6ExM38MvQkAxMaJi2dPUxpSsL90A0wY
oQvC2LEnaRC9BYiB+N/DiunejOgPAnpg91mr8v5T/xgCwZiebjE7aXR2W7+hpAnlA72Wvoau5MsN
njr09LpJOZQPYHHIfQATYaIZOVbd/IBveyAAHKXVhSq93DD+DbhHUWd8mOC3LSc6fmWQ02jXlL8u
/29DuMjvzO6TY6VgZtV0e9wwKzvjELI06sYeriP0J3dSc74HDZ4Fjl4W3NNhsn8jlqVbV/0k5LPS
FzaNP/pRCCA4/A9FJrLWcxk7YrJM/Y0FgYqDaxrMElVSjO/SdVxcv38g+wK51S9FE+27LO6wB3Px
gsmIL6kc1Z89vkYGzk8KYbYcasY4C5OTWFZWMNa0DSZAlWkBcVWs8JQNeqQLmCajA0BfX8Ffd24g
FKsGI0YuIL48X1UdDNmtDFO2F9LeUKBj2EKnxqA11etbiYYYV5eSrKCIqKvbIGnZjDwOEgJ/edkM
kxr0I951GPC8SwH24Rv4kyvjkS1NgffIoD7Qoys2dK/HHWmeBAi+d9A2rbyn1zpgEsNB6roPXemt
zJIt3YeY5pkuj9ZwbvWwfCFHln4XIhbegG9ClMg2mR1ambG+hLbrwExs0AToXr/jZa0Q+oZ4IvA7
5GkU4t84DUhcMcgkxtCsLHjaO4xIcmWJOwyGmnxwwbRRFrUFvFZ4uh8dge6dJqnO+87jBsuq8Yd8
VLTCHW4pVtxFZAV8Up2hGniLF53aXNXUkQ2yWS2MUmHvJazO5YK2kN7ELceliZgtWamRFwDKPqFC
VeBHYgUUhq+JuH88+cvdgrd19c/m5RUT+YObyB1nP2KE8fM808qLIVlUvsE2q5HfaODxr2K9QUwd
gYbJbNmyV3HUvYH5NIRJln4SQ4U/8JDHGsZQi4tcWZJHZ8bS7gUZAIaNuXfDRqPvkDMxvI6H2PKh
+LCP3ONfm1KM17l36KcH5xyq/yOHH7qRcTb3m3n2lAi3JxAfVp642t9LoNUvLW1Ck1VUDzZCgymY
aOZRYN9mSGO80ZTfaE1PMISMi5sQTOmSeUA/EVtJZl+uGJ2Tzay/G6ph9nmur2QWBRcXc1pwKU4V
m78Ac/g8VN/41AcsAJ2rLUKorn7Wlc14a0OIfM/ugXdkF0kahnpg0iRXYXr6W5oCwfH54Z54h/MY
IMtXkFkYMQ2pIQDR34WxN6uqB6r9Mc/+CxmkSJzEHUX+m5rULWFtWFNPsQEqWzp+1rJWYbbutvMU
HvZmQme76CdxcE8iHD+RSdHKMF6m64awpxhEF91vFqeTB3RlNVVNl3i11dq+gvmmPCQoA7rKMBfS
tvzTGLggbqapf8/Iw++jF+uf20PuZGdN2dxMkHqdIGrsjE99DbVFFVeSzcHp1uCcMLHKTfgtMHeu
6EwNLRRds3rrf9Cyr6QPjJ2Cd8VBPsx8QHZnF770EyLrjMzVGUH5UqrbtV39FUeKUKZ+snsCeC4Z
WBO7ppDLLrZkMib+VksVUO7U7zwEHoSi+reK2SMtzfMLzKKCmeOwbjj/n6HvywHSZCQIVvN7LNAb
6neAzK5OECMfQMpa7qTWpSwNDB3bBsUhVhEdUSJxyi58KnJXSr5WB5nxLX/u6UqhX4jkDK/NHctv
6n9T/citgAn61Hd5T4sh/AYkCBA+N73RJx1dtCO0ThhdbVBEesrZZe2hQ4/n6am0ZHthAKEBBFeE
VqhISSzBJXFEOCFVflJU2HTeqC5GavGirQBdLfRQa+7qpnlm3UittAC+2c0CfSp4DOpT8ZQehziI
/T8l10bwt5Qxk82S9pwY57KnlLGUzw238bDhDB84AilDMk/L8iqCwswaNwyKF4cU19aD/QhJNIVT
iWRUq422LoH1b9h2U3EPJy4COwTV+9bFoQakiuoRU3KtTs6nEhBEp9PhXzCy3VvmnZNfEVb4+S0J
8NmtABmsKlc79je3PfosHbTRwYL3Dn7hxqLWOyYQS096YVfUzAV65UC1br6C1ywzm6tDuZhWBt6z
fOrcnbx9hRsmn23uxV+wzirbWUnJZOGHX89h46Kmufc+z/zSdTw236PbGGaQTG03iz9t9Fc4dVqD
zIEseb1eRG246xTnFRxv0h11eAB/ZHEgzT2iNkzfozJSkRZpAO/WyNsRlinXuHY8AFp0qtNzm9sf
nfpS7NjS1w1sfo+yKLhxk5XeXONs9y7uLQ/RSxNPfCb6jUQQrS0OicKqCoBw/jZGWXU2n+RvWP2F
oTQSqhRNkedsGZj57Iw2og6fCU3dvzfB6EL1xJ8aLBdqVHzIZK5WkttGOEC3z6IIgQ4WqpV/mLrK
azjMPnK0IicDmQ8ie1raxhL7OjZpWvsJqnJmcNzzNT8U/v+YjkTWWGR6N6AYxRrMt94oHQPkYb2E
5xLsvwFb8ejmRVUgqOHrPd8BwCKk2xrK+2iaSa1Uk7aP/qIX3Xj3OLmFXJiiXHevKaSzQbr8cO8p
XfsWJNrJdSP7Mo9aKEzdz2ERVo/oZucIH5xM9td92/VL5TXYyjEBU1nbP8s9FR9XqkuttAWEheOt
MBRZ8jQe1eZrTctOsATwRHcQm8v/b3bshaHKUVwgNHz4iX5R2woNHFwxWd47HwIOXjrCcYCf7qgm
fl2PYk3ZTh9ELQMkGfTguD/b7uihCsIQ7W4E3c/TieQw9Mr77Gst1wo1eYzMNDHhuuYw5+N54Vyb
a3oMgoKex8XYHQlAUjo4vKEgTsyzjkXfyojYwtI2kkT020sWL6CHaEfpYNDLS002vZGTR1990AyY
b2WLSmAsVu/Q+Je2IaxzjGtPvaKikuYKRU1i4IhNysoncBKhb8N/rQ+PqygtxH7gKTA/8ZfLkuMM
5OnOg6OllK1DNsCDamILF4LLaUmCaKAW/i/1o23jeF81/EVEaIaEVj4Fl1Yz+p3sMrzzpoBVjGFg
oC1gp/PxH/A3J/tTTnb+uJSydjbX/ChhzoUYQ5hfenKFTHGQHQpRSdhsJf9qSatylvv6rUDZLID6
gzwk5viv77Hcums0SdDEa2Q9JfVO8N2t5A417r62O+j/1Ne2DrndM3MMNm/febp2A+nWXvkcw4KP
XVlDpciZze+YfZ6Dq4Q+c6aWeSE/ex7GKaYcUrxEPIX+lQ38/SpMY8fAaNyM6C/r3NOmYjpsQ+Pz
mmL8C1iJRjWfW46No4WMK3Rc4egK4ksGsft9h9j74Jf1yfAV2ui/WxhHFhI5xcWGy/br288bQQU+
94A+TUmoHVzB8EvWskhC+GvayjhuO/5th7Cqygfr/twmCVVLMnxWQJgn8EbsBahl/kqv6JsL1Nmm
dsC9LLx/lSA8FFgmGlqPu+G1kF1VM7LMmB2pGEFfWIrhJYCOh/3tf1Gmjv/n9yGgpGUqb7Auf+dA
dalguzbdaKtDqPSFIU7YbVm5Xc4Fcj7BzYII3lqkUZasjiOlwU70k0gWjd3hd+pFZi6yHaEusLua
WkiaMKCXBC0AmA53gQh4KxIa5yWdfOG+UHRPRIdxsvMtXU/w31yG9q7bgv+7w4RI8j4zTBVIUJjd
bWEYk1cg28tRnfFeY0LsXNClb7BDZjywlUbuQldRfMGh1zv/O5ouZ5zMW/QGKXZ4xqRx/GrmQii9
KDq8Y1OKIZXZmO9w3Oq//L2kJgANIw5GFDtfCfLcZNMtQ8OW9H4WPzvQBFM9iDEw4fJirZADDlHS
dT1X+8/8LUjbYQe+J5g9ce+ygF/1jgfhxveB+Rq+lejAbV10kIET+5ktKV7sW2mk84M/NWSEQn0S
Ow7JPnsHlsRuuql7puBKAOcHUZKGGXMjsjr8q9qc6liY+DanB8gmeAscqqQKqe14nsRdXKrc3for
Aj4s8YhorOqpVBvzwTYOTCGLaeVJojn9guyR/c6bPKyve/i1Xfy8oMeHG8HGbugGzRb9/iGyGwqO
FpLNxYz+lqIo2xPSLI3i8V8Vk6eMpQaX9dASuGSUUx0Op3h4+cV9TaQ2hV7tq0m+qSKvRqct0XwZ
7zYLer1Kuzj1V/tJ4/5J6MV/uL1mfr7wRH+DSP49XId4h900LWiDNjX9qVw2bzYt9QoAMKrnJIcL
+4h71CskHiACbziQ8lZE/WW+omDH2gRRqC45fb200sxQSO1JooA9l6xY6RXe3eaAD96Hshg9gnKU
hwQ1ED1yAKqg1O0HyCLsF+61x8wl2/yETvh94NTTjiSGrUJTtncc2VAo/w0FTQ2lnJZkNFpEIpr3
Ca0+xIZ0Bnb+PwbB4eSHdblV42dKwjzeUahWu+LU0lfahssEuO9IHx04FXtX/FvnFaSrXRl3DzGU
oCwB9nC4HMjPrlKSF7C51aCFCWVQvPWr5hQFVChBYVoAi6Z4fEF7uDzIKG7MIKivWnKF6+56fpbV
O3k2vJhLh9ZLkB7thADGFlCboAVmEjV1+z5NlT9gjMtH0ZAfEPRFVIUrNbXTPUdBoCZcp1FcLAj5
7CE3qcRldGfrjGPxFyB5z7NpT4u4O/teonVZorsbOImA3MHa63f+9dy3pYqRza3gjSspzD2/9VGw
D/SKPgXTjlyx5BVtP3CqS56GJIaWfLU1ViLje/mzXMWF20WnFxiyTyda0LjHdYJByVER6rvpv1Pe
0IzVZYfA7R4tebdjD8NI5oalybIwXxg/vRVKUbZkgRPPDUNNpecS7l/iTW9P/yomiiNRn2OxPwNn
/Bde6+7EHy9WxEqV60PIlx9z9bjRkDaVFLSZf3tXyO10AEQAznibTWeDIoQ6gmou0k5OI1zQe8nX
UyitJmaAaYGrQxZhTYn84aeInly003CikfC1h6zWdDjn6THQ2ZrHpqEABSlor4zilnzDT9KC9LIs
F/VKbamArzu6A5gpKCPRr7efk/bu0a70FBti9JFhrUMUsWR1BS3w3Vjj53etcv+eN2JyTkNNi+cy
4l4WaFN1DGYrs2+7JV2Hv9wv52yRE6nmtuwgZxxAZsAbjLCmwnxa4SZmOPGfET5MGM8oURBJSqJn
0VPSAtmgtij4zxZ1CdOUOBAQFdfTIT4L5Vd95kaDtgQqeAh0uRWYJq2K6cE68L8uADMEgqwg+WX2
hgjKrF2fYRyLPY1w5VMNESzZrWMsw+DFtYmLznrCdF+pZHYcwbbaz1GiLYjRnuHJq13tZFv8ZoqU
S4j5DW0TbWBHP75bAdZs9gEodKwYKGwMu5THOY5sSIiZLawH1l/nXuNMhelK80C7HqqTmedWgQxz
Lg7fzwKkxLtHjCPvNE+rv/7vgMqKvQGlmAQlqiJBZ6gU4LklegjOdeaYmnBj9BgxUds5v0Pi+/lH
2OHUKY0UvUpyqJ4WQmN4raCneiZ0jqJk8aJDbPWzpX82qMHXE4e/wm/PWUmudlEntSQnSnrqAt4q
Ip6rMKeOz7MEc3Gn5jY9J5VBD2kUO2t6sOYLHRp4+HRq2ZZM7zTDoW2sJz3pXSDHSO+rWz1N4gjp
I4kpplUmzM8jQ/n33gRYaL788q5oP+kaQCncdIRZeoySnbC9YOqQRN4GkDX4TwmiKQOTd0rROU1R
n2dsLAFXdWDISrZNUCorHHjQB+9Yq+9GhlDN+IbG64luYuH8v4E3Q82iAKQwQCexj7EEW2OAP3n/
UiRvfiUzeMGYm+hOaZUuXZwi4pxmm9S83Vmct0jp/CRwsdc2i44J5g7LHtmAlvKxrXzDvH2PqN76
LvAhhPoyMdSlvSjOlTQYRYtpQ8KLXit9h+h435KI0zx2SZmyr7/WXwYMH8B5672vhHiAeUPoM7gH
Ezw9MqA3BgZsD9sRwBAoGFQxQN30/v/KbGMTeV20orFBJNjidUuXw/B3c6qyhIAv7uHFVvXpkg9M
hfGFqRViOGjaIipieCCKn/Nc7zZUm53l5i02mmsI/IKTP60EPw/do1reTzTCgX2AJwF2he8epHpZ
QiuTWPiApIIw5hZropMrg5KbrR5Zsn9IpwnXI9ukikprltAaQFW602V/+x3L+98Y75KGS5f0ACqs
IKuMQjpuAOdKglPGJd932Nipz6nuAep8upK+6mI1mNxo26yb3ldM7bZ2s8XvynQtM6Bp4XLYXF8J
X2BNMB4A91/JgauPzKCIWd7V37mFrW1s6wmGdI4OqKZhBJgBWnzHNfRwQHDzPkx5hgdLSGFRJDZM
NYy6qdG2HKO1R4VVQWmsqKLyFOlLPtESNPrhc0i8iPaoVfG8r0Su5LyAxSf7fW9HUVc91O4vcH0z
TxVRepNudHlDborU4QI87R3X0Zqr/PkfHnlYX0ziUTLBcKTSIaUkWonmHRuofLPlyFpHqjhe7RYn
Bl36nyz+FenxQQe928YBkUiYI7ObYoLEvHaDJc+ls5uVQootA+Cnqfl1AmSURMM1WNX3lru8dJhQ
Ib5RUnbmRhOrYkKbNqdhzLZNQf7jK/+HxUxhvuaT2hjKWL3GDf2tt1dA7qLejj+/7FJe0FSKmXvC
Sqf/MR2yvwhDBqBpT1wYu5FfEiD3F8at9mnHkWMP1ph4dsrHvyNI6VCVuynkhaAUHunOTDnjJo4p
amjb+LRZvO1Lt80W2rtEAJ7t4fvMLur21/YIjzJCKPH4MweXbqsj005hW70QpYuMRKsnmWXuhJ0B
l2hFh+7mVIqvgnKRGmIcP3aQRbo+jaHVk6/1Ixx6C/FdB2BlwJgEfmrlZZpUBD59aUOKKZ13fMkO
FMXloRrTmJYZww90b6OLfj0rlAVItyw1ELFUxQhAQkGwq+Ia2KDk7Bk7jGo4/bPXdBA/kgEQ9pHZ
/DMOboc2bXtZhoDZ4+w0BmrCR08XmUb8OWaW8AHRVPgi6HysmEFyO99A8qOqIWZdqIjQpkJW/ZCp
OTDHbzTZzRSOBF5RYxdZz6ruE8qqm9pFfzykBTMJaiE7apVGLJHHw0CRo5z+9XgNM9npyAqQ8exX
R49ERsBfTFararErzMAWHM556St+Awwdic4FUW+GbFzT6VPNB5eBwF7jf9lpwP/kUNwVWwbT70SG
uMfGqDm5oLs9QBM8RVlSvmEJ//DDrUoDnisAiUnsk+hepj1gWq4OSeI/xqXSSPukVd7wCkIms7Q9
23z0M0mm17dYIixsgkF3VTLoydCo3Ht60iDP5t2+uUWPwwp/TRF1Oa+gM3ccNueDa501KTTVV1Cs
oRWb+oS1gpoCLkYAM8+Z1IKmHuPoUpKttfS/Wa0b8O0fG8MXjfcQhI/1EgkMmrvSduxJSMZNwztU
js/N7KmzFx35JH8CDFbPeqx03nSf7ADN+q7jN97KcC1Zgi3vylaSTkXT09W7yumX3rQ1xYZ5FLrS
gCBxRm6KlYvA3UbS9rQTsILQ1dHdGUmdIBiMq6ENYipWWrGkqqf9IH4L2hqw3jNbgZTMcsJXwC6a
wr79w2A95OUuo1ymi6AmKYG3XS7CSH7nQoIOTMfv2zw7ywoAmchFLApByZa19blMAm9W07nxFWF4
eRbpHiiij32cJSoQbtk4n8hB9/2x8+yXOwgxoLWjDOQRvmsDUqZobW4pO8vRu9c+2KALyGIw2N8K
6fsHbhirD3mtHxH412sjB5tHtbBSiZXVPXXMb8otV5/HeOz2iyF82U+BJH4AmUs5HVPlQX8LY/ye
jhNh5KQ+zZlvXzSL4mJ8Xc8CK0HwZB7lNU6Bb00agm3PeW0btQuBJDfioEPIZxV0z6PUWIlwzDF6
sMJGD+UGgl+BGMGtl2QwEKBx8uee+zGivxbFwIGpELlsY82IdwwmzMc5WPs/8vQHyi6ypvKMuSE/
TcZprySorRuGLvLteyfi4wzXEiKgV+zV8Ma1gIQKBSEyQtFXWiQkGCUBqHn4xSoVxFBNUXOdWbDP
o4EJkztoDHBIfTM8LLzlRVDhPT8bBMTqCewLeqBWuQx4or4BWC5jM3kaWcT/DYnHkRu6svdbJ0Zk
QqOpfgE1Ls3C9+UFE2EFhfS8yi88VcFjwDEGPS5OeWEydB08tVUT5iJhbsycp+niodRd3SfYBR0G
gLtmuo/Y1L0WSAWRC4XaAby5fsGYBcOG0s95PdB8YN9Ik+aXWt20RqSNS1/nPK3mZ85K0PrSBDoq
XKcCHzkHz5kJt4OANPHw9GRpOrYDwQJV6oq5iGjx4LSbh0ABIYXP/Apu4uw+fPNOWTuk6JaWrQx0
eMogqjjHvd19jk8MOQLTBoa8yjqEHSub3SOVPx+f8tMEeP9Mtbzb2Z/nFs6I+CrCN8GoGYDLMXHv
CwSydFuyu/cl8WL6mf4yWBig41PKKBfebIAVMltpjYXbhyW+wYeUAXo84tbL2WCMwjQ4xn+D8S5C
JFHw0SyjnnJ1hO+Njw0vwI9clcAyPt5U915K0rbyvQeYSLE7fnftHqlW9eyMPJ33JZKxqDnUBlGs
abbXsZ8EDVtBZXE7wswbBZ10BGybm0TQ6DJeLWMULijN/QxKQQeO1O21s/1DaOKMn73KhPzjyFdo
stxZMJ/2C+DJ2XGDbTOo/T3MRy8qw4N7EFwJIF8LYmEB7v4KGA0myDL4sj1r4L7YhY/Hln5FAw2q
0uVHVRashcNBeu81tNtYKacAn49TpTHbuEPLZZVgr0wdaDB85EP3FTAXvNa5EMO84kPKVsllSGrB
+LGDWpmGlJEoWNdiXcpTafeeSGChseP9heuWYRemJmHEd74tRKtTTSB3dzjgPLGtGm2w2QYhpvqV
+16Pe7tAgDaWwDhU45hmeHYw11CBALCPHxPMSJajeYrGDkovxE5+bjg2dXXv7AilCtAiOSLqTxBI
jxz9w4SR5ZxOrV0Ao7Y65yFtstGmeY+hMoPQOD9UFfjOYZUd0frvzkvpkATDFSjvEKS+DXhpnWsj
y6KoMEm51TTu/bGwi/plYxVgMADqdh2PJB0p8fCsIi04kRom60OTVlpYChiNKoUARfthyV1/E56b
DOXm5ua184jiItbSiNnQlqgKbdQiSZtm3nzZsgQnYSOOCkSMKVqi1cneSrOC7njigx/Too9wZkOv
86WRpWpzEm9V91rKrPiXeChumHjWScN7r61wzkRV2Sz+d3ZdMZFsOClhkNcOt/TC5LX3tIeOuc29
8V6JdNg60TVlCyRbidf5sjK6anm7XgvYqrlbJB7B9s1HM91SsCCjFimTCxDji8sJ8VNNSDKe5LQ+
YmjlaG2TaXRcq1I//rfUWiJi1PJ3XTzPHc7bOay5aEgbf5j/KhthY4vYBL/kLMxSd6+BsHNJMmwA
hjf2fUhDiar6OQjCUoXzGoz2JmSlYt06idmsz/+tnGUwEwmP3ZwqszDXtZUelQDqHCFEOlZnF18E
idCsTanMtCbcLaYPFrQ4whpQ2jCA8L+SabQqpOWBCkM7J450/b5+n8F9f0Dfo3faVBtECz1iY233
Pm7oKu7iOcNhk5W8D2uW2Ty1wBWdZaxYgQcT4b4sui8wJMYKdNg/p0mGzeunzeQxniEn+MBEnNgT
ONEXedh6uS3ASGfYjE69Gi5CJtGQczGLr+SVGVVM4fyVwUfF0ao3S+PaMe15QRRR5ogLhI6SjTOO
nIk24eGgAD1JGadzLRcBK5ycOHTicZToU3UO58G4rMHIBnoeSLENNIckbs3NLd8kL4HeANXZNN/8
MMRHR4Zk0ekr7gB5WuDSctPY5Bk7n3GZswjmMQRlRfHpInwONTv3aM5ySeeTA3eTnFhJqQM7NC5V
tQFSgiXTiAT/8jQ4/xP+xfTFk92UTsFx1tH9xt2aW992edSK5pJX0PrMT150aoKj3R+rSqWEsJtZ
D+rNElni08Sihu/UkQrQBaj/FuKdAxNHZeJUVjGbbOZ+Fju8oMLvooKxjHt9TLV0JS9j5ZPV3CU2
QotRgA6kqk+R/b29qCP6Ugd5/NM/86HKQBqM50ffhpflLEn474oWWpBmqnmacv/PN9oZtigVa+mh
vadSP2WTybqwkFvE/oZDqguu8TzTdpqWkhV8YscfxBrLe7DNySsHv4xvcSPzoYGy3/Wr1SXucg0F
D5YgrMIz9iawAM2E5pYoile/6ohpGgzc8itJvrh2DMKXA4MR2c/50nk4+73hWo84JzpjK9DuX1AN
DUdIpYGPiD60tU+PR6jIwxlSidngKYe539yeuawJW7IIo3uVXDtntfxrYUbA9sWmLOdjeyYJNvz1
I1JT6Wtp9QYQYzVAxmVDmOZyMlPNsCzSQSuNwB91CA1/Ig+m3PpQp/AfqR8yGtRmQZ/KBllc4v4f
5TSIARjyljTpXx1gqeDHJrX0ivhFvnjSIqayOEtp+/J8GEK/KK75DHXQbK9whegXUOj/8wNl39xp
m0zqC+rscLKPiTSlP1uySE7aGa7+N6570kLk5+OwspMsD3n+ZZ9P1P338EGeBL/Q3hcXxOC4PH74
2peJnJUOGuzuIGwWF0UJgeW1X+hpec8Gv0FxwqIVP+u8f37v2ugEFMmjPT2OZvwHN3lgYLCnZVzS
/tQubh8zHo6lNxL62PzVEcGVRmKEq87TJaftBZATulnwNG2UK7zvQv5tfbHKFVUBTdbMmGQh1NaX
VSJ87Lcq7iuR31tkcSxM6SDlBmhczFiG3H2yk65jjdQOBYgUGETo9ws1UMuveWPjHHQ+BHjkgiwE
Rsl2Wj0umpQzodJKnnxUy3THIg1ZsglHSjCZvbqJwFDK0RxnHw0URQufEHPMfs+XsBksQzUemXi6
0UHynAnuPnLoxxISZtBr/nWr6IjLTsFnG5ywXZCFAmMErPiyVwy73DW3fiye0fXJbLY3ZZX0PFZ2
BTW3geMe/vM800luMKyDYjDJB5b5fzEilNUgMnXrbqay0HYX+csqvj0zzCpqqPucwqCbGHWEDTwp
Yc2NchOxJLmg0nBU191y6E9S9oCnWRUIkLbXgFBmmFsGMINEIzJA1hslv3UbbmzO8pEpmp+07wSg
QEcFlYiu5+xUBfy3PJwOb5FSzLNZ5RVsPNNqE9QZNsYYoYcLDetL4LiqiLFtufeyVZ5uRSuUFuCP
WLZorlaFbzPZTQwzoUohj0VnUsIGhA3/sgWoRPRw+WiQMkeWoGgnVPvJaPT9EgwLac9FDS+Plsi1
wzZCKW4xLMbd8zn1KSUssWz4v83EKzEodS1DiOdO7MHc/a8ivu8vL8rUpu/UH5cK1YN5fZdETAEs
SQ+v2MLBXg9hCra3W8SzJvp714KUR1q0zebGZXGSnyeSThAmgQul3YmdSAZEsh30boNvThCHFUtE
AhnjW1X6tkEQdbJvO97MMZNVqiDwOGkFFtFYH7RM/hWmOHC1V8vJ3xpeWDDaL/kzBaMI1WuMYgEe
yE/BXIgwWAMFoDlpMObpJFVTnTGkYFpqWqhrrKA+cyn5r5Vi0/raWiAl0d7BcLlY762Q2Ew29kOs
HoYwkQl9TwyhKcI8SirkByyxDgZzP1qtgzoplVJDcKffFR9ZPqY9us5rWxzDmUHkusQdImuTFq5Z
v7nLrjm1ugWBfx9QlMNoYU4yoSn4+1qj3EU52IYnVaw9sAAaKF10Tf+xCNfJ0Pfotr7ZxyyWFMit
aJ0L1nSmJ4hCcyXwl6J9CmyZbf27nRh6O/743NO6KEPVqXsJcOPAoZPRmC1swtAQsjqV1mvNheS7
o/XqnPnl3gIuBMJ3lEWRZgCR6pNpw3VD06fFDfK3c5/7Mb/rNhcc16ZqYlBZIdUAaU75WUQlqipH
AzRXB6Ji3FhedLgYTguYR5Ik8yQPxLAsTHwOK2JfEvKM5CryDkQknh/vXCysjaV5pT2ebq7aqIpB
1MUw+qWDfct96UxDTzoydE4g1MTpOu72uIy4s5m21yVQqZ8hm2TSFnjRRqiZmgFd9UpuPq+EyBzc
iyOPZ1SzQjnHF1MSr6a2hwIUgNhm7dQZplj9tG1AztMpB0C+zGkIy66k1BYJGwEXxqTmFMT9n99K
1+2gEe0NbIEzva56xv5n/PkOX2qcRaeEmGso0IFQa0gidFbR25Y5cNd44E686bsXwTdg2gL0LPDO
FK8ISxBBSrak81OSFqlu0J9OhZfvbzS6LC7j8yNwxgg+HMgcy7cLi5NJNbO8GGst+teWgLSPw9wc
rGgVm8fiI0xFK8w71yTbcndLhI4W+33r2OrrITRHdhLKsgFUgDPFDWwWzVh8PwCp7N0H9odx2cdE
mIKWaMNpGIDC0yyRfMSWxIQQMdzpLnNZEYaSsO6FX2sEonNW4o5rQLjTzOsO2xBSG/GXKSk7OTB4
3sbvRBAtgPzavyk33dEF71H9/5HffiOSFVKkwQIgBprEvu9fdahK7EEDJu+L0Tn9tQ9R+gkXf+6J
nQJkwUnD0tXvx9ZhZZKf/9EXwBOIHbZSerhKk1/d57/ZJBXTSo3uwzuPA6PPBAL5NvQzieZTHo8l
ArBMejbdggW8KclfsCicUBfeeZouK0WO5w4x5gN6VdSOXhVcZ8yHCb6DqRWn6nnnySyYmwCcyPDU
DAQB52or2qLcS37Gagw99DBC3ex1mnK8k80tUXZ7S/0gaiB+s1FaBS+QOOjeSBn+yl4ve8jga2fy
7g3jxyn1zMGD6EmaIk9u4Uqfy1JOcpslnsqw7ADwwv8+pHCeh/QI6YOA2mpa6JRuET27djxl49rJ
cuo3lqod4LikWgxs/eWW+au8KF26pwjkfKyIxJ4Q3lQHvYdDQ7RggIaMHA53t3PBe3UX1pcJs6Ss
1GnOIB2rxsCMO43tmJQtDnOIiKfikpkf0NhaG8ujwTqOPZ9GRkj4bQcgjqt1UevVmQRpZlgPF1fT
JoEaxJc/vJedMxFCf+eV6sWnR2yMEkK+ztABj1bP2ODb645gth4+vuIcRrXf5B94WpeG9yhpQOY4
7JgTyGx+z/oXclrmocVH1XRNCfU4G8B4A4whLGZy4S81Ex+EhDonmHBQRwISLFaa9p63oEchtt5u
Hs3scSxOG3eF3Q0VWzXW9u2lZhJFtEcG6KlTX9C+F/Nheg4msxxrjsFkxKt9mJbbXCPO5WCEOyCl
HB263RAftGilZb97OBWPuieYzNznW2w6pYiCqGiWUQPmGQKfE+rUfz7PX2OSqzZztjWoQocWo1ta
ieIf9nR/8MTg8xu70MUAY9fEp/bf7MF7o7iibEzPTXhQndJdiP2lubVIam+7tX55gt0RzJP5eS7g
0xtgGPDD/uXajz+LTskpUPqd70Q8IMlgi4cwYQpIjLNnW7ykmAFjUesHFiPFvlIgIetwuIEQGr/2
w2zbvvCXatWbk/fFPuTGcZGSYJo0xsB3PGZ7138jKkNKDSRRe7AJh2oZ6S/5eNOrIoub/PC+Y5lo
b+hfENSCBRTUgxtM1f6PtVX0fphbX9ew8C3v6OmosmgyrC3kJsZ0SZEvueJa4rfRA/Cas23BsozX
yPV1coX9TxQVW6iC1B8F8Sy6AhaOQbQWFmY+WqXPsJ0m77QXZnH7++0Hke9uE5RbfF7sd+oZlmhj
2ZZAF+Q2xqSaC+fhKukj8L5xRwQbjyzuRvcqeaOPsckT+CJRTIAFslwwx47pf6Kzu3s7G1JQvRC4
5JkoVyoaYICV0usI0ssV4i06zX9MLWFNjkbnrmV5/AFgwotiniuIsjbqnvKHVG//BVKKSPaaV83O
HiD5SE57tvFad/upbasdW+4jIm4HXajpbA/CbeYKHMxBzl5ZxEmuPX5+BkcsYGoQPpqZvOkXUR+s
HCQEmtxbBNeGjDspxy4m6WMZEj0dC+euf13iK2Fe7v0rMPa3hY3UBJ7zZdjyMuPjo0WAFlWCFcOp
Qg4Hn/w3Hjgsk9bpbazSPKMERpK3crR5QGQ9hZVy1KcwsL9RgAh+LSkUNpTVvTYN5fYh1cDRH6lj
e/RqExIpvZZ3wiiX+mI/eTQMJVEWDJJzDfSi0cF1qLztx/nivqin5xQaF4srTBq4nlr5TOdE2ZBG
FQTJFAAA6YiY2yhS5WwTlSiLoIYBLEQibixrYcUMMs9xbfJ0yVGjJY+pUAt8r0yDvO39TJiji88A
5mdfw9NGcYPznYI2KAawZXBF+AYPMiD1k+QMmEXWl73QBzy4IpdcAdK0hcwkxh5cSe4PNB68sh4j
tIh97xRapGwB43/o6j+79jD3b+J0cP7q4HRpNW1QKSuJMCjqWFrMXrGQpPTIC2HGr6CXOH/Wrq06
70ygHZK0eVLagONZKjqd8RHBta/RyIJOTPNGv6YFizoloiZceFPrceHlLNaKyqg//1r2kKtiqF8i
2VZZHHv9fOnOIFkczhGu1IVc6R9gEessqADK1jDopXvQvpxTzVWtgDUCQSuah0enSDuUfGH+ORg/
V1XLP9psgI+i19Eyq7Q38MwydpQZu9KBnSXO2Ae6SXyYUq9t5nllZwjaxLF2HLeoMA+F1l6IwfkL
o+2Rz0HgIgwCxlhLKyw/BW6ARIrTmGRrmHE/T9M7o+PB8CzNVnvPAGXn2ZVjjKszdJnwMt/rtD3b
YmvniqxIo0jfqTbkEeonXBWJX4DXsNkfXNYJhLwuXIcZ/wdNpJw1PxnRtD6OYSz61lfSniNGAxbp
Dy6hP+geLYuTl60yoPLAX4MayHpA1vWD8V1tlZyvLeUIpxiLkAuO2k8Nin/nTMunkiXcf7E5nhFw
w2ufldEhT+YdKQKbmptjZnxdPuKQeINOAkMYGqIAedmr5AvY+8DrumrlPjejcQY8aXKn69fBl8NO
usisKxSdKYosJLld/DBWNLxE9V5JScYzIfd1ziarlmTjPfprZX3vcvId8P7x2ZRvy7NzM5ZgvjhU
PbItWajz1Bclr9B8WciazGnGRjHlQv2MpC+l9F4Sn/Te1GrN7G3CXuJic4hoWSp8IuqobE2cR5eu
HVQ2svE8fB7kWgqZkooqUteK0ucKoFqhoW4iJYxKXuLIpAAFv67fa4JgmoRUIDamA0YhZcI+OP1K
idwzEW9LS1SkpzDZaLQT7MqOOh7T8Xq0eqq0+bMEmlTXOhARncl/BCipcC8sbPjV6y2BckURkmO3
NPVqcyN6dX5+SW+gWEdz7B0zVfVg/vDkC4I1m5/M5Roi6OPS0xb9gsbAT2JesZHfHGYuCs9f6/y6
LvlREaTt0ft2UTAW9PZEtIw7aFLyDt09sbI0PfRncdK4thbDffSDKrgSXAVujwB4gVvqVtZghYBG
+ZulxZWSHiKsnSFX/uWW0TFd7G3NxDHTGg1j4Pu3nHLZg7XWfOeiGAmem0WCHmnZx7D+RBPs+elr
sm8n6lHHzOgR78n3yGax51OQbqGZmtDom1aEYu3jBcQAV1wkgGyaW0ngEXWvmOyb9G2wvFuRAS9D
aLzuRk0fSuZabR/XBsIvCR+4QGuyGMb4b97qtBxkZgkECH23jkgU3N5zAlBQaP2s2nmld0s/BNPz
gBuDNfmrbDBCteNNMzKeEelez9RVZlenolB85Q4v4wouI3XLnGbs/K/ASgxM+IPxfbYbQjp3dI7X
wMnIJfpWJxNNowT+hjzfz8SVha1+5CFY5Gw3/9H5I5oIcINBgVwF+OZaTGvm/cgn22agoS9LgXvm
280MA/e86YwLiU1z5lAgFU+xYMBf+9x2D0jNsfawnqMKxMxfzTMpT3DbsvTn7vnTGsQZ0oM5eTq9
nr6IrR219YAfLzy1GBkk9BoKOpsWSj+SdCNxX2g9M++re4jjS8ttIZP5dXHQX0ZpQdKHDYvxBMpi
/D9i49/hO9g0oBXJjX6Pqx4JQo9evJQlGNl5yUr/zCsoYXTFVSr8O5X/xCZv1Ote6b1MC1Jutawe
aY953qQf8aZ8cTL3SXNsrde4mFK5te2yjeb/fyv37hv0FL+75NLh36CjrNcQU4DngABgfoggGXnQ
qcay6WvSxt3Qz1N3swJfTnHkwroknD7RwNgSzykcOMcBVB9Ngvh9l07TDJPPJO1FR7APeRGl85mt
5fsnYrX1spReboSN5FVTyD0hX6XjcYkhdKdcyRCivZoApbprdh+ND0tMAckEtR6mnZ1iOehefdcS
GoRS1bWnNcz1ECYJgGJ3WPXwaD4eo5HHPjkGIBxRjf8zCYbDfQnODKeIYeufmwRzT6ObI14LvDDR
xFmz+cnP3fbdRKN413K4pHzjfLT6P7mEozrQIqP9RbmsRpmxRuJ6alqy1jUH+3JOmAionksTHXQ8
8lN+auLtno1A4+NqGiZF2JDLxL54XBlwUtUb5G9+UDoLhKOX34maTt+I9gojzofs+ZFtSKJUkpwO
bEhTtoEm1CD6PrTLCN+JhNh7opLToLU/piiIEwccEdNTqDyJvD+1ZlGBRwRmUsAaFK8udaB+mpMH
w1T66pZdYvRp5iWuU3O0Mn0sVsSzg+ac374DpaLLVFi/aHbBcmQI225VL9zNS3oBSSQbOX3bmlr6
guuAIfjyNsvVcn+UeoUV+FnSmQbCh2VOph/PH2iw8SsMr9tH+iD3sXRy31IHcOSBnzPCuXkghJ3/
/+ZuLJifWtNudD1gv2HBY2svtZXoGvlLw5jKFgbKCORmbe/ENRIzwd/RyXfRqK/+HpRzcIzPjirR
C9ewyS5FuG4KJxLOS55wrxefXlowKW3WPKww3jXnjRkbrVny1OMqsb2VUfE9Xb4oEYVw0Bs8HQHr
IzCkV0APnJojpOFpTqmHDsEhlWrdyN9XpBY6SBDCzOI4xUD/Jx0uzaDbMRQQj/vQB6iIlAtffplJ
cHpnY074CtSlW9Z7kzPgEIHzh3EZazDwpqSU5xNPbB+THGQ2eqh4soergQuAmRVsb1ey4AgPOj8U
X1AW11x1PhObXrvgq31OD6iEFuVyo95EJGd2M/ZlYCuvFYSem32mnYmXozpedAkFuTjw1g5zdHrw
WW7A9X+s9NssCuFutXSrbu/JTHFD9WD9FXmHLCCkt91OogantHA41I7MH+CXNXjv6t0E1gVjuAtL
yk1rLIxxQhiC4vT8AjuocHjgf8uxC603eVf7TP9U06r770MoHYtmfAlulY/tvF5FNpzKDEsncudn
CKRfRybBDCvkV1O4GbeKUEqvpIgEqcoPlcvoyjb4pKRG81hJpFx4ZwdaW++qZOkJHboJWA3EySR2
zuGjkqCRQoy+YEC5mXAMUVgI8JQEg5h7hlg4zUSVnKtFuJJuSuuTm7xuJOUwj0pCo/7SmWG8pR9j
DIOUwNdu4l5poLPoZn9AWDECY8K5R+2hCwOlbrM9UNrNoUPrfk2SpnHSVAYEEiMe1P1/f+bLT33Z
yI6Rb/MMmehZrlmbhEkrk4p+vw1521Znv/jbxC70YIRoWdaO6PmlVKDu4gnV0SK29sjyF1ghVhQy
YH74O+nyDkj0VAn9JGW0dxafz6MC8gJp6CPMPrB1EQskyTmtFFlchvZGidoTaOYZsEKR9FK5H4kz
EXkeEYWHfpFcn7nbzztKSmA2kPqvOppfuODP58fN6OJQIHWmfS4Q4pmrpVHnW0pqXwfoVzj/XtHZ
oSThoMG9NGKzKTem4gtQ9DqYQJCMj74pIgI+pIxcwihs2wDd7paPJ09c0OADWZxnzOzR6YidxsoU
J6FpmKQ22+CkC+f4d5zh37iDzZ83ElZzKycYRkLJw1Bpc7dqw9lzdfdE04kT+Xke5qNPUrhx41is
hisVa8VfhV7xYo9Dzfkdwi+tBpmwQhKtq3AXJsivq0/zz59VLQN9UyULPUU2rS4hoN0KDN/oxmgR
LRJxLpDZAjd7gZUKjZKCsI9LEm+bFLkbOTtf9lPu6/i+Lk0XypJDH2CwYLNT9Lzs0/DS9aOSz3zC
VUs/K9752gKfu8+6cDgbz6Q/3K1tCBNOBO19p5s4CUqYJRaf+low8VIAjQub0UG9wMyZF+8Ym4sE
x6lailHAxZyOQYpCEjLYOukbwIPTqDc8rgHYruUh6AMrUKc6iEPAsk91ImNeT2GRl6WuYqzu3Xbx
ojDeMHuu1jZnmTAkCSl6pkd5xoFNnrqzjm+jqUmcGMKkRNkvm3iCHvSyRa/0a/maVqiTTdTlTAsi
nyD7czTMkCntOfx81sSuKB94+GkuTe7xBdAtVGWM2+/8rfs5xkDIxrVSFA98Sl2Yfdb2ImwGae2x
HjXmnpssSKIT35drAdTIC6vWf3tMCh5bdEvahmBKTpf9CpTBf2WAhf5TGsxH7ZOzaFJDkPIeLhqD
zjozgrM3eX+0ty3H/d4+ZPHDhAkF9XnpaTdVoBr7w3qGKCesySuDD3w0n+LwQvy+zqMjg6sDQoP5
BGiT+bT6HgKxg7yMiaioK9DGMeF9qKNmICPNCgnDkH1muOHzMVhXkQENy3BpfGARCoeltIDptFBa
4Ec0YcQD8P1fx/TkpKZKnFuvftlBtJW1SsK27s2XVxoe0t6jgqFF1dWiPrkd00i4YfabK6CyK041
Z3iT07dIT/Y7vsbTHVh2+zNZdrvd8Fkf+rWyLLIlYYYjMZjqH2TEEaYKg3dJXm3ev3s14Q6zBh38
PBilv98jiOYf1HMVuZcSqmJ8REN4rWcu1bYbigR/KpS0in14zfbo+Y4oD6imndV4L+jQAo9Sfj85
q/DrxIzvBJzG8TIVwDPJe7R/xtoDAvj6veNhV85IReif1dtxqaK3HNkmIj62jga4ERZXKM0sVNTn
xDabJnLLlsu8wMusXUyuFujyKUOZTIIbMKtZaa5eRj9RIWaa22ZxamCbmdpZAP0nN6j21VWeTk/P
857/m+Lb7e6A5gLxh7xPbGAoNGSOpiqOzgngyhU5Caiw8PUV4TmgTAe/YDVI5Awzf75JkJBNf6kx
K43xedzUe0jvqFP3C0v2zbHEzAB4p4l9tfW9PIBgRFc3K0bl9m3GBQpn5bJYsfXMDfpxQc2q/mo7
3YUuPxkrXWfUPSJ/1IFMzZ5N22Gxz+ihRdlJIJcwpU57TQAZ2gSoQ0P2nsXT7bYqn54RAzKm74Pf
H8ksyXhbPESTGx8MWWiu0tfgAvwUr51B+GLS/9ggcO0R7vApn4ZbxK/uJLG7q1eusZiXRHguEq6n
kRkhFrGK8QgoOiIc5CmwFYpkbh+32ZjgFilE9cC7abnS+BMOe5EhwN7235JXGtzFK/eO83/IbakP
CDNcQTECZTlhRVkKC0WBvKGUrwV6Qw/ANECBjEQJKIs51kMGTaBV9dm29S3OauOk1lJCqYXWvVmK
+VYCT/CkjzkxyQcK3h8oOFWLXmc5FxupJ2V2k5v8YOgUN+LDs/D/4d1No4NFwTfPPh2kJ5znEfnW
5p70iFHImYaUZBZRB5i1j41lXdTAeTiUa7jcd9Qs4lHJ0STS03oIOPLxlKCwAc4rSgSIn0Z1FhbE
c8mXmQstrA5mTwGqhGshtigXvrjVAWbllPrBJVvpnh6LTpw+IBIldwpWLBJ4E5MVIbegrcgoWvBZ
ggd2F8ZnsRtG7nxpkn4WW/KGhot+y/hfTcf+Qhm36yLNc7ILfrVcSwkOZDVAyMiUZ2gwKLD0zDCm
385SRB6vQVkJWoTE7TaQGLCEmQeagyNB3d2pLDeQYYR4q1tsNqGFzfSgpRLyClWOblYy6O2ypSZp
+x/TiHeBfOK2N9PTx3L6vnnS+mYwO7gTsprhWtSsK6A1aBpHtWBnxEdvc0AgMmmH9Yhs6cE5o6gg
wCeE+WnI047I216PMblMYUREP4mnlh97LoSUQSTnpKT61bMpP4GkN0vJXYA5rk57m69xUKvnpr9Y
YsjfGPWXI+gOzNaVnQPf24a0oRRRz4czsd1RWHeWAY5IluJwx2M8zJyABr5cda+tdFLT90psMLhH
ik60OPrH5Xt8trPWvo5mvH5fvzdMiDvAiZ7tLhcwM8D9mAdtPYGqx8tL6J8kQSr48QXR7aDJdHRg
Qfxbeza/hdZlYqjrbJZj5lLkmSmrUSx8kloNeC6L3PiM4+0AAJ7ghSSiinvMHxv2YMxh4ZnEzXFR
fn3iordneSiSNKR4YvTts42kvKk91nz6yy9q8IQpBYSui744Rm4h0AWl/SnkOTW/cJ17Y1opeDkg
wqHd6tvvh2z9SVstENG4Y0UwDR1VAA2rONWoU+STa+AfmMRfxIIOdA0heCcc9DAcrqZRaW1y6Sgy
ljq2Ii2B1geehhh9CsPIrlNvhdSd0J8tfNJSbxhjAH3fyHK6fkDpcd8qzG37zgTcNN5hWKXcL0rv
wS8hMwcZtIwiqMki++AKCvXqZeMZrHhCs4rGkbeOswqyePkT+G8dpWRxmoxooD4LfRn9hz1MPZ7+
VPYbg+U7Tfxx/q81P4T+M9tsHgbcpkN3A5dQMYCCPyQAIXmZRCzNoKUWyo25IcLmYjov03tg9T1o
2kttNDP3zJw5J3PQUwaELu+EVjleDVNVxMkYwDryfgb/F1rdQfCIlzwh8eAHPlsPi/DX618WE2aN
P0/Mg4i3XGbGFGwc1PoxcK1hY6mj++9c5fmZLYv+3Cls3P7w6zREUi+zQHPPUyH3fGvpyhBOrIdu
kbFrSjxUow7moiNbHbEOfWARzaTCdy6VACv639BEnqH7eo8dhE2Nr+z3i4z1EBfmYN7FJcUJ0S+Q
MWYSTztebSnCSryu6QdXfCM6zp14ml8WoRvUIfthryJmXvE8JSwZfxs10jp0swmnib/FFE5X4KBM
Kbj0xFg23oHfUkP1UpiXGDWCcwBwbDYklOuMMOBgSJUanRvVukEdTOq65dtFBsv2kvgmVLHngJRR
PZT84geLyKDyCkd/eM2Ik7tduOO/fLOxdyImHbdf+b332P9SrAqU6XXgEsPiSFX7SH0vnlsHFDZX
rMcBx5V1eL7sdUtD/4s9labNWuLqX6FKpG1pbTIwtGVQ7ExEwYoCb0w5cfASo4ENlRF26rAALFmQ
0esaB840i6RMjYugdPTVuT0l/ELRm8m1m9cusrRJMOw/wK9pkhvHJ8gvWzyrvl0MSNAMIZicGxX7
1pnkn/bphpi9MagthUA2/5splLy2TKWN/BjJlJ3JZ5B0OGpeEx/uxlTgetm37uc9KWwYGjtHqkAO
Ezi2gfzqhHB/iiccyrE7vW+zscStToBH2czfZhPcPxMISe6l3LeHrze+F1+szNosttxJWi9QX5IV
H23WaxYivGl4BGtO+zrzgqX4F6Cjgy5GIDVb9N6MfTZXdAzGP/PhbJphTv3KLU2SICUEhJ5yseKh
yBSziik2aVgg99eAa72PN8WpctwqUJwWsn4SgzbWnYZtqCu77x3Fj33yhcyDBOVXHFs0O4iXbXsr
Da+8qcuYKl/gMARY8QENvSS1NtR/DA9wCBYj6RgkVlgomtlIkBIv8G5f6OaFlgyuYuZyHObWxJvQ
LmRAocCFGWvvJ7g0hkTi5GjybaEGavs8rPfn0ItWA59nqriEgXMbW0rwOrjpOcXnUDGSi3XiT/TP
j41CuBxHzEub7ebBfByd2SJY+3OomNGJzRrYKg6tbN83qPixeENi0lSzIZXV2earuYc3UNp1dKvx
GbOXK9vy7BjjHvaXdEM8nkkXEhVOXcrOahluj0Y/7/DdJsXOSOYo3wwp+tQSyLgo0/4AL1OLMN4E
eq4cZyBGq8JXOVGGZ6Y0Swin3YD6C5T1ECnILKBhzl1g5grg169aZIdbC72gO572VO3iLNey9VY5
5f6QuGEeSSrttJFIvW9orpBPy5Vk5IinhI1VlvK/y8hCyIHRSMZqaAVO4o5rfd7N9lUrbjwCnhTl
HYNwa8hgiAg2McMFGihXt7EiihltWSUoTt7Vzv2ZDUoBjjCZ/UavBlV8+JTc/7CJsmmp5xstebnu
EQ+3dTvuTs/frAvZ98+s7d1fkJ83NVtNVJLGdAtdJJV/jFjaQcJCATspWK5tVxRhZkcPbVZvz5CC
f+Q7iW60riPonC0GYNP75B9xgkE4BU8hFa9pyBWdOSBDdYCVZ2vzDIRmAU/cDs/3TacUnpQUDNbB
Tuh+SWB6e8M8umAmmXNNaw8MPRO1s2dhdncKQIP4rvnq66OPa1eFsqPzZcL4Hq6ovIwQD5LhkMRG
qgn7rBhR7Iyp0yMJ0JakBgbpD1KyXNqZI5xOIjVv/5O4b1YmmRUbdkUBtMg8U5PF/k15NXQdGuWh
iwwMWHniyyX5y5Ld/HI7TCVpiRLpWC9os75YjKxGJPRyDPasbgRHIpccGlSUfIFbeL7bOjEVCM2m
cOGdA0HU1ChiuxwGpDS0QS1fQyEFKf1M/vvkB/yzt6Y0CUJBbCqdLKvt/MWwyzzUyvd/71fj/0jZ
m8LCiRN+JB0PbPFPHWyUtjYL67WwAdCEsVxcjJA8/phUZePdneIPc6pfc5NyKrpuCW0SdPYtjqJB
SWeXBZXPuKecvYxxM6ix/x7Kb552S3ys6CifzRpOsTy/JOwVX4feU0jHemsCWaP4osc5Z8U4XhOM
WBkzwWXsjt9NZdbuH8Ir6oG78QCTWBqjVjMm4niSLR8TlsGCgBu+I63RQ0SRxR0ntOgrEgUJ0LS1
VakiFn3JPmy0JqUjKVa/JDD7zHTWms5iyCL93u04Wsd3aeG5uE8SvgKGr+68n8pDPBP2tQO/KSzV
WitisGGoheiYxKKdvMQ+VGlurps63t5o1c8rEQ981YKqAmZdrb3/y31ANXMD1uFBCmYpcET9irhx
EbRrwtx5NynPAMF0cS6aDwi4ROYxzNOvc86H7lQYDj1TktATbG4kWOFDxxwt/I0hNS9PtYMEJBzs
SitkViND0Wtmy5huokF57rfEa+3lmw738aRu8NvoGtKJPV7ALTIAfRcszr3Ov1JZBbbeX7cGq6oV
h2AjuczOPzjm34CF5I/XcheSOkLPIx/oHV1GhU6OC+KqLzKW+yjsjCXOpV+bM8XWh9D09S7xsmm7
9a/P/6DvnQYG1Hpo5kFKoYzWzo+KNnMzbNRWl7ssFVJ+Z2M/VsVY3tE6VndQa+d2Kdsqp8Slk3vT
R1lAr0daWdW+eknO5LX7Tq8sgl8cex4a1N3RrJL6LQ1vW9/6FOnYRWFR6IaLWyzAJ9NA133/0Hb8
Xrkn4bxNX8K1kD9sAzjiKw88+I/7evsmN/jmNUEHP7pNKHiORHQjQpcytGQqi47f7r6xLxVHj4Hj
jk+zHdIzVAkaSG1xQ6vOe0sz8iiwl13QDupXJ04JJfFPXy0+Ya/Y2xYGcY7dyyY7AqDtSPtY6mX8
agkc2pcfyyjf/1NHsS4oWaoYVc+fKwYo77KK7duDHo8Dra+oscWcnKjdru3dKq4N5MkhcBBsxjJw
y89rqZk4lriNi149k7D8p4vkRdo45eyE4gXok/nR3JJs0HPUoLa+g6L0yqrtL1UVNlO+tokWDpNH
6zblNMSCey6lFBIwmWo+fAqi9xRGLMM6DoNf4Yqa660Gf5YH2yEWZXlCjpT1ZUItzGOXVl/gaqHy
05ZGrfeuPVz+R9hXHJUctdDmgJpItBWOfwRzBUa1/CFNvvZyZAblnhLGEpZI741SUVy1e/RF+m8E
1bNzNplCQHYqwyVP6h4O7JpU5Nbk6xXtLQSZ4gQA0iHeZVyzArMzE1wxuIm869Y2bCadunIQIUx+
oN/8nRZ8YuQu4mLjSx8OeDJf+699LyA22LezUoRogd9q5KGpH/2rKsRJhQaakh0jZ2c1ddnLrt8B
94hHYLr8E8Lkbe22c0+6MDfyrefvZDs3ws7O53CVYEGFA577KNQhyZPtEGAdpPcWolFaY1WJYgNU
GBFkcCbKJZxdGpv1HLEjxC8g1PPsx0Pxw/GnbwBrbccKHEHLRjpPWyCQ5xuWN7nHdY4KfZFeZdlg
ioJr3o1PoXqzSqcSeHyFUiUbadAyG4BbsdU4ZdUL+cSiKEuxhMojq6VtyvGGT6zCH0DXbk736Xlc
elw4xrJoSGXWICqZx4AV7wlBNH6OuNXxr08ZbCZpalLaq9Re3D8WYJyYN7l3wxGgX1ATqgwryrCX
eo7TegoHCJ3zuzuZbSRqwzOaRQkjyTQbongHuJUdYvH/wpCb/AYSwJmsQmZ7stN2iIgHdnwmaDtD
8y2JBRukIOPOcKMDO4jKJT0/ZEPRoQiISqVzGb517gH5mMrW6mRoGEPinLtt7drFPI2aj9IrCVUC
iz5Ewe3yXVjZreZMvCJ1w4jQ1durt5X4Tu5t4OoLGUKd08wGXEB1PPSWG1KGw5Fbnsg9FJKwuXmn
TaeqCA8b1wOvHztjmuR/tCnqVO83WxxPlAqy24dlXlZvtkzRPtMLcYlnK4gd2lPrEBAk8BVMOg4J
MlHyhg/OWo+SbQblPa51qgaONGbAZEm+r6Mac07FmeKxDCsogv+SUwqdGdaIR9fKxm1J7MDPZTpl
WNYlg3ONmpypuUEyG4fWFYZxwQydGxCVya/rA/0F5RN1AnFnYyI+AykEABLMhEmEC173RkMyEAxI
XsCjac42QRuaxIuWYbIdFiqVxSXQ6MlQ6F4xasqvmQSqK74os73woWV1E2/HUAk9OpFTPozOkduA
l+kwmWaDFrIjMfeXNv1seNVzEyP5lf5/tmQB+w0ut5PSW5BbPbaroV8TxLMGUXRLNt1ToOqzdAAE
kOxExp9KfzVoK76ShfmCtappUitl0Xv8HgPrHQctEIWlKIw9D6q4UCgClzkUENI8eGWrRnTFc2LP
c4kIeaqDDDCqSmIpKXDiR4o3smX69eFJyW0Uffq/Uj3cIY1TdcFUUE1Fa9rclDlW94pnnYXVjdW0
NR+eBbFJt6OHapNOIFlluZePfAc5wd7z/WmMEcxnH+qr2KYk5pE/l9rmpy0RGE/4zJGxPDCGJ+qh
mfPgH89mmApxCR0VANcikRrianiFWYl0ixoZXNc2vsRWpsOdmIWraKOGdoQJXT1m+Pb8YSrMt41L
QHi4HF3lZUmIkeyRIlSK9Cx36q+Z7p2QVd1Tqzmg2y5gBYr5FdA8DfVnfx4H+yTrfyG2H63i0NJ3
eA5COHE/xM5WSznGaUMGkUMfEHoRRJje4PQSk5UqzpvDKG05EhRozprYI/9Nt4OmVktmXIstYGUa
W/f5nBq/yVpB4vOUgyYU2gVdt3bPrzaJut1uk8ZrufYDXuWpGP6nflxosYD0VB6QESnRLK4NE3kI
96skeg8a5v676taZcCuH6c0XNy0o0DQrrHtVI1oiD1STWAcd3R/r4+y3GT5428YQHGE1CCqQCbm2
6aulhIm/VzN7VWFpeh8oVrkY6jwhPW4q9NpiG1SloQl/LbqxPFD+hcgCXiVcAi+2bPk+lbvoJigu
D33tQKZJ2bfqKaWzqct3pejDAGpcR9125uumeN5aJq2fdDVmM1KDFLni5+WXK73grb1BbAeuRFBt
eUo4XQgwvz2tWRi8Jf83DCJeTi/+/kT/7rYlTWHVqaZFgRtONsvxP8/jxIPF7bRobfjJfBCFYwnZ
xUC970OW6zsffEI3tYJw4z8cTFtYa+xfnlOXBjsDH7MDvb1BRX8w8b3gPgDDZQ8FgYuQKru2TLBZ
SwzAOA8CeoUWpNpfz0Q558FE9xDtWq+27kWfIVhm4fKimqja2P2K6C+K4KGlr9Ve5z2aEUgqjU+1
dNieONmZcVmuLJzFfnIlzBzOwFVIknYkRR2RfNT6q0CYLcaHWh44s8u6gval3rCITjZ3ei7+Lq0f
UO7ERmd1BVma60bkGWGX2B0Q2QOrGx9lNSYR9wz2e72t9sD2B4FWZauTN3HUIqumJsmReE0RzwgR
hAXkjxt1O7mH6QXFroxmdKTjFHPJ4BM4ECTG3ZhB1oy6B3hTse6bDSkFo+iD2fbgK3yKyPR/dOht
RmE8poJ4bNE2W0WUW5dcc++exJ8M8GI59DaanpP41n+yPHP72BJBf341u8V74K2m2IQd2oanToin
/ewt2Pw92z199v9w/IJjO72pbT+ITLmu57CeVKzPLz8sP36mmjvf0e4MroRQnDKiQkr80rkum6Ln
skSC1NCWvPprik1b59m5SJM0nywThiW46v1OotJaDxLyj1VbcvlifwmGHbBZUPUnL+x5Jlk9Amkl
eYc9GjjLXGOlP/SPfFCIkdwocmVkptk9ghmJnke9TdTwNcf8UhbY0YbCY3tDsOQuqjDikT9yh/jA
9u039CCldvZl3BHvD5V/Ix1CIobzcoUdY49ctKZ0BIgKsvs51kbDuYTZq2BSor/iEoi5t4jwvttg
DobqT9pViE8pZMGYqGZ8dqFDNTztWzeMmxyXwudPTBpzw5dbWAxYEmNxlQU5oWS6FbSH4PVznDix
fYgIZDHTIxCRh/PQQQdBy4y6o5hEid8Ynx94OTuniIqKRcbSGXqAR7h7KOLkTIUC8Ll+1Q5/Tkrb
9l7SegnuOjEgh/vF2gUFeedcAE04a5n3HaBCvrf9lfyuM6q3/Z2fL+hP5E+PblSroGq3lRHUgr82
CxHsRYqpYSkPuVWPr8izJr4piDc9pZADDvxKkG4rOltsV9mN9Bd/BWyxJ5YfTWyp3Zz8opJda3Rh
Chsr8VcI2a2K7GZGA4B0a+hFWfTY8Tq7J7IGMzZHNZ19yjf9jGF02CFqYca+SjZkt6DdXX5P5UaK
m/iaqS6jCWlnrzERsqrG7mL0hPUnE6GR/WJR8SRdW2ZbcAVGK6cHcYXu8UsdxDNztAVF51noyZoj
vAmqcn6uM3FpIIBTWG7o+uwAaIY+ri7CxNojd2Uy9ZFW57sKlPOGoJ5zQQ4KuQW4zLGeN0wFn2nT
TsWgZYHBENxM/mSlCeGRKSlzeltX85UiDVwL/X4w6K5G5la8ecsZvHRf0pSF73/zkSQ60fbI3+wG
nmErK0AgmkQqzzolpB+4cT4boR+QhhDb77KBn7pXYiRoZTPC8L16PCYFkvRSN4bsTi9Md78OyWeL
/7l/JaVMBv6dtWj2GC5WJ33kDXrPBKn9p8DRZz7/0IO/4yDegkyTGnkdUtl9gK/2N9iOJwlZdAu0
UylTKAKQ2WvMBWwmGDGnFKYfoFMp6WwP8JrFIObzW50m0DnSC0HEiHAhIFXtO3rZso/EPVNKDCt8
3qKRA74eujrl4npeO+ZJ7ppWWlxJThunzXzRDFKytHwK6ON68Wygswtl4zrxcHl3cKwGcNabtd6c
eT2ZNo3Q/Bl1+q+rePbaN4hqY8ePshk4QppOFV0GbOmYL8OeoOLLDjneNmnmtnU9grRhnvEN09PB
Q3kUOQCi3cYfMyEt6ZfWRqy4ECgceffrfCASgx1hucPmFTuEjrkFg2OfQhRpMjFBD9xSOG0k736H
+/t0APp9EQkgS6BClCDyJHVCe5wqy10IyLajrlbS1mG1jtV6gQXfPuqiDMgn0ssv2Brtp0+6qIKk
5S6KlZA8aQyrYncwCQphj0Ktdb6if7JudTKTKnOI1gJkJ0QHwNZUPyOM5EIA5gAUF3UtHChff7Wx
IknW4iLqLq2KrnHVD8ABgCfwSruBpoE/1gsp1zaNcdKolqFV9MKdLpfvZ+Fo5QjfLpcm6u3AHeWu
WcY3o+2t3r2qsj1ITvwlC3zEzotWMMtrYgOKGhYoe6bzzF+H6KibOzElF2hLr3t1GlI4RsqXqJaT
mZGJqEY/VNg2iSrxXz8V2P49tnbqfp14TIWgYH5hDBgiuDyoqNjtu/dlY6eCvLIyWSgnU/gIuAxS
q9XjWyamzsZN/Ynl5zrGhsF7BjLMcbGXxq4SVu6TxB9v9RmQ+5c1NjaVheB/ebt/CXGfIpmFwNbk
p1DLInqzXUpHxl1RCxGHlGLG7hNgUPoRtW0tQ8hwIPyHUlwS9/F8opgqZnXT2OBCtbsElUW2XzbC
Uc8k84hlofhMUP7cN6zbtFyBCYu7ryHf4kaJtw6qNnYdXE5Mw5biLlK6tpH3g+hrTOzmz67UoRgp
/dD1uFgxfne6YBVeLVs2qSC+DUUuZhqUhtZ9YYmaYkxpToAtdJK4rRe5/hgHQVmrhC3PTB072aec
hOGwqN+Gd6boVjqkrDujzgmVDzZ0//NNd8Ekk19BtlBUn69nnEsKzRvxu0CO+oxOj8/2yu5/HyAv
1LSL3sbUH5FrUE0KnuqNyFaKHclX9AxvaW1iuX5tjPby2VYZwdgW/v+znK5TJv2jWRWbm/9MrHY7
r9MqLwlxDrtfl9PPMDFSXxremBln34JznSFH4oglgmYVQZDCmwcpOapvnIazTBH8jqmL2mvEnusP
xRu9TPqsatbM5kXOunu2FGOO0bciq2EoIkyggx52TriNGUdWrSlBpzVD1gsKHo2UfazD+EULzlzK
44+zIiXOF3ne7pJClfRH1xFYWopjWfUC1nZ9dk5UUmiJhvTW2mr4fsTapDbl4Y1IpzDL4BFfKeLp
ycsj8k2ootVJ5+ujIcBRIOpz20fyNrqqnq5L1CFL1x5W+CoOq/D/ZEKjAZZcYsc0LhKYPIDcZAu/
rKXDr1xQppRkvQZxym4achc3UHgLFWG572NhL5k8XtQipaotT7ZqwF1s5eXeQBgupdyqkcN4c32Y
OrqAJ3EGDLfhCUefJVl2ppqfj/Azf3hwMTBd1WX7EtkakuQTDYulBIOSKkAILadgiN39HlORaoXc
dE24FIN3IzQzngATVFmDNj/qSLfNKJEI04sOU8jxGK41AQWAPQwplYmZu3B78Fp99CJ/kHGPqggW
091Est/+uxgZV67/obYVS1uJ3cqmfuWBgGicdpDy7Fn7gI/yOeeZWUWhRtME62k7AVMYeWajKtVO
b6BHoVYLitss4N2jDfaoGDeAuMFkkbjQRfIEGHo2LcPg7ZxIF7hogjf02b3T9optrQUQ05cPFX2D
D15BOKVuyKfcHvTBB9S4/agIoFbL3wJrv2YFGp930mJfAdyPqya+u7nIni24E1tHpc7VHijEeZxp
zmm0fwPrSpDDRRET9aU+5ef5C9J5l7cgA41QRUiISbeU1lfJVN8KtB4R/XR+8RypjbrGgZxuQ4OJ
KLyK79EgfVXgPUlhbXIguQ6dfOeIarTXI0FWBzIsCARLYiUfRRwR0LM+hFPDiKw69G1F7uASmdTb
RxQpuW4SSImHnyAo7oKvJrboSJxYZghDyIM6QG17YQrbbtBWyphm7uijg/fSD88bkYEFRpeRv6Mt
5+qvzZ+qnNW8cBcLGG3xmfOYcNpdXFqxQmDUgApi8D5gOXRdQJQ4qejJINlNvDmiiEAqhHdD4bxT
OqhOtm3ripI4gv7c4l+YxtSAcNRuj5IRpxs/YYqyFkiPlw+GgVmbPI/66YWvNLl2E0VoTEYYZcFe
ke9LALVOPCghUdIKmn5vCdv+tcrhYFS3/f3pwgkOFpsZceEVV6Z+oyefGm7b033GJfI1IRZ/AuhK
PMEPRBA39JrQ3Pb20ltFy8ZuauUzOVQjGcXWmK5jGugnYO98y6T0+Rzmn/8vTvt0+9tyYybm6Vz9
t8s1OovrdJeQp2WACRR/llzJU2zC2hu8horZvD89YfIhLAE479BRHrgV5vBbXF2L4PmUX9vmMkHh
YIBwPLctmymjTrRJw4TP5Q3xLNQZZdr0NC5JPAoBLSr1etSGhwk5lkz4I2yV20KoRA7qCh1MxxOx
8jTxeTHQZDYlvNggLdxTDIPSi5/dbSUkMbniXqy4lzzLT05AR9xTTcV0Xr9wLS1de2CHfpWocbdU
VseyKGZJ/3QwAb9FEqqSs4WYuCyVPMVdIS+7DpVtRofadFtvAVfD6wxERq192J8zV623jsJr0IMM
HMD/FVdZPHADr5yI9Uy7wQhv1Z80Qd+E3dkl8hYLjDHjnjf6Dex6GJsyU8AMAXtO6gxR7dvPayMK
tNp4LWtdlByzIXRarcbaG3Rk3m4qxGEly6wJO1CZi4yXaE2tW2k0S1HjNn3OMcuKCQwRW5g+dCh2
bB3zWraFYOTT8/weRuAYdKpTGswz1rxSnV8uvH4qhcQXtX8gWC/9n9KoxHfKbTLdKgjLHq+v1eyO
w9tBWtKtS9B+6byGZ9eTOKcnN4wFl89vb7VXdmktz2MUo+Du+REZzOFFi6SmG7GN/GPGdBHwx78s
MZOx1h2erC1+clhqgUF7J21CN52vNI0Z2jc17JGzgoeZbvjzor28+wVJiMpln7jgszDE7TkYDKjS
qP57nj7ZgL62/zmEH5quG6Mr5eCwRNUFoP9CQY64pJgITpBcoX3UbihvF3H83mx79Ca8YHdUJkFA
2hm17Kfz9mHaiMncfjhBOGW0kHXq/dJkBesBy7KQ8V0ZEmKbjLLuROniMt5SBAEePrTRNnRjiXQn
bQXyTKpcWG6PomfSsuO0+kic1qARByb/G/DDBVSmJdnkUEhixThUlht3nBamSbsOdm6cbpoarAX/
6Dl8DjoxUm/po0no1qnvbAyUZ4e6JuV1cVuF4S9pxBwvw9/3xfA6DYbwrNQr4bPftcrwv4/FMy8N
pg52hFvXUbjOQmmiKpBktilPoT3Ci+T7nSMX7LjVDAxGe+35+MRNyGdAAfB0JVxDwfSPutsTKSzJ
Y+0dwf9np4DiTp9CGC54B/mv+cYXQTjnru2rlGobCmBIP/ZPsD/CgfUvF1mgwWXAjLY7xVqDCTZg
MuVorToFkyvNd/y4b3wpI+XPDo3lvjS3OmbCn5Nflf5RM7sgB1g2pKrqOdkWM1/piYIWjLvylw6h
Xa9gh8j4USnRSv1u35zyda0ttaQYK9MSI+xrQPy9urj+s9fjRCSdIgv0Y9nrPQJJR56Y87wuMYa2
hq0B3tmyrCu+eEI0HfvwKjzYYsRR0g0xMgizFpkSSnrAG7zwELvhNgujXZ1bwWMOy+MyWJ5cI9wH
ZxW+7VHmQBZru3Zn3g/mm6P74OWFDSbqMmChnhjrSNcmIboCO6AT1/Pg86pFST/q/sOrEL7l/wlg
GujEouVKlLsx+yNI9WSqsbuQXYoKtpixQTEZEe9VJTcrm029YlqJKbDgIZAD23uD/ZRhyVn/t9na
Gqj7wd2UYc6iuJmnnjjRU8/zqBSVTP3FN+Jcxd8VI+0CLyOmnIEbU83Nfs1LOSwvYiPskINJAmRD
ECGENH5u+wU0xBYckuC+r4a32D8ikgvHUQ0U5nKt3CZ2lICr98BTlONozAddpSgzzI0sf9oE5ADI
IaSiPDlrGvZ7h+TUnx+CFjIy8NlM1qCiBYrQ9OKxKUlpivxpP9bCqqqnJg3eGP4XwPwqxuZu+u3e
U//gH2xBPwZRa7ndGhQQcKT5KB4IxTwpftVrAmY4M4VhWMUu2kgwA+aXMA0Z36wvu23TCNYKW/zQ
oZap5bBV+YVA9LBhDYp7F+zJSeAdefp6HrZz92qfjklKMVZ6rfHiiTo6PENJ2hWi2bDTra/EleRQ
pHRUTBK6Z/u0NCY8zIgf2d0wSScf29nL9PR5pUr8R8m3Iu1C0y6nGaj0u53CFoD0nIHUag6gjBvD
JnvT+Hr0IhUV8QIprptlFTfwZNTEzBZoKW0JUC31yjnG4+R0nMkhs5f4UEpOI5cXMveaf1wBvJ8W
TlsxpCSJbiD+4317relYJC02JUs9Hmz6yVOVVfHah29Kp4XxM2crZmaJlIgcbVjFVLW7/o3KKIgl
0ZUzvMy/8ThJHf9+UZuN5MysGJN/2HkvcA1692usfomKJAAs8UOoe+SMMQH4h2CWBFx10+sVUe+7
I6W4ZwllSF6M/T/0rC3hYfXpC2AeX0SeYNmFxbcjtEsnBcOlPyFGraqCPgyzUZ1cf8KGKiV2woWR
6NKET67M2QwNkPkwF/a2DY+Hy0mDU8n9MVBllEZ+4ZPNGISHfMnpsoZ2tr3w0jTttYC1lG7Ys5/k
AyO6DaAVd956QYaxPWJd6tXmmm6ra+4wkq8r50VcrxlntgVKPv6SrPbHCoeNqM4O5YQSA7n91GSg
iS8sS79cIjwTXoD3ob1iMxTif0NVhKUvd+VkWDsmnG6xPfQ+2r23+g573k2BMIyXlVCb/Y0KXElT
pzhJPHaVyWgr4MJeuqCAWDTQvjAtvFjSh66PIDTQTSwXUBl3c00e43Rei39EUnWBUcRYitygr0DI
VYDpw0yISLH8q5+2bYSpMm86hoxMxiYm68TEmcR/lSNYIeaCsO5VlptZgaQeu2Xg+DRDBf6br3cx
Ooq4ARZsHPVejqrJJIj/t7GWS4IGmMZorPGKYujWr4SkEYaoGmSUXH4DfZgO0jZpcu9JKD5IJ/jg
75DrTq0XZpQGfGH6zTp2cwVJJd6tHFhgGHLQSTxXVGcTTmGB75gc4veVzfLbd+th74oUI1stbr+A
XF3NgO2sEZ6UVN+L9NV0Hv9kLFSSOCjhm1KT8NkLi/9CSqvNxwOa4egkwqA8oGlA01IlQvFcFc64
6ZmEf7pNjVK02b2wI3zsiubvGB/U0cu4pyJbIyScSJJdIShqzwetWpe501qDUmrY96tDOaICAe2M
qo+e5H1YB40+GWUI4iFQMA3z5DaM5zHNgkTdgNt4t1OFCkJ1Byb+7ZJoYBOHjRVkMKy/gFGFQgJU
2sB3FpHUC0XdilGECg0ZxGfa9mcOi4Ibl3fmJiMxF9WtcRg7rPpTLHE+yV1KIZRLe0NY9KmsIpVr
YOvJ2LELSziiRZK+SGnvE59gN2ZDAJ6NZE0EX1nO+RK1LY/+rzAjRtfgtU5Rq8NAtm5bNb/X8GFd
l7VanI4mSoeF1F7ZlJaUOL04BPQcyRbRRotR3yXmu3AweUuo2iyHOUOit+e3UrgNbkC8mHIR1fCb
Kv/CoLsZsoa6KdTqz7EapSoR0oKJEcCkxN9NnU38r9mHBC6RRybr7JblRxZll514/IVL6eYqpWVk
oME6mIjoY4yyKxaYV5Ex18fFLr1txfoW8mqu6RMIfFv0zI6S3yxlH6Fn1YVGyYqT9iKjGYdKHBD9
xJk/MMOkt+v1DYjWiWkJyjL/SrjB7GkA2JmQWII6QuGZtdCFwAJWkNk/62yjM5BTrDkZbBtV8QjN
EWKasaYjWOIFJxFkFjY/gIcLVQi9q0cfo+Wdl2aePZB+XUaRWhb+4XaXU/zcTH/UbSOJMGioPfeC
2jcpX7o9LirClvJ9ED8Gfzy0PNv+5hIQJjNMBbNcfaT2NAYGJKW1bmBtomPTDuIIgH1C8fIK5D9h
4DklGuVTduOdEeFT/gMGzg0+hMhsHNK+jaNx0r6LEjdXuswGzjp2D5hvJo0Gxu4dHI5amv4xVURh
vNY7SgRFdDgHb/4YdpQpWiZ7Vj6oWdkV13+MdghJBOmu0anmoMDblsHW/1vV5MJyqMybtqAfnKqY
JZBMmK2AlYIaRL+SMEBD35GnzqSezvQk+FfsduDlZ5vXNjF2JDGTT5uQh61dEIKkOKLqSVqYtc/d
IgdsewvsgdVJwDFPZME7v1MtsN+xCygqIvWPu5bpX3obBLxEuFL8WxJzOgSLznKWF0DvrjfCKTbo
u+ZdHpAFCSj0pYAlEA6pwsOZYnhN5QUiBM2KBqqHcCph4ObLgXOs7gkMbh9oc5ts+tdYbubVS+pj
kCl+sNdcqTJmJLCboaubJuxFHaaFj7cS6nRpf241C97Y+5RGv/oODjK6tK9f2WgQa0BNI6QuWRA/
+muID2rGjMhUHILOywlGyRW2H3zEytQLDDWOzDLqRfJLGB69obrHGoIEE/IsrvliI1qUGnMwn/IN
gPaZi04EuXC1yxanmgo10tpEMJgAdHEM85pOJtmZOPrzmKdXzG4hxoSc50KdEvn8hEVYFWS3ke4g
bofbLPj4MkWyMClIn9bC82R7pFBzPPdq/NkJe/xjHJCPOp1pwErHO8jbEACcDFen2oUubBkf7Vvh
/Qqm62wYWVVjdaQz1lkdQ3mQQphA5xUnyGjqJVS3dm4YfSrZjyp9d+1VEcc1GEiaG6jeSyR+CROH
DE4m+GlixHNN4Ogpb3RqMJJzSPxpBLRGTS7B5r2+yIzoi4ffnA2oDdfFtTvFaeKw5O3hj0AYfKwa
Uppu4JXY4IEACAKfnP3pbHE3qrS5owQqnWRE4z2kRaqWJnXs9kYA2WRSUSwSzE4XaJ/4HsLhRzwD
vozPiHqsXRHv2gaE2ItWzsTfVat4MQo0lT/g9WD8tMjD3We1TH3qU78k9+pOGSHAF5FGPePksdcU
4G1RC2MvhPBvM6qj800vNb+TTm5AC25YaEyNzbi9VER1No0yyyhPWUYPY5lxViIMNmbMmrOGkLJF
S42VBqVgbCEyu96y5RhJLZHr5Jn1TtqJ/SdmeVKF2boMdBJ/YsVU4wW/EB4gtBckbMa6Kq/ccxJC
3d5AxaFh+Fi/wt0jsqSVC/ihS0d4dyGr/itbNNk2IKVyLWGYvn6bdZl2VUqo8r6riY04RCpTYLxN
k29U3CT7+ANOFGbbNbIr7HwkRrBDlJOtqq5zmfcQilKF+6dpx0mBJJMA6vP+V7PA8So8qMdA8cUP
RW8hmDO8t16pCGpt/GXyjSe7i71SYbAtSEGCPi3Qtni/EBNExb/+ahRdZ2uwAAui/JBb/YUSsqlh
Wrprcrz5ChgztKB9dUgmCaCYC9BjKRLRBcmfV20k7aXwb6BOHuiZ2rfc+KD0vYfLHMVCM1juXK7+
6STYyeFyGMniqzbiuPI9Xj75lIEK8SPyTxgaChVk21MzxT6jG4vR55ifeU8YwDPUaU64brYuuMyJ
SdfXbQKo28Y0QIeOSe1hPjposhNiAjL0EMdRETM6SBMxKuuer2ZIZ1iOhAv9HZUAMhbpEVELoEXD
RyiixGPp8dijQGX0xEfMkhohbkZyIx4a6oVxl+0B/BbCIp1kCIcTGG/7EG9mjrhBLtV3I9LDe7l7
rqQmNB1zQyIDug5nYX6T0Q0IRcjDQOFnn0VeqHMeXe5/bVwFBXefHrbWX4S/g0klYQzcp2IbhtBG
TIHyPKqihjNpTL5QJpRljBymzNZGUAP39y/nCkEoZYRU9aoSzGScrZ5xo+1wwUPdRWJ5WnmGWUGq
8A8CN89KZvpEFMa1+WCN3pWmOEQJCCNs2DEjTQHZzflt7Eb2mePOYHTr//GXr8KvcElmW5qaQahi
EG5Ndgf7PgEeqClVgLQ3uDYwstRrxdFGQkYpAPYaDbMIWY/xYmNuhR+2hdGDP/ZeOfxkaP2Jlqn+
Qg3S7vqg/8J8OMfgL+4SZ6xj1hbXw4u0SxVicVwUwsaAvqqxNaFDQLxyEh/LBrLhwf3nHc/meEpD
C8tcUA4+jChICvzjQ7tqrXAvfPXeWAfCQR8XCjhhSLmx5XQem2gfhf5XrQ/y1z/GEfzXLXhp/Z8s
ljiiP8NL21Os5c6Hj+NpPyEYdLnwFpO/XfYfWikHW3eih5dp4+HdXvEGQ5SJOOcjrxG0ak4cEGNM
qqwkFZEOdSNJW5838G61mP2zBetFq1knz0327bPTqxBBROqf/LlVf6hubuhs9ntwY5jgMBl29Arm
w+v7EjREo/pjBRGaMo3G2TIMdOPjS0ga6U0UCJ97h+A6W0OSMDJ2nsTerJSUIb1o7HmZGirk6rVe
x7PVX4G7bxksotZ7fLf8zn8nnZQsKZ0zrWQkKF7sfp6zbg6NlUya9Q4zGNW/Yk1BbZ150ozWNCvv
MYj4RED2UEyNv8ZVNlz9ikxPAbtLcGGZ/GGSl8C4z8993Cr2Ezn2JnJZu2GrDbM5U3kKEnr+qJ1t
PVR5GxcH5kis2S0eOp1NbwZFhZQ9SVuryI31VTMwT0wUY5uaedTuaT2N9iw/n2JdQVori/QdQjHb
l2izDUDQ3lVqwQ9lKVTH33i7sd2o7I66Tg910OGIejKtcgwOsOz5TVjdKvTv6CVlLR354D/MwcNh
VL8EIG3E6FrXGj944sV2iJIK5JFwmLpQIT8pjQ4ae8oSmHDXqI6yA0sV33x22IxRQy9GkYPALhXa
HOTBDoJpXtYUdTOmvD1Y9fna1KsijmqIdu6+CFFY8oRLLKtFuKnpAKjh4Ggkzb6q3cEYCcxI/Prx
2bPLP1JpKAqWO3zdpMwiMnhF9deQ0RAQYEpEtCDwI4OVC1UmbSZmfGEAlzVNNWHyKyirfqzrOnWn
3piesEuXGUZ96JHZe4JTWnhK1NWUMSM8B3f0tl6We8gR+o2l6WI8HW02ofubtgGnbfDDOZ4EQCiY
43MK9v7O9nQwpzR642StUX49SacN2Wp6OoFPeqBCVqc7sBEpSpQeMTusi6Mvr3VIyq/gGQBnQ3RH
ZC4WAuUaFvE2e6Yjc7za6iLDtdhlzZBQ7VpR0WXepvZFJ5DtdmJpKhS4376eqaaxTHITcYwuOyXY
SXZv0DiDsJkba8RJod+wViz1mVa6qHdkNp16CsE8tTvOaNEZAC99RcFtxULhPyGHKuTUl22x5a5J
94bkQUU/iLGuUxberc/UElBclUp2w612UbKj5eSoPQappyAS9TB4IRsPndeqcjAgUlg6wIy4JYcP
vY62lazyu1k0eVzWps6R9e4SiE7klZfgJFJ/g1qH9IwvFVX7DKKrU2CC+8UhlNpyYVJQ+9LsvXbT
pP8EhqIAwC/ISXbyQRVOPMmAI0gF7zr1Yc+oOtLEz1UFStsfVVFe/Qw/oumlXo66Hcjao1ZQ+26T
EK2pBFBO2DGCh7o+4fnzww/C14O31JKakBcAnRoN1kMkLfmXZ6x0HYpzbdTaCKqo/U1w8wEQQYOK
j7c2bZQ4mkywu898mruTM5dN38VgVTt2VkKuFYsA9qJadI716p63EmnNFAUnBGo8WWIMf8fnZAhF
cG9RgyfMo2K4XdtJpPe35MbnzuqIyHrITcFvyjszynBJLg+J/BFOcu0vf6Iaru7G6+GVSFQr3oke
EFh7n+7oypX3RjEkmN0zG/+XHUGVNHfzFwQLFSOOZQFa58I/GqTq8baoS7aIr9x6K1M854gPaYLu
Ploj52m4LIJKNyaNWrupQdo0LgpZjCANQNq6TWe5dy3l3wHY+fRIDczxyqAToBAvBvRz73QXl0lV
3+OFd6rHQJB2NGwbdPUc/SzuHziwz+Lf2RKnzE5EnPmqTvPh+OKPtU77B+vtm1l0BK77Ed6EoaSV
GeFoDGOlzenzKvPJ3oAe8xIdpbuN1USMEY6HshoqDET4vRxd/hjS2Yox0x/TDFwqcuwLUG9sYHXm
DwRj0D0hdZ5XWkN0rffEiIBczTCP9/kxlDshlnCOvCyrGJI6X/Vz7DYU6bBw0wNGnXcDFBQt99a7
2hX5bzC3duqoLXwzrKZoY63WCJRYQWAuYU5ZA29rx3c1NfxCr2wdP1D9Vp2lu+KFf7COR8f0TmMK
Elbs8fPxI9R/PXSx9lAY5tLzsi+bW4BrR/D9LMZaAkne6AjBf4o6S8T/RVlAE6QuK1p5pqc75lT9
R8PKqXreDn7iJ2GsQVbMP0ko/zmtgwl7DSODnF5J1KRJkuxqJKTwFVcmQZbvZGPbmOVUeHUy0esd
0tQEIowvEX/4X4KrNkFdICIPKTGHb3Z0OwzOXPp8bdHEKeW0/Vpy9fhm557FTVFlmuICphOIhH2H
Ow3zVgkxqbEpi0vD76vqG1nE1oIJ01bq/sA0thwRNB6sdAuSHTEzbdPdq1y3abiSEf2aEooGQKDY
Vl6DFA+fSXfYeWhKa0SW0gE8lsZXDQoToqzf55zV/GwZgqDIVKVJwkCxkbDEK7jkxb5kiSCjmX6e
PwSfvIHZMnO6VnEC7+/lsJBW6KrlY6KUHsWQ4ZDTpePMBFAbCi3IqJWu1b61NRD5tFgxtiXgJX7L
7uembMeo9AiCJ0DVczbRe2orcuCGqtc0OvleC2HWMTJpQaQAxPimlTwtPrTNYwTQIoz5804CPVnm
xUWBeMeP96E8jDfemQHkBOa7wO0/y5R1KdFa9vnGQww5CVC15j7sMXg4avPiFA4oRTlquewXO9Ap
aJ54zkg+URXhOK44AEQupIDYIfKkRY86VnQv3YFFOUOpcLn3xWLplSAG9yaEokT17jsK1nihaEBD
WsR8txFyQWhgYjlCX1t1/k/vjwdZEq0eBq/Sl/7jGMkT5XkFmUXYL7w92JpV/Uf07XCs12FB1c3s
+YoqeUbboRjNZnIqTkfsWcSS/Q/bxlQvTySpGN44DerbVS1VGhtOD2h5IW+QTcsls5gBs0CEMflj
qC3y9t2cjEiCEnfDtfjqxyXxLpodCgn7cDipkXn+WpQerugq3oEqTgHzq9yUQJccJB6HoH0vkdZc
RbqjInEcJRrxPr16NMeSd1RyyqoBhoHV2lLrFjSEtnu+y7izoDSCXE1uVejF9h9CwdVkL7kV+HgV
lY/Swfxh9wsw0sYZ/QtcFKzGgqahk/AlvsXi0A2pwAJyGAuKkMVw6/iHaXjLXwA2nMK28Ut6Kbv+
wy2mgvL/XpKkcn9i0yduzkXSxCGG806LCVhssAIg1M65tQfoEUjxSyd0jf51GFzocxVeppUiRx/R
EB2UDBFpF2fHpT5Xpkyr6RhLojtMX1y7OXV3EIQQLOdhujMKlahwa0nmUbHGjvslTI6dOjVPT2m4
pA66k+TI+0cwNWcDg5rYQ85aB5xTZ3BxD7B7wVJyL39iYNHeFpD4D2wpB2JdX0NVkJHO9DR6rOPx
3VO1q2Dvox6N0XTpvVzflg3nCKJOMWvP9GmaAfpd1uk5tuLq1T/oCiE2ngc3NwjI84lJTFWR1BFy
swhAdxRBhniXXOfqfn1WnM5OYf8GyCXJc6Wwnd4xz8U93ZmkVl/AInf/Deul4YyNSHJeduYFOakQ
B3J9QmMtfc9TApuZ5kRxtIFJNcxKTn1t64x2jgtkKxi21PNcGLGAyzWA0pTnoGMcUs3SUAaXns/t
++ZgNoyGnx8jppOTxMDE/Jv7o92GXTALgSMBMImQ9VDSqPIgd4sSUykJA6kj/ITVyGZjljPJJDX8
/hSBIVc2JiK1DmKThLN2eTCO0EMnBLzFsDGxkfBxfCuwrzsRYWd+g6L+PMJxHzPhKNJEev5n73/N
6kfAAWviIZ0ZAOp5P6Pb58XCEoC38kP6CppCrXm9bWhDdsrFY+Pin2k1OCPCTX16MMy6k3/LTfXl
+DhvITnRPSae6/2iE3Pwu6q8qPcSKm2ezuTk8XN+QlYGC2yRf+2kUi+gAXlRV6AcDyMAx7YR3lbb
ov4obf49iCGhkd2ZIfwYzXK0CCfolY96DoxGypmYrRwdBNeeucQi/FNNZPTMCZNEqAVwFxyI9f7A
gk4QnTkWeCwQjZ1LbnhKNDFKXVn3DVgzc59pAnlQbcAcYKUzd6fLLoraaUsu+DusztqlPagh4puA
RDo9KwgTz1qkjQahjKbIFQNZDbF204p69QIsc4EpBGsbzSaaKNAcX88fGaBN5Hqv9asu4jt2cMz/
ryyk3K1vXGRjZg1p5cUGtZK1azmIZtp8GQvvXyrrScSQrD4vuqLNB2X0wjV1lEgfYXLTUiBzseN/
ddAIhLeilDiw1jQlcgLhkxYF64zEAwUzR202zfwjVJAuasU7to7055FsYr8HsEFEJM4TacWDSc0F
ZI/Vrs1UviChiTfqtKFHSOW+fOzw3/XNIGqwnBX/HUTU+dHDzQ2AFO/2bdomhfCACLU9ewuA1erL
QUS1hpctgnjXw35NzcnvP0Wcq+hZj1DqcuMj1umg2PwLhpwCJrQGv/Zt8aRzSmiujCoh6SEIqtiC
rhDFDrqJ99+N+Is+wqyffSqmvV/yE3/ELop6bnuT/Qgu7LK9ulbSXOqqaEKTBUtP3GjcxSQxDuTn
iIoeXyTglRAyhNNsEss+2W9TBs6bO9i4OBGL/UTVoWAON9O5inxgxAnj5srPcqWjKF4RH+wHCQbk
/c3fBUQ8m+ofX6XPAxZ4g3RQPzuyO+KcTRLxKXNtKLmuxXB5GCBNP4l81YbUz5Fsltf45WlyxZMj
ixFxYlFWWaFAbYcUiGIKHQC2qQDdokDAD3dTSnRtRHEh/OB/TFniGvF0qTiyexDgENKzCYksTAHd
uleT1fl3P5wItMBy7Q3oYFouPfXyBkBNYjh0PcY0Q10WDCHqqSUTRAlbRnh8Tk3+rabDCwabg3Tr
cfhp7HH3i/YCe6GZPhARPU2ASZUIiP5JqfpMKapizsCuZ8+jpnvX/OCG0HqDa7B/ucp/hMRXfegc
azq3y1IGJgx3DGhhTB2Puus2FsakZ5Y/lNtR59QV4Fn/Xu5sO2335Jw8ONPVZoHDp/pYDV76ijIy
bt5fM8IvsNHZlz+Is3wfrKzUWh51yZD3vIHGclWy1yEcMQjiezcygSiJ85jQdDJ4QANru7Llubpe
9SFQX6Cx7PWQ9M1b/YPHOKe++d+6BPtwXYQN3Se1SJtn0I2Tt92Hes3vrFgD5rYC5eInazE9EQ5i
4PwddiuOgS5uAJ4vJH6bN+UKsTxJQM8GzATKGLkPzgniBFapWMEm6Nmv8xRomLwyAX8V9xiceYGJ
bIj/XaSSelWBokq8YEC5oaUh8wllvw+JwKu8xVZMGxH0QfDCFkmpDPDRLisHLQvwSLmuEvFCXmXA
peBL1Br0ikCumEbMe8CyPQR8yZSRRU23bgEy+xUS3KejLE+Gqk7K3IMn5ONrDyglJaCd2ZYJBBqv
KS7pvzHd5UkfSAzwsy2iSn8covyeiQprMAT0znVkcfqBJEZKZpi6KKSPNhUPy0ep4pr9j/pE6gaK
/2HKcr05qSEzATWoiPhDZQVO9Ak4RILQEG71xOJ5nAfQRlkAdDQoOlZhvJxeoTtV0UoogGwlWaYk
PT6Wz+PetIzCGsNQeLU/kM93GUAJTNbnHkFH69j488oDHJslHZrZ/DAK2IC0yMlq14PtjtNAGfEG
IflYibBqopEZnG6xBSZlY1uRgESabX4EUJNXQ/tfIL0At5f0Ys3T9Le+zjmszK7DthKVp9vfWnvw
2Axv7tJDTpyYiWy/A4NQaYYotoj2FphtqU9kMJjIN4R90Mkq9rP2dhoN17pLx03SMT/HGLhBMDH7
izNrmqj4oLBqsyBqkEpXNqLpS+cJFfOC0dY8UMQ5HTI2j+0JNawdA+Y71YE2RxHVgBPuVNsjyFvF
r2cIIAb7y2TJ4JUyvFHnXi+T+0uzAIlFiftXLh/offxwVDU0UGz1AY+t6U/oELTQqHSAkAUn4YCW
a1Eu2MnZ6a+psg6SSwxQXc/qhROwdCnZbVyZpBbvGRCIYkDcYfnlpqNdYSIWZgbOIhcKWBrTqRyY
dlJtkL3paM7JviXvNt+N+Rfp/4gbnORaxDkVWiPFKUOFViDH1o2R95XWbr5wuCI9UsuiLiNKhgx4
+DQCc6CA6qPKulXvjaD2MDd3xaenIlWjwBhSL/pRYvTmBhRU8GrFBHuOlCjRfnEtsqMC4K8JW4d5
Rf3wL3HFUHYT1hN7Gj2i8HXKevjxOz/ruNKun5ZuVV+JmyN+ntPB3zz/ohrHyzrVebMpF/9DYTXN
Foca/ba6n6I+N1betw7/ovXgeNWMc11VHwwcHBEF+3xSuLatmUUElPul9rPVQ6zM7t6cbffTxpha
QJ8ZnPuxb3Vcb/B6/objolG1LSgvYBONVVTRNJX1io0Oe7vi+qiAIEVj4j1HwApPMvF9w9SY7lq+
TYBe5pK1GfNN5EyEyAvJxFrMFgn3QBrb/GrWDitLdCqk8TCf1bk/yU8Z2PFwjcS+AqvOOlnjBCyC
dLcRE9i9diULekzzcE1MYX5R0Tv2naz4Wo83hNRpYvZLC7HxAYE202+780R68vjCg3wom31jkpdX
/3UMadNq/Dl8bzJ0qdZRgwMKFLNKq2u+mUEADm9D+xZof82uZ5ycvr0WxlWErnsRjxh/33lZg43C
bU7OpxYhMfcTHRD39ICGrZwLGN1HOsqB0wub1qnKYjSkX9+1u1YAUKbLwwCEz+8CGL4dkIlEvqwM
qsR0gGzU+aaDxcUelf3KN3TJ8M6A/lC+7pwJbNMLUEwGWXNUj3YJVyWonpFzDJtOa7ubYEcXTDzO
Sm0QyEwl8vy292LNtmWUpzvHxh7KPAZJwkWlGjiBLK7cyxGIDDHnGMabke15UKHoZ7/LC8zHSq0Y
kJR0zIj28TevjQfuUfzYRpWzvkGpmOj3HdTCw6VMLcr0ZQJtZNGwJ4C/ZoOyJnFsUxT5vJ9/l26C
gE2iJMrHr1znFj20BClcyDVTzstjjtOMjXZEUs8KpG70MjMvaBnUfNSgFhtVU5S08zSAOaBvdONP
MRuFm5QKURmY/OEcazsdcqmrpqctmX8kbBlFsyKVxA/K/D00uDykOpOLDUUa5Vv8NXy/rM6I09Ik
DZPDyem+BfuDFykYclWfd/f7Q3rL+3JbdIqc1W9+vmZHEnjZ+Zuz51aUnBcxFvyctOT6CvXcJhmx
CwMrcwyX/31rVEQ90qz8Is+r45fYTUYycHzZl126z+VnFZTBh8VvY1hSa//ioprrdohHPvgcKpQU
7cdxlVpENCJY9dXbCTwxl3z8srxVPX6MnG5Fs38cKXypQYI4Z+s05mlpLVia/l8FZr1souo91Ulj
C9tw0GqZUhJVXlL9H23sTPhYogQ+XuP/bI1mn6i3ZAyd1qbIHgEOtWsYz3ofVGCgaR8SUnHhTXLg
9/to3XLeZCvFI/j8evXPaQxVwp+JjPjPLrNRsQMJTFT320X6oC71il1hJ9yNlsrSC2907c5EmPJz
4ID6G4oH5YYx/OWqCXIWhB685i+XyyZ/foiG2Ds0oWbhK5xmn3BfWwpVitV6ns5DNVXP9y8bo99f
VY+3wpaFnaimtUvKL9DardE1fh9ABZtzZ5LaRTmOD1bBuP5G+zklMioslCuMYjO1OFNK/JoF6y6P
HPBVqfcRByTWQ7t1II8dixW7Jbsw3ZPdd7x2MSbC9Zlaiu6tgWs18F8gogUbiWXQRd/JoKmkyjsd
8YyD9pE4IvPGloAT6lRRpbVys4YDsSlJ+9BcJAbH39VWAhkVmlx/lrWY3rutobmlznX56yaaesHD
ll6xF5cJxbChuYFufM6qBicAi92gtXoGffxGod4gA7R3Q+4KXtoef24ikJ8sY3IcniYZq4RX7hGn
ciBkAvxWQsqepgrkhL+ibhObDcKG7lDXUA/A4lJFHC76UeGFafhCfEnB8nXL+ERsARMsybdqS70P
WnphPad7W0i6ZSOSrj7hYLnR2GerLTb93tKN1K/3a+7hx6yiaTxS7fa5Qxfj0M14k4J3VIKxKmO1
VZ5XiiYo3Ra0oQxY0T17RR7MPK4+JNS+qGBxC3bNyxUdLcN1p/cZ1Aijaq0GzmRG7buHQPddW9an
7BdoFgFpIUTIkKbelMMq9t4jROrKxYwBXCYDz4LlnIfv514mOdrDgIMAgZ+Y4jljmhTeGm1bRtt+
cujJD61z2/QtUpAk1Ddke77jZraDsdgqEmzaKWZp5/2d3vSs/bE+mPU9w602iAxnX0AMoAMa088h
Min12+1MBmlAanBcgpjccK0cR4o+bHnwRqvmzDQBu7u057XMSdVFS+He7tgJ/UtCEf6MfDmQ3w2D
58+l+d5+bEEN0/H8eRzk0I5VQUWu+eFC1M02XPMarMr2YQHfbJ41MwRJEBAFrYD3O9hT532dnsDt
eiv1LIZnPcTadp1pw83i2MtgHjYjiyGEL3owDJ/w3Fs/wL6MkoGn6Fs47qO9HLsaX3o3BaG/sYPS
HYRiIavjT52q3qafQ5wOfonUSoAxictKmyzrBx3bCLH2NVIAW5YM0c+ZsqirWXoN7hhtOycX4p8e
fzTAB+0lYxtXOi5v3n7pVSfrHqegpzmRRzamnFdkt1Ppolz/zqnvcg3//qHUbRBuPo8ApiOgv6JN
Q066CDV2GIKei7nOOSPswz6k8TFqN/eikmy7g+mwbpckFsuAu5rS/JARv/WtH3D5//5GOMUf+l7q
bcIOtfnwURRBHleQfDLanCfKQTLcvKpJcrDYQFJPY+lRduABxlAQ9PbHEe/eORsTfz6mbAO1YIu7
mbfPKbexyGNaR2/o72fVuYCsPExs/2jtaMsGQ70uIiEOfj9l7O/uczLwz1gv8aBs8GYAmVvv2Hj6
W8uYbmGA+P3owwivjfJxHrBBZ9k0p3AyxUY0Mqm3ElOFPnhcxZAbi22IJ4uGqjRHXdPZIUqJRcw/
xN+OERLOX+iExqqBadcu9bbC6JQfwcGoWQx6nw1DgWxRncUv+Z3PWn4WYeJ9enNb8vuA61pTB3HC
F29tU2cpyTYzl4W1elrXNM1spoeROmnE1hhXshCcuVfHRf17dOMiEwerjZkRCBxEuj75ZyoXBRt5
T/lF25O7asBSfZYFtgHuqMgJX75cy/3D+zAJh7OdR4a1Kx2dCgHklWRAwcb9iFraXO+H9TLsda8s
qQ+s/4Wwxcx9vloO70+RMO9YNqZ+nd60k1WrbM82fxSZHzncLi24rNd0Yfg5epqgg/8Ky5KNdj5t
9M4DISw96XG+CkFf+4hXn64jFqvzCaRQ4/eXNPkYQOQHN/+5HrisChF1UryG1bAQK7tIhuRbBdpJ
lVhPyDqfruyBzG8XDO7cWojDVuSNYo/zUfE26kAhZE6ijZ5jpmQvKOrctQfzzUgcxJb1C/b0F1eS
wXb+KG6DP+is5Z1uf1kYh4vZAgj5N1SYHRXD1xAA0AH7j35MinK1awYfpnK0MZ4/CQPT1XtjF+X/
MQHxbLuAphrHOjfOOWS4GMfsIs7tXteWS8brU2LdKx2zcDTJzhQv0K9J24ZMDuK5K1lBJ5/7yawz
g8mX2sQX+gReho4WosHkosNFpm3sZ4hOs7sj7H3c7S4Guo7z2+93LRFUG8nDlTqqijHGl0YQvpEh
RuuQoGwDJZoVb0xVUI7YeZnIWcpy7xK294CVRr9nEFH4W9JA1ZNLj11pFaLPdJebDczatrAQgdd6
cxBHuDLhYfqQiyVo6SmmLhp1KA8dMEqJGfePCg9+9fUZ8P8uaLpl2zcWiBtMPjab9bSjhGCBsfw6
tye+CQpbFflvZpFuENY6WZjIsq8my3osxddGb3+VNasa7HH2n/wRzHcpRP2aBawNrrA4LOOVDVc/
cFl9f+b4TRUEOgPuJAFye111bhkiXoShlauqYLjVWpLsCcgODDhGUAlwswmiTKWWLVYzybns3+th
ZljBvImW4Ub23JvEfemdvTuN2LIIdCcx4Hu77LBh9g1Q4G9/8vpY0LA81kQzm/VY+qxrK2W5Ynph
4fX0q5SQJni3RfPBZ4RAdnx9OpXXI2/xks0kDhvgEzjmMlG/bCCnpwNzLpJuqHxnlyWWVJ673zDj
mGqppVyrm5yD77hliDVmp0S+G8wNkXVKgFIgce74KbwHsIcMUY5e2TLne6ddFfk8PiLaG5jjmRnS
tBy2PBHAP9X6mAgnaGNFXnJdsZ7i3y+X2hyaE+qOc8TZ3184cRg1VqJmz793AOgBx0sOdNerPXgm
709nQgv1XSPxjBcU9VOsDDe3LbLFbxoccAwvwx90GBtiomjzvikOH0hiuzttG9WQdyjhqfoOFmsQ
rm5td29iiG9HhOSm2QDTCHQG70kUjUyK/yeM6wb1isdfnHTr2X6qFUpBfHPQ6G7CKsCuSH5uRh+0
aN54m8nwJ7p6BvUNLGEw/2HhhZCeN/r8bJYVVKQP2snw5f+EztQk9lSiDGzd84UcpWLZm8/I1FOQ
re4Y+ezPC05SfCaNroInWMh55PXgOu3T3njmldbK09Nhip5hwOAxC/+3lqnLLmvYk4FovqJVEpp0
RuZK5CWQ8m426Je9DByq2mLpxA58UL34Xy27D4djtjM8OI8y6sGWDtt0LCXwPmVn8F6YBwNUrNIY
FPQtJU6cRqzJuadtMsaZP9kbI4PZu+wzty5CHgyXg8ZLpLjgdYY0m7U5mM4R7KWm+t3a+XooAUCt
bm8xxBXI+T/RhrxkEDdERo1J54RBlubeIVBd3ZinPjd0M14aHwFX34lZQxZ2c3zZB7mm+OvQh+KD
t+wa+Xi94a2oaFx3t1m/3TivPSVlB5NEuXaVBs/ZKMyEpKTdrwWPIXmeI+Hx1UDetVCkdaGoxtaB
1GH2emDCGI0RvSQ65bX+PwkDLPNWHzK/Kj3exhpf9/GodC2Q1yxlk6+hNvtTSYXHiuftz375wIV9
yWXG4V0t7Dfb2bVq+xL5T0wJD2fmzj6T5miTg7EJK6uhlNsEAHP80JYow2+rwCq+IzDBGsxrjGsG
yY9aQl3ZAz7UmT/OK/MQq0i70UyiWZ2rnsN6iBMCcYF4aCM+qnI5uY0eSD3dmr8TgPdy03ybpwy4
eFLw7dgPnS4pMIvnOqGBFY75diCG2mt4WOS0QJy3+QdRr97J7bxjBqd6sCcTEnPYFSYb/msuSBlv
yv2vWOClbo7Fn3oJCh9BCLQgM9yBUJ0jkUdzB6Shl8nmD8PUNgeGeZK3g9q62zg3id+eUlkfmd6q
fvXL3MyXbQpLZCJDKWUAVO1y7s4T0Aix/NTp7/n3mD6Cc9qtoqSL98aD03ZIix7bpWlmAFiLxh7/
WfO3oy/7RJ/YZCaIp11HhDle/u2ssGSLcSF5zmuXJfRO0bof7FgkwCaIYXy4K3SfXxmRN8UtseUx
ti2iaz2yyqi5tVlnIJrPXjLux7daws6Yc9rtsWgcrv5KSth+fD1Rntjn+6PNtZBO/VwC+SyA9APb
VEmUSSSwFLX+oyuAeDCSZzOAip6jcjf9U1UVFHQi1PAwnCurSF7p5sFUhd4XWw5T9Lp6XmpWZmxZ
+sBvoj+E0rFzMyn6fujo3SYtZcOe7LITV8CkjoOQY0zPkIFIK1cel/20O2qM4hFU2uJKd+1WQokf
Kfo3rgKvvr/9RMh8Uwlxzie5fj1AM3KDpPJXIj2Np2NijHxxABJ7Bb6j9OuOKyOJpcFv2SEy2t3d
kBgyp1hQrsoGKWq2X92OBNxejA0AK4iWxyawISAxmbXwx4zUVLFtckRod70SnOCpi0JBPhNKsfQn
lLcPVUoLjLFRuA+gc6NPsrxSmIP6vt9WvvRn5NUJHDRYHo54cKhloMBHLHryktuXHqJMpQi+a19Y
641F4Ay9THDA9VyP9tXwTUJY5dZMWJC6GN3U3kUETNy3PQuJIOJxqQD7qskTJy48f/GvSIADqNiB
FQsp22jvEBN+g3QVafhY6fkBzX3FAj5fPRNWM7myElwSRsvyJwmhYEkyPe4TE2buh0NU1NA2yLMy
ke2fEIzRIzFrQGoswSgNU6bMbwgGj0g/JqXhw4/pNnzS0j/cFTduAwas0dRzUup1lwFL7MkK63Et
dmzre1OVAHMgcFUNxlXO728XROagK2GdiCtiiW6/VvYXPMXCJFiILsGlNvU7HW7FoVIhHpVsi1Bi
9gUU4jzK1A2S/hpOldh2MQ36uGItA44pR+zz79O/or29hkEzsHg7CWtTd175aYC0b4pfSrsUaogY
G7qdpgo8sQPHbQe7ZXQIwqJCpNki70kuVSZkxsuDK5AMp9XEVT5lG0Bg2DdI+uMHSH2gdKGAI7tD
JbkvFSP5/UxMBGvL0W4WIpqeHxPKTrUwVrytUuVg/RPPFWGQLVThuSG6x/BDkRlSVEN6kLAW5UA+
G1ghPUhrEKerlOd9+Gt5s7NQSG1HrwnQX38un4NFW1D2Ql27FUCi7v2j+8wTDVr+WZarfm/pC3bk
RiE3q+sIuW2c46WgdUzjpf3mEpDu7kv7X3wz1onePXEtL+RMxI7oTyoEgL6PyFo9/BCEAp01AjNq
wjDKq/rWY54eL69ajWSnddjnZUr1JWH3jeLEgHIIbLIjb/T+DdaCqOBXSkvf6EhVd2/v0ohqrsIQ
BCGytqkj2Esxz67kFfqLS6bIYbcG0phvOMVijxUEMjzTQreV3oFcq/iIxwjWH4DvnHPzN6jdbE0s
6ZY9lyFKtRFe4fobPVOVmtQGC1cgRIqIl/sir5LwKBkYySDL1ltI46kdLEUe319LYdP0oDrKqnii
PvNW5v/H0zpBHnzctV5+UeXBdpxhTPoRId1Zd3104a2Z2K01pL8fywHbrd0s/hGKPQ706WDUkuhY
XU1K35oWkTQUnLkvFy36iSniCvt8epZWdqe01R1Rgh3gQrhL2WzFN+Q56wTzCLsBWqGEEAiYZKjg
c5VaDR+GP1HCSomiSLYMV8FrchD0E67dieVb8ztE2Hx0fdqUjlACe3dvlNDpt2MmYIbR3vj5RBiF
5Rsb8XmRk/NRanMpnmOUbSHXBEOXtS4or7KkdptURMPXdAUk5yB9ou2NuJe7IA37b5NzJuODgdks
QH8VnIWOhw/NkSrDhIUmzQg41MHhDiimPljjLTZPddSQyY+tuNljXYpxce9cO5xD/bViQJseOBVP
FvHk+W+OD8+gpeQiJLp87ykaQs/EEdZzOkbCYlpq9+JNe6BinQWTfRjK3vYBmvEEuw0BhEjHZi9L
eFF5aDjgBwPedanGYznMWOhgR9kSmUuD01zGhMXQ8V8mHUJ3jdnQPBTGCrWUoQLy79zvqhgsXwh4
7BVRpbPgKGlEFQrl0PLCI8MPtop5Vo/kX39C4hZ0zMiZFdec1eKNrarpuHJapLxhoCZnVScjGNAy
hUoea8ohimp5w2Bbsz8ZtgyHC5ijfbRPTlrYE2z5X6q3yL9lYhfw3sD/VN+jzQ71wVwM/Q+ADWbm
rxufjIACD+UV2gnIDocTsg41iSrQFiBv+xtAE2ppidScbVkduLFyOkZNiBqr6jo37Sqtue8Uz9Hr
b4sETxViAo685RJbwtSzy5PEdwxQZJXn9ZSt5klNq7J323LQcdBujqZQxN2PcICH5QTF3ik9kIn+
01xq3g+yDayW4IZJPJWuATJs+p552cqnIGC1Z8NQlXIsD4+NmssMCyHJyouM3h3TTKNAOPcEkBID
oBc3VNUJXacMpPYk1aI2nGKUggkiavsM5VgJ7iMfbyZfM2RUXr74jpxY3AN2kMBB9KusTq6E6bI9
52IyIUiyMgnk46jcyYdsmaXB8ZAV8G4CjGmNLdxBcXrl8bFDfkcsBQXqy2Xr3dfhzHrhrPhW0Yx+
NenexXdXpn8FyKidK8O5QnZfuIFZg1gLwm9c4WFANL3KyHNC7Wg0YuntzeD7Zwp7FZQKLZTa0zNl
hogHPIXR3S2hGmgEFcqg8meRyXio8O8vD9HsNvXeUOiCuQUFDYPyLoY6VKrLHURXalsQ2wE9Hy0F
lcGzOsfQaoDsuzRHI+Z8wvRm7D3gOnxFXGKlNuu2fy6s/MiF1Ca2d646tEfIam2jcm4DqAtHt0cs
fQJDkysO1N25mayZHjio3WtBqAXG7xvN0FxVt22C91hBQZyooRYIijnUMXws1o1Zi0RoZmMhMEXu
Acs/74whLaZQrzFFm194n2CsfQhvRAcWNqCcBeHjrDVE+KgZAyXaJM7eRn1bjKJZJ4oFokehV4sN
XoYIS3Oc0Ac688B7ojLLhdaYh6ixqHfK2yta5RD/PIJvr8u/yiFGs0q7two0x9oPnmDGYHaq67iR
X5nscjpig3HIAIMMPZkuZV9/My81aGt/Il49rnNbwwIjbcUoHfMljhSyGqfrCq4aIS0nAbHe+5pO
qtTfSrt1vFiObVWq2NobH82+aTKegUNvReDOkae37VpJoGD3JXvNU3x02PWxBjjhj1xrpOPupPHk
bdO3SytWFvVZkbfKZ5ZoaRnwsjQBOIZiN7I7R1A/dN+zIBp4kkgRgeHcRGj3S2w1nwTbzgXg0yAU
xIGf1QxUUUZxfZHvuWvoUIur5gTHADRFVbgfpBJ6j0G4TkasVZvVx9weZECzxS6s0Fqdi/7sVtco
P2TIWZ02wYhX/qKij0e8kwdSg4B9VvzKlTCq5GrbzuHs+X7LZQyxFYk24we52p3zGKqg270QOMG6
gIofjdSoyO6EVVv/slqrnFSqy0oSCELh2yn90OyVsv6SUh8X6Fxf2qt9y2RC4K7VhENDSFgBTxED
yjzVw0PrJ1HZ5xUYls9NbtDlgoXSHC5uhvc22Io5kH7qdULIFxm647coVztrka77+m2u0lebC+wz
Ik2z9su8/wO14IxHqLG6z+Qmoe3gqUecgU2ujRbK9b1cyMFz7En64fMzHqw89VKNfAKbxM0HD5DX
QSbs2GbljnkiwzmLIDgZyq1z7a/IVseXTnXsO5vmPO8DLio81eHqJDtZN+AZAMppRuhKR1hRialL
2fA6I6kVSrDCSNj1zMMJFD7lsQG/yWIsrVj4/65rLjpciF7FWnok/C9cqtX8R+C6YS5JV223jAHW
8gEqDEKWA50G5Z7digeUSdMeA7cRi5nWqm91IB+6AyAgqBMgNtDcekHFAaPAQ+DbCaB6ldOzTAfw
7se3J5pR6C2juhC2G0lHkNgzlMuPJb2oBjosswWavd03L6aTPyxcDQ3OfGplcSwYxeZof7Y4AUx1
JghZCVSnV9MHyXEThkbZY42EAexP6kIUYd5EfGYmJ69KESy9pMPSRmURCG8rR/xdgQ3AqbZWinJF
prKOlUcjZIKbu99w6FYVSbp0cIRI6y0ZUb7cpBFg+ao+4nBD9AnhXbIKs8yUFOzzuxwY7mpVdZuW
71SFwaQgmy+r5qjnl2etCVQkXrQtQHfdSunOY/0G8leD7Z0wVHk/WWJQ+rZSie5tdIxTXpsI5B3u
V/B7oWWsHeil5t3HiBMZelTF3eavqzWhsxHMQ03Bq3wv/94M/HIe6RTN+ePKKzUEdeY7U3M+Zmx0
VH0tznk1UzPITiI8kN94jYTvz6/BqFL5EyrRLu/0gF+zrg1rBUgGI761WLLEnnVnDfbbNxwhuHt8
xGcuh7JHRHau1X/5wTPVk48DSysr2BlG1Tj166lWsKx60bvFWgK+M1N//6kug/nODLlG4qLCg1yk
UouAm6ICmHDNfPHXpdUcZayY7yPN5yzmGjo+7vP4UZprKumFCjDTC1vcIxlQ4GpfQeuhdfel0rX8
TyjPJqHOep78/oKDSEmwEufS6XYvHAVECrnC6rJgsNivK7rJq01nDKhlJcKX58l0RGpz+o0Yaciq
dEu6TEi+H0Zp1v3PNmoTs2jytyLufh2VQPNETJomv2HkJA0FDnqy4GRAg0RxuqBcuFP3/1xXNXkh
aWxyfiOOfnxfhVZs/GERTRweLsSUuHUH/MZugCKjxUVjnOoQkT4tU+qkk0rSw+wb8t2EdB6TcMi3
bJiyHX175+wtGotGtLgbgA1RbKwDahBsBCTdlz2f2+6r6JVBWGXNKpvC2Xdt4QvpFVTnVWikGg3W
Yg0zGf0UKl8voCcLCMibyTRzHWGW8O4PZDZCcBY5zvTNJSuRzUOg6kt0FrPIk845icT21ZIYGOef
sPzw8EubtwukPpCAVZYFlNDmjG/QZd5WO/qiaJKtfkIPRHi8QM77ZMRtTxug0Og2IbWVEjyzfPb3
1JMANonGFx7CVDxSJX6Ncq+SZqWYrU8awcNNrKu6BJW9ry4F2V9AzfkeqYcRc6Qn20ZvXU4Y6aaR
gdvTYSWaQa8BfiQQ2hT/zXk4afozeWVh4yLrQ6twvRz9Q9JnbDWsM04IV8IM7dbxTmNFCaIH8CCi
SGNMnqcnpMH38GfFg01mSd6Uhq8aabi48BpudNJL2n340ae5wFNBigPT3X2ePJ2lz5JfZ00OphL4
OJwOItpydiiE3qAYgAEIOMXCadCW0n7jJEFcXiVKTSCqbfnsrK0AX/52JyQ7Bely3928/h3w9IVL
kdLxS976OLXsk6GzijQLTuEHQoxARBF6lu0Fiy/jRrGoCVJV+TiVn7mNeSsrc02l+cqR1ViuQx6g
2/Yy57TBrl+EPB/8qBuyvwcc3vG2zFH+Y06c8XBsxCnUDMmmK6xSQGX7X2qGzBrH5P0p0pg24VVS
oAgVlgZcqr4ecfwBDsx+ENh/g1JwvdpsB+tsoNP+KFjND7vQfIcTQWbijbTUEYRk+t6lwVMjHJEB
+BtXuGFDZJUl+ZXONZ9Gzzs5z90rBBsUYny7MzdgRF9Et9IXE8Qgc6p5cCE2vBNkqjA6oXnZrFMu
mVe+gks6N3kwXxpznSc9h+bSncApj1+DiuFTa+h8qt07q20y9z38EK/h8pQevF9yG8vAvXiEhf90
yNZMsnHzOZF8UFGbswQ1FTE6POmLurwGVL8U8JBR27NuR22GTI475HmYOmLF1eFcP3X6MP2aRZbu
sr0Vj3L5XjBK7CjZJe7ob33S8NGgnxb7VMiaI17y6Wiv8pMassRCxYpQZ14/e80JUs3o5NmPS6zC
upik+biZ0G9xdOApxi+3XIoZ0sQ6zGo8tgeBAcyVLCvajxtFBzz0pyDnyTG1aNilQ//W5eINC6LK
5zdhoz02UzbuwBMimH7fbIYxgv6D7/wxGScM2TqK5C0KqOZuCwiFKoBZVWSQCJrnrAMAtS5ImBPn
ZZl+Kj6rzv6zE/lrbfgisVSSbviWWKX85pYye3wKf5mIl4VAlsZ2Jz+pyeegHZcLKvZSN37jaJNg
Fa5R1gxPB5k7CEf2lV1JQSjDV9o1td6RMnCEJ/2WH0i9YXnpdacBDtGH48+kWVk2gKdHexa9OGUC
KCBM8NyQnS8LCqKsPoJfEuulXgE/bYvX5VH70VyJb6Jp+xGY3dtUjemEIQgP5+bJ1N9H7i6yULAK
9pbofr2KghvVvifsr6Gt10spDfIUmuaF0aGIZ45KKLCcDZgSdxw6zR/pZRpAmDg2Qhmym+/SuXjx
FagD97v8zCYdiPmL9uJ6AjmWUZA1Qj2IzihbCLb6T9lDdSXa1lxQqGwp6aGRCxWGI7An1dkUkAea
aXdUN8seJDk59ab23QDGloiViaaOK1z8x572+s4MjkK+7HbbTrZclCgCnRDTVwucP2TsRyqzetA3
OXrivKD3VErQ7LHT7w68IvdLg0yr9mlDA91B3A08C1Ao5OxATofGITfodjBt4ZTWarY10PBfavYG
MqnBZNDyHpq9wTJFCcoCsqqylGONoaENPuqh+tI1QiZRSEbNz1M9J0rbmnZuQJO5qtgsWKS0mzbG
cvQs6i9lm2GBJyqEG4E831PcONliPSzjLuFX8qddM2Hv2dMjGZUthfpVLmbVWg2y8soK+4gpVAdu
l9EMV9M4Kz7iO5lycETn21d2oliS/MxWN9861oeU1nfEm0BKvrhdIz3lX9MeJHUmvrmM2nicpH4T
9xvfcgVKhyzsYz0hw2i7pW22X4kdbWOOMO505O0bOgmbP/EVcMsJ1rQmIRJR1hoWklsjHJDlLHrq
SEM4/dJrpkWtqf+Gf8ZaFi2Tb5Id3P7pjc98jNMRY0vwnpFmA0LO1QfzdRJ91n0BJvfIGrpESr84
qdPeWhwspR0dvNNOv+7INDq4PwQroIKvw1vk3yQwL+LC1z978yAeLHFZdzcJQ1IvJCKYQAiY/enl
/ntGHbkEgBxaY9gJZDCMxpUw9vsKdwn7Q931YEkpPNEIk1vfwjXw3OW4Dcwvqdhsfh6dakE9Vy8m
Y28Eo1V0R9qppP2segBSwtgSbp1cuYiJ8raFy6SAnoGNXOS92lF5CTZLlj5VvXULSXRXn7mjF2Q7
/lQt1YmFoP3vR2zeRpvNpLxqueo/QVGV2Dzy/XPO/pQRCaJR+fAbCaH8NC5OsYQIS1pHcZwsLmOv
XK2Gw92wDohJ8yWbwM0Ysg6aVoNQzodI6F1GtcvUSU9Pf0FcSM+rnbMGZBfy/2TTR2MznNweSCDu
Y5fv+Z34M6UxC08/JO+SolNPdytnRF5TeILeiI+97TAvgJceiXobfNH6+c9WitfpNNM10AjX2+0J
MXAiPKgHG83wuPnYd2T/XKi+aAWoEWiSyUXpOlGO4kuMh32Fa1TFcOp54+r2FScTHFvUO367u6e8
WD8T/01nxyH+sc966k2bdpFpezPl+LJBXmbvg8bGGQ5QE5O4iZdwW7mrGrFqoShgFEnTtnux6b6w
5Pw7QvwD6VGayievdR37eVPq34nUbOmFJo+M9Fg9uodD4lDVOh2vYYhxANWnCLQlIjcahCusig6o
QsUnRLlsL/f90ClhYi9CsTykK7zblZtGMpmJfk1aGm4qD6HQSwx2i4pNL1DBVqOl0Grx2l5I7YQA
o2Yz4zbZsJawgSiIj8cvQrQDhUJWdsSaYnuQXewdG3iGdkvVhx1z+VtmP8uCr8SB1VxpHLE44G26
lFomUE8qY3MdNI5qD2alY6FgfuyE8ailHsTqz9by+vdBte56XR4/LLTR88j8M+kyKFACKvqq/9AY
CuPMTenTKLO+NkybUurR1CTx7LMJfP70RCXaO8YXV4KjQHsNxfJJLdjbYLupEvTt+weVDY8xSxO2
Q37jz7ATGAmMcNRVide9ZOk+g8g6mX2Go5UABlavs+5bTZLhRjcAmeBYbrXG/GyjTeW6L3WHUoXB
bKnSORibi2Kkmh1yF0T3kZzG+W4FHHwaMyvVHu8jBxZ6oNZK5RI2dneixbyE7TReTV4kkAz/c0ku
uCha+8OMn+XgQW6BefzG0Bgr37r7BUCe+0TOISVzA4Y0LJOQHqSIXSqC23PnPKia5JkuTYWEqk9S
wvRO3QNwh3pU3FmD96IcOF/oWcEKgoPDKDR11qaR0H3wskjaGQIl72UdLw8/74FAoe5DxtbFsAxq
soBlJ1w2l4HFB3jkiR9NqLVqK/ez0dB2AM/MHNnwae0PkC9aq+pqYrMDxPsR+QOwNaKd4c3HIgkM
3DceJTnaIGGTNGYi7UhfqnPdWBExv/2vd/1+hSeAl7LPsAPJloizflrXIjhfYxtDVsclTV7FzyB+
peKwAMIcFGsWr5Tb66p4APr5MNbDa74ZdfB89p5uGPdijij4F82GJQRU64EP4Xjj2XhesFR1qLn+
C0nWG7T9c+mQ7nolHJwEM4PCUHZM2h+0E3KRUeCZg9+BD2bAuAsn6wHarRRHRMxMOl12mJilI0hL
jLyMpKx8/ieb/Np1iOTLVs7v1Ct9BMr2Wb6A1tTtJu2OgxDvR0kO5Jiy52SXvSfnhYr6Eb3Nl4wu
kadaraK4LC0zYSFOW++iR+afMCIPMct0lfQg2B2TFoTg/7a9RQEVRfPBBsx+q9tgtNss8TvfbUsc
ulzfK0MxHsd19NgXyj0dWjfsenq2m9vT+7rcarKbMFbTR1aICvcu4Ruaua3NmTce6o8BItbjvVP8
Lbj1KCi3ClGa2IscPPmqw7jlef/J5KY3JgxC1eoJ/BEO2y1LgKD3XYI1tstfLSXhbLuqqiaqd25f
BedUeqa1TMUmcTeFM6+rAGOisF/NUt+lBauq5FbiJjEyVQUKc0YEUs9x+0RCefkQDwBtKgvK9fEA
VgjX4+5K1+uIQCPRjvndjatwQg9rgEQBzmgWZ62U9vReOK1e9R0q9yXuvIic7dg7dV3D6fvfFdqV
yK8N/CjbgXmzAaCu4t6PuLY6L3V/ZvZ2bfxCVke0OSmVqJudtVXRZ684QprYBkvszfz4xB6gB9io
eJ9bRNP0tLO/lEplQzm+9wIR7cb3s6C3UaQ3SiUN6Nf6Ng4Tm18wBA3Ee1u1Cl7KVGKqueo53u2U
ZTrlWw5Ppll27l1Dvhs4NpU8XjmvnBeem+mzfgnMqj9GPm+MMrJiwAsXbp4MLSWLRedWb5xvwINJ
gUsHgX6KGUmVWI/D7qFkgidipk+dy9In5qfllHbIuJ7qgTg0eEe2wkP2pIBu0r/qppd6D9VoeuVS
s/KWkaevwMYjEqKudjYcSrIBd1AooAjg7PDd1jK8pev+HClyxtSyGdQRD0CyLCCGZnKU0ov5h0hI
tYcjB1RIlJ9r7YLnfGF/r12BqmBFrizszzi71gZ4O+r1RpMAk7d/9sAZfLHoMQ8Qz53qazr8qYzW
5dhCRc8+x2ZbbIIVkSfL1Xq/g0UYfzVnTrfLkmbyuRa4VLJmhmT75ZUfKaYtpJLSDek+l2tQlc2j
3lMofd0cH+OLzIdhp9yhQ8biLpAO1N42fhwpPXDPpVMXS1wdH7oNw2ICY/Cce2UrqDYn6U6KUs+Q
vlEkvsRfE7uyBJjuuJQs5uvhBRcoQUDedrQclNyfQ9f3NS9nDnI+kxPI528IWW1AbvmiI1JplGp9
GEfDeEwUPDphXBi2tFkAuIsmfBhQ42eAT0KB0HzG90SORS+cI64qc+y/B0OP2K6isfN78If2lCFg
ESYKvKzv6lGEdL0MspLIIY39fXa92/8Vx/5MwtHWLk8LMCVfqJstYs1QZc0BbzmlYeZ5twfALp92
w4ZdwQjMmPRREENkGK8L2vYQ93a06xS79w0f1ifErlGDJJs2X6DlCXM2l7xPJv1tqCTWow6LlPco
e5KHpeXphE7T+mcJvJbY2GN2czsg4KlNnbrsWP9N0ke6dOPd13tktL6akbPbZo3hI6zGg4BYEXLq
G0PiYlKKBOmB3dFxYIdU6RiAouIzOT3osswVzCmicyBX78BEhyOBC1L9HmbjNbdP5sADWcDycbAi
36jbm7TkMbkTP1+qQNZKdBWsodABOrFr0jbSebOGGEwckr86bpGAvSN2VYjfI+PaVxbTjLRAP3NA
FeVQHxoCgAvTzK3Cw0fUJy+WPKazXerwSugtSjWqvN2OsWzm0UcwQXTUb41jFSGnDRiqOQIaNNlz
DHdT1kry8LRm0dvNpLibCM5NC8IQQ8kRS0BkvB1QIibgFXOaPOyZSy1v3fWEYGWP7VqCfaZUExcP
4bYmgySjieYMXun+TtPEmoEobiu+hlmJmWDXyE36WP1LXPPzAQXk5SXULhvDXrGw7vT6mfrCUDGy
kaQsaXHJ4HkKW7dy40kGkDv7AW+2rgfbJuPYs/kYBkJVd+MC3iiWthi8KzZOhffF4qb8IBNH1Hxj
s+dAIJKecaS4PWoHhww5xMiLWBumSWMwRkyhzD3LqYW9+QXlXR3PUjwH/4sUejjel/TpRqEbS/b3
PXwUlz+46UjF4Y3A7dVRfuBCxTJfxfCL+byRBKRXWfdBgswklKqHOxz3ArB87+Qn6r0/p7KA/el0
7uXlbWSJcLwx5a6Ij4yP7sylUR/71c+C0Nf8uYTZNSdM4vVsi5+zSODyKjtRpk0CwVW9XKcw5Xuo
gzXso5UBzZ1CQLNdYFi5evBu8EIkdxeAGobPGLerz5qV8vScLoOMDyAIQFRVtAiL3Q8FmzI3Cmxm
GVYs1ly/2QpRbA82TUeD6KOIKtY7rpnwjvwkHQRrq5EHcv08cGZVl+Vy3C0KDpluEWA2EvPQkit7
RLy1u+5k4ya1NEB9oPvcQH5dGGFfBv58h/2fz0YOO7sNt/8sGpoTmOYTdcIP5U3CIPmKl2yHE7W7
cGIFUWtanF1+G/FEEV9KNCsy5T66ke5/PFqWmix23Hr4sU6xp905X1U/qf8IhhscGw1FsjMwtPZa
Rz5PkixQwhCSlkn8XO5XPlPag+CtDo8Mps77k/5vDqdBFQNgltvv1rAOMPg/qVdnmaNcDuPRejmO
AqQ0kKgGrMiJCKBQpUSoVkSLQLgmtH+De6ZUeRoPFtwO3/Ri6ELuI/ZYYgaXo6jmCLexu3oKqoXF
w7g+9O+jUlCxMArthriB9VtJKUiH8/lSSXJLgZ2DoocMYH+NAhPkMxvGocqnh2htNJWuEXe7ZiFL
bfsIKig9cUFeGmd+KyRhD3bvP11S4lkVzaDJowoz6nthYeAeCytQ+maM4kOhsHkR2fcIAK7blNV+
2ZrFl8PivyJqvGYDwh2PVnj6ofrS2AWRUCX2BjbIJhMLTNbi6OzJIYmYMmJgr1FwezstTftGmg5r
5DHgkaTePYW/TFFwsOEZUgsTICIuZYKdMwLrPrlBzCFcT8EsUbwjo2KrRw8RNaKlzKzepYlu5/59
rhM+LhVh9sZ9ZMGqHEwKwp24RebeqYPW7AlJt789EdUwOs4A/LHBfr0kF6DDyg95A4dbloUMS/UJ
BZy/Z/QU3kYYQYiqmYCHJgkR8jy6Jwq/V7dUge2H1gmtlJJ5IfaPhsjGiOIcwMD1CXIy/NH2uEtu
aOxl3ozsPFjKUEQfpKwqNO7cwnXW5BKeapwLojxO1RHS0cMqA9TvERh1U/UfcNZ0WBoZZj8+PnQg
QtbPe3ZSbN1ft4qSxOlvHLQjJEyYk4UhoaETq+nlArj+9JRbcdyE8gzhNgQI/phc+5zZYhZk+kws
KdG7dxi/gJxPeUMlZCz9J8omFCgTLnGqP16g2EnXIEPUf3TwxGOej7U5oUyXBNBPTH5YpN3TJhA5
FqLk0KviluKeBsxcof4XrYaBryRE6xgh0nrb+niVcccAfgeYOtIQnDpin7rKeBxO7FAwDpEqjAVR
BqVbwTi2v77hqxvs48YSy5s446DKiVq5d2hwOASStlsCdJII0I5THaYfNZ5bVGzM0tFQTZFrW3Pc
1FDzZKuzb0YwtthpKZ8GjGDkau0AfwEEKbKHK/rwdLd+L0TE6/pdxFDf7p6AYsL7e1tvygq8Pkxk
8IicWmyLscRMotxfR+4ubVEs6ssN+2KbCF0YyW0iUaLhb4b0yx85PBRXCzqXQ8TU+t0Q9fmxUrOh
Oif6F2WYb0nQWo10oi4RKlr3SLHIzOKXat4GSuNXW8h2osIt8oXruzfxYtYHYKGW+uiZ1DOzNRfZ
GrOEjeYs+rNHGcjUtZLR+7Pc6h6UwZRI0kUA+zOL7L3xjMHbmTnLAhA5KI5HtjVSoA3D2czbtNO1
sS8ItoCUhNwZVe37qzJNny3XWpv2sOEHdWr9whUBU7NxsHPz73jVvHGaZIw2/MuaTmGPmvJAPkUr
VUJrhGfrHL2V5Iz6JjIp+MmP7fzwY4TwtEjz/MI4XENvf0j/dJ7ETj/4VAZbR/CqeDyPb/QMdThe
skpos8vLjOaW51k4q16EPBQLVtLthlfO3RNKXP99TrcBnngba6zDE+lINoWaJNFsGA1JgXN13DIU
55E3SYpYM1ycUHADCx3mMW054eo7KjbnaSF7x0UzQfiygJCxTFz3VP5Fc2hYrpUqt9w/LR9CMYOl
cFR7U40gGND7drhFVI8PiUpnF5r4mgcOif6Nf44sZWpT6eGdL/2Cmo1a6aYPe9rDlXUzmgeiftzM
BiFxgXziX+GH4AthCwjoIurG/ini5IxOf4FL6JM1762fnAD01zBORQm8xBY+NMYac3yOkF4VCjQ9
3r6CdqwYmRmBYcH1Joyi/ZC3pLjlX/4zt1m/cDTeDNexMGOxqEjPoXOAWUcGA1O8oN2LTEggRWal
jt9jkfZupFDEQU7duwbSlo1B/k0YIXK/106WSR3yR3/qkJdbKAExcMNyAkkQ9WmxOLPH/l2hX2YU
ZZID54TuWhGzRZQ3iFwo/BU6OIBhOMcDQQNyEc3BZIRNx6isDLQ63C9i/edXaIZhUq3FEftslmzj
VnByh8y+B/KYW63hIP+NjnclHDYtkEaetAdqKsPj7RsVsocZgTSz9mEjhxXutE0gvBbWzHRV/E5X
TAymV+ux/S35Kl9N/y3coJKXLvu0UvyBu6s9uo/FePanJ+fUGO9Ufv3OMfyvrK6dU0U9/m7zkYMO
6d1qtxIDV1DCCIDKCFObyoZEzkIe/Ie/5r312xh0ozoBWC/NAookTIVPdvf+W9s4n5Nb+sY+4RYi
nvdZDEBhY4wN4AyhJ+iouDkTOj6TXo0F7y3URxsOYGMxjC0EAOgavsn0nnWm5oGL4+2NeQ4R8dX7
/sXck0jFTrYkwSWXh4a3pNBrZqA49QWq2Z21EW/w56FXAhYIVclYtn7R1INn0AM0JertS/qLLj4o
Rc0JWtch6ybEx0G/MsmCXeKl+yzf325lIvLhck7c4KRIzei4uQ+NGzq9ryMvQU02KwkIB/MlaFil
qHvVBYTDi5F6i3u+VMjvIDPj69BDfX5xwkJTBbpAeTCTpqTaMq64fap+aM4tCk//ryypVzR/i4Xu
wJhrsZfuBlNMXrnTQvUVo+Z450c2fDPPFxF+y2OYMX1G9cTowqVAFmnX+C0IDsgLGKbRlftDVudM
1R8tNtfUtrPd552Mu6v1BEkIllLU7lsjqqFJrlnn29sO+ISTCaMdIqj1HsXaN/oiOJ+xkYdIGeAz
ObHbb/+u+d5CeEn9sNEZhBe7YKj0oJ15CG0VwOEZ2EDPmayN5Zj1qypNYdSWVVbdZ8/JpKOSNifn
5ko2sTYRfTcsWskU87kyJBlQKpK3yZ1G5YtOtjKuk1rGDPFjmj5o6RbwOds4LbySrF7HoKDMgran
h3qYRt3pMcI0Va90uqBNI9ysSXB1LjasvBZbF6w0QHtFLb26NMEBOP8023ipvt9mhj6wRBKuwPSS
AcXKFhNcsnXRonFlc32Vn/w2fEvlmVe5TQ7UX0b1hVaTld1Shcz7M8bhnJEiBJWauyMUxa7wMSX8
hv913qmEZyFsN2BoACwAQK0oXGCne0y/xo8u6AmMItXxGcyW6OpFdX+NKqLVKKxi+RoHjjsgX6gj
XPKqRNJWEBNLUkSNJtnNmzDTvToWFIhyb0f65bSKznc06qJnu+BXnO2Uue7kxJpRSIHu+jWEL9uj
tyDTkZ+SLDaEvAMQ8xk7nOPbUsnC0dah7tmQ8/QmWCqudjvlKudbIigfaGFZ8FgISM5hx6+pHq6W
G30yBh/oE18kPhs2b2zuKB+czuqw7pWKJ+91Uxnjb5MxkHeCaNgMBix89D7fZM52Ttpqkvq14mKy
0hC9/N3RPubcafmJbGZE2Z2D99QrkTQ9+K02/uH7WfZkQFZTf7AF498pPsBt69SmJ/Zv54PhS3zx
Y7ttwqp+WhpsMbtFmpkKlJfrP+iZDfMVukT0CKLNME23l3g+ZbU/c/x5OeavA+v5QyBCK2VRb/IN
DWFEXJuzQUEs8E/FKY4Maiikn1URapw23/9y4gZXZcgte4+jOqZx8DFumAMQ0ItyZn/iHlJlTFui
+4GrMJgNr+C/4YbcbFoin8gxBMf409reRV90f+ukuB3kZIllFw6l4v9qPIA6HUm6Ktq05zDRm0HF
vafxs122kb4ghkfymdkYeTjTUg6HQ09CFoGARm+FaY4OE2bmaUwg7HSdu01Fj8IyEmtCake9tfNC
+Jf2I5KCYg/GSvAfISpycPi7E4CTq7JetLeS0gkPK7E6Uaz0eTWQMDpw0mlQ7CYP1xZY+ekTt/Ss
PihykJYRamtz+/KNZ6iX1me4mlPxi+OEHSq6uz8pTAB5FscUVuVyOJRaxXUsnSudg3APpYoWoXJo
uosUUs6lci7GTy7NWu3hXtXCzif5mhNu36yMUS8PJlyzIAHOjXwar/3ooEBz+fcMnWVa+jR9PoU2
8wUznEslQChdWBFASeWp4EkYScpto/IAmmZI18wRDHKDQB98VE277QPQoHohW6bd0oSVIfm6oEdL
LhfB4nrEcPLAb16gXNljwe+4RtRaDLogX3wkjwJnbbp0Ipnddub0x2L2MMh0TbNcpTuAVgMg/c8B
Sm5RUmAiJBdP/hYuWkZDb0gntWdCeFRb7UciQbYmS4hJnZ30Ap7OVfJ9nGQ/RdX5D+ZQh7lP2kge
3Ev+JpLigTQ/L7XmXkEIxnmkwe3xUiYpDsPSQyec1T5uDTQwGIEexcV241FXcNxDNtVzlrR8BHDZ
rGeBv4miQFsTqKG7VEoFAd0BrQsiP74NRz4HkMcFiLImKLlxsWHCPbymOJs2p+7kgX9tqHjVuVGJ
u/gohpwAsbLRBZovQNIlnrcK59LAPFpJMu/toMDNchpWv1URfDLlzOVLjgbCQZBhpVxX4U0BJ9J4
3Xvt3EUW92n1fWh/c03v2VoRwGDq57B3zQ8LYmgtxfGTFLjPf5/NM6Fn1vCvfaWY/NP0LKrUv4DJ
JuLvCFCvK3EYRdCCVR2tt2VAblaAI874NZ8muBZEvWHFKev6DXmMDNFHoYpdraAZdhW1c3hyfPpD
WJvTTMuTmQfSgpShTJ9iIHRWI0DOe+GgYrT0C+6pDFKwn0X8uNlYHFthmCXaUn3d92R40qhM7xkJ
JU0X1c6QVH3ykq+BtjaVOOz4mQLhra9tdp9uZRr9QnPPU8HkWLoyALT+2RMc6h4nT4buCc/h/sUC
vtP3aFVM4TlJjBCjK/WvKBQuj+N1QKvPBLNqvzi0e1fHdRFJws6SxM9uVy6MOzA2IL3rKKxZb8xj
EmsvO+m0ZPh8+4WuMrdTgjUmFhjQzfZtqNSmEqqCVJ48Uy+q67+pCA95zlkK743/TbulURqlacWA
VvZqT1SXmTzUir7WeMy0cuTz7XXmEI0Tq4+Gjgdx1z/jQqmqG2byvFGUJM8277y96lWihX22OA9a
/E1YRPjsR0qL/AU3Y/DTqqp8zuQ1aJh9PP9gqXhysKXyIrsWTc/RkhoGPhGfJ8TBTh84lrl1Rx9S
zAUm6HFanOqgbV9RjfQNKGjlGhzpGw/7NHswzmURye3Pk4kwqHJNSHj1C1FumudveKVtmeZnkayv
8vk4UTUHyvR66Bb6YQ4Z7J1OpVeUox9CN6R+X9MG4hJB8fYgXAnPan9vTGJVV+rqGMdLBWut5uPj
UgsP2dzu9hXdwQ8Q0cOoC8uUuvnaPGXM1WE7uYSg9lvhAgmreeMcUdO0n4Cgjyo6dE/4BLbVBNAe
CXTIuX4TpWO3tS8lpy81jCYn5wz00Yck2e9mIrZpAC46KPXHS9kVmSWj/cdJY4gw4L0CGqCbrMEY
aO8jZlurJs9Kr5lSIDKFB2dp+zJAELWDExNDsHxQ4yXb+BHCo5JTLsORL2k4FgtrZ1uhfXgw7mlm
HMlh28GZ/g49GxiKGbYCR3Z54u5qg1CrMTaJdvJWdN8gSEv+ODtD0iS0e/m9YggQolo04eTmbeUb
15jLNl3bxN6mRuHq1pPqsTyZ2Fr9L5zm3OsSROva38i0NqFCLtxqYmL8kiAUUmpIA9DDKIa9cUCM
+oVGJxTo2hQFPEp4bRg2BG3EXfkGV0zsHzvkpBvwIMz2Oe+d9emok7RaDzM+ik7Qqh5TTMlU5wNi
SA3vOyUNQ7wRKVJCBCYSDF1FNANn+9fRXREkhJjGCx4ay9SlCKtmECt4KrCuS7Ay5pjXKme0aWJv
oBO1GyI18xLSXZ8f1+0ZsjnFEU/kTqIv9AVZJ2/KEJlQXQaNzH7I0Lra3z8nc4RSMcTQlM7TQSm9
PsHn/6Lpe1+IggQyQG3THKrzA2lRWmqF2E7sNuJGJ/Ot81wAQY3cEdTR9W83nEjY7wajFMsXMYl/
oBOUcxV10RNWSJcFO2RH72SL71Vc5eIZHJvrovAdBOuiBVaPIQo4vgnnaKVmz7gDn1y8mlSCB3u7
uVl/POLmX4zeIHqx0+9p7ftW5ikjQOXEHHKx+mK6cpVdhw8wwD8vph35PAeWyv4L4ildJVZKKWzh
bQT2D9urRanaYBEuh7eH81hvpzUguWLmnODhkIaQzJY6Go3HIpTGDZ3nXTMHClscmfycNpKxlOqX
6Nu+BDrPrKuOnrslUil7eSwt1t67C5vdEL0xl9teq/dibx3JpDyMiTveQWsuLz5sLN9qLZJ48tEn
Jjsk01dbLNalyKjo+9FMXzdvuYgn4cKM5G2XK9Mr8QytJZYOlU1Wi4vaQvUYSl258AWVKweUZsc4
bdUEMPQyvGk3rgE5WGXtA7F7UdXEw2R2QeGeYZ7igmpInxGSIdE4bogoupQoeipdDtvx7VTCWk9B
n7nxKA0yW5iHS0EnLmyJab6e+bZY9EfuSAl17nObvDBnuY5U5r8oqOMS93lsE1FVOQZJhllEd/Yu
7MB2hlEi8rka6ZRYaYawb4OZiMACR5qk+ngg6qG9+yv74r9cL4ouWMI0ZndnbbFvJcJTaKZzsUV/
1aT/D1BFxdnt6L2WBWzJnezDVW1G3/Eua1w8GibHWyn+W71bhuNk3bZRiMpet8V4tEG7aQzkEKR6
1CBl3/4llrdNnHxfQpcRYF87MSLmUQZr98/286JXCmiM8QyFWs8d/FxfVBJpUVTb2vvwTI3PAa2v
AgKPvKuEoaAhps+KGbvkU6B3L31p/6n27NQFgB9LDsb6TXYTpznWvMqvxf4634gQAslSnUYJJEL5
7ILdw5b0JxZfpHuxkdCmFj5FWRUuocENwxVIHXdR0mKpEpvtKAsXYB8v873UwWgp/Ida+WRI1aHc
/nzcsZYu/09uWHfQy8GNXzsn1WmzO5iD0JN09pZsxSl3tpa3WFs3wVKm/rxr6TzFSmeYRJ7c2Gyy
E4gEbN/malCcnoV6GAbGGoeAfzf6ct1fiIggF13J7rYRJMJCPavA/KVZoD9ofEob1lN54XzLTNjL
rPUfTzoqTOmmo+KzCDfwl3eaDnl7shPd8UbYmlgEIXcPY65YnNtmqhxys3zmUg4DUARGLpCM1d6/
j2JEol/Co1sLOx9wKWaa5i6a+FNUkiVmxZ3CUbhj8dZiqnsmTStpbPCJVUV3NriaFIv/aAVfYGTY
3d7AQlfsE523SsoX23lWEcVzbpUO2d6BmvQhAO4GkVQ1mzZBij6f17MmqdyP5qW6S8qsE35TKrul
KpqzM0gcq/wuBO21h3ER76S49Fn5pJF65muHoUbyeg6HOluAxpOqHQ6WpVslWXkK1oOLhLSg1wnw
1aI1wsz9739xdAIGbcUOFNkUkJKbZewQxYV2pjmfQy0Q6GKAb5w5eOhQxZjFFqoYgOx8XtpUAy5t
VKoM0rFXa4jSpJ7i2umdsU0pV8e0QeXWdc+4Q7PiWkECds/vaJTMTTBoy4RAW9oDyXAU5/kEWdlb
MSaofNLg3HK5FnSaK7hurb1L5RcB0VBAEDUzWIEoaIhjEzF07q+Wf8Vpj5L/VPLVF5TVzPlriVGi
9EIp5aZvlshOmtb205n96L6rfatMM05NRGJRmXYkcSEyKhMDn1NYPk4Z1UUKDoKiwiPbIq5j/D8/
2qeTyrhiVwp8AXbFcYNMsqK7Zcv43HF6LM61seLFxAtWxvSZ/ijk0bDSq0Rye3zja0weKSQUXVBC
e5UwIiikS+pTNBp+Sc/UckmHewdWD/bBe30Tc2w2/7iE4wn1C4czHYhXozRrSRKvBDZtD05W6V07
vbdU3qWC0nDFuwUJzlwLuhq+u2BCkef7VW5+4Or9WIyEUSoT9vaiA0VVAqD1SZnmAyQpyYofaRpU
7Lj06rCmADUyo0OUORUCGIQOsiWoM0WQRee0/MHbz82r3K4eERWJS4Cw7CxudN0UYv9xiVI95JL+
B1btflIBObDtN8cmQmN+VIYROgjX5vZuSVuLQJ3OXLhPF61xilTl54GPfjSn98SzOkFvGjTphq4b
1/QKUrfjmpDjXo+LzZSUHK/O3iQBFtM17laVSeWQnwVok3Kx7SchZt0g4Il7lLRohZuUpoITsJ5l
dbDrfUZ9NLeF7doYiiwShLfUWtts2GBHmvt4FzBrlFO7GgdiaLvQKQLuui+Rk6XpA3Bz2EuLADHA
YTXDFGgUpPCqPCB9f/DK8cgmD28HKfzTDQ20sJGjNGuEfdap+20l4pUBbajzdiLXE7Wi38tsuqbQ
8fQJsRCrz0sk7hBbEBvyWvFBufWjGhxxAk44cBEOXJx0ZNu2n5TmyghobAqX5lVNMywD54Q7boNX
SGj6vdt170+WDbh4eoUTwCdNc6CfN1E+JHFlrrayuQFsrzienSqfHUq4fH4yTWacRqZX/XFVKHI0
nuoPapFSe8VoQujhahYHXWaP/ZnYr43wU+nL4bJcAGdKQv/ktHD0Blh5EXG3AiANBDNYsD8xeWZh
vX+NXcsC77AIc1++Hu+kLMtgsIGrsJJjoeUAAKj3WvJG4gIm/iGzN0aYX6JU3XaBxMBy9ftnenor
CTETzn0uMGTSkN0vTk9IqqbpE+zHcNP1dKFcM1BPrt9KG7HLNs8EcOBq8EYglgWDQHa38YI9UQGR
rs13QITkZyNXKekgjWsA0aL6s9sjXPZS2TfXGJgzPfdYfIMd8p4x5crpf+3oy5X3/OyB/xJ+87U8
ImdU14Hmo6Yet0L6Lr1s3yNmhU10i/TYt7TkIBX59acmNvct18pFoM/6A2iJ4ZFdrHQdfm5cegxt
FYpEOVwg+8gWiw1e7i5Cg1jm/UyvQo5Ra3qCX6Y3ml2f1GfrcPNndLCuxbwlTLwWa/QOf72Xx9o5
ToAl+NkwSAdzAT8kWl81DagDFFigOgVrAQa6fohvu8B3TcjzZ5cJtLnj5L/yRSx/4aPvUK97elrf
rzGW4YYhONAFyffiMX83Pbp6KYiF/qQc4eRnUuv/WCkoMLAbS+YxciBJz04ZEutaJvChsQHpCSfY
Cceub5pNhvVE5u35vd5tVVhbF72bLwumtaYamcz0t+E8Yczch9OiaESQpkhSiO5rn41g2uwb6ahp
lXmemzPGNbFyYzncHNhuK0gCfIjfUf7delED8fWMVPxU2mhN+A8YHUq4RvciPDy4hdVl+Wex83Sq
9qU/QPn5WPLS6KRuYRDemtuPobHcfID8L5H+cHc6EePev0TH3RtGLWQ8kVdQX+eoMsUERZvf3ndx
7JxblT/pMsB72jgCOSLH5igaW/SxxNCm0oXHiZJoWiXgvU9fgHH/ALvsfhdTPFpyKY0nuLVmQkpy
7PH7fhjp2OdQFDZDNOTUlFWAk7WnpohHgzeaBq/N9sltFHUQiHcLbsvb5B7w8kHqUlAlzb8zO6aM
ZpPy+McxanCK3JEq/Nc08Mcx9bv5k2cmO127uAh6BJG15eo5F2GwiOa5YhiC3i3do+uj8FaL134i
rMGMRbKRcqVHIyFVKccDQe9f7E81nZ0lIuBa75ZqPUA8GZl47yzAYBMOluUV00hIyD1fDY4uI8zS
Bi4ee8iGq2JXJMjNj20rFFsMPlDxWiOtCH/NtWqBz0k6Gi8Gb9U8OVlziyqwZISg1cuIrvMf0Otw
4lO3RXgSX8sMaUxojONmV1p2/ITZhXBlAhNCYr5kAjy1nTd3J6kNEeUYM9Koy7L1gGOTcH5r9Mfc
/XVP4zGw3SnANW/mBsZ5AOEseDocUHEhfF/f8G05dEbGojrXbzUkP0RfmoDc0tL6oTJhViRZN5Ek
EpshrVZrRfovjW7WEK9VO6SrTECOhAeq7UEMMD5/cp2MMXfAC2etz5cLzYeyrdhG2tvQjHXi6XTV
CL+fhL2Srk7qs4XHZZsRWeQOQsoVc5Vy+9psteYbSCCi7LPjjsj+2LTJf47/WAlv0HR8rLrHNpiT
MFA6N+c79mJftGBpN6GbUHyMldiVF0iUgRiLOxFPBS0g/M/HNw6VnzziGd6rxAkHmyQWFhX+clgX
inap+AgitNFrE1+SIjYGnJjzcE0p4cTnQH/9pqx9kVTMh1QiUrBrPNyt/yh1stNq2UDGUKvtj26X
o5P36/KS1HyX+xNuI0ABmIloLyp9a4bnGbegZh4OnLXdlv+Nny0o0p9E41M6cT6UBrI89XzIiGLQ
iIs8P40KX01WHIMMLOMY2xrhTX14G9KKELggocNFjF6EzecHxfttAI4k6DVxqjDTzGUQKW8/gO5v
qYY5kLBCyayuqb4uJfi3LGNF9sWmxfytxLsTIGU86bFUfZtC7i/g2QM3QyTNDP2Co7oCq2Vpy5/Z
jMIrj+LgrBIE24Mgf9LPGRjgPLH4TVqlXjKQGIQjJWijI27KLbuMQ+oC6vTTditMrWmr9m7p6Gck
zcfzKQULvR3vJGvl89BVes2evFemPygPEgYy2elmTN5TdcTzScj2Ts+88imYs0cwaFLrHDvJ1Uc/
fqfmdj1E/zkvkV1QbMvZu1K0hz61MvWkk7ad49jWlNMr8fQJ8WQWx5h+Tn5bQqRLuftlFZ/SlZpu
iUPapapRqUkUxPQPKewGz7tSCB+uDJHJ3wndS3rxEFqQK6pueaGoVbXMkowbjdvUnXWJgYZ7+B+r
g9SGtiitn2aOCa2uDZUK1pG/674Ft+QyrgBozb2eQOz4HZRc7qmZSJ6KSU0HijMpUD9SLNnpXUhY
8zCmv/qqEql6Pg9M/tWwJw/kpkQMwxwipuyiKI7RXoL0qMSrtMCx5XQDflhZ68cQhxn1E5d24xgZ
cTCJa/SUM7zYv2cMDy0VXhdpiZPZFqfKqd7naw/pDiHj08pZMVZaVHySofeAP4T3utyJTCUTjvEx
HU0Ta8kpjsAvJUbtF8EWAf4Nj008tG64Y292/wID5QAexCCT0/tEIHdK3Hxk7bznMj7JyxYhAI9P
Fj8PblRO1EU12bkXtcqNBUySAb3olgJ6jg7infsDi077RuwQhcapD859JDHgJ+dJipuqyIX3+eX7
1Mh5BKiOakJCwrg3blbmgcL9OmFbCczZBge6Wn19FB1svrYh2aoJCL4jWxM+AtsEEReSHhlpMyo+
7dVUaGeDCxV7lkvAwekHjeAhGi1i1bpMniSY51L2WkVAcpp4TyRJ49mCbVj3wfZ65QRQ4/vQwgr+
hs04lBocnuamxADGjqfWEnVxN0a+E13qOSnt9pBF0acXgilI/YwGy7PSrKMnX8SqgxyjesIPB8oZ
s1L22S+7a5ERUhonz12uQxLE+sMHjJWb9DjFwRjrAg5AQOgsuIHAlKF7SOD4qnWx4iGmLo8OWWqK
3MhcBe2SgRsJDrenhxHIRk43X9KNO/gXO7o8FEGlVfYadUowfPEhKd25qxLu1q7dnlgtN62IXz6G
a4wB/olCCuVmjQPJcSejdAZM5S/fHU8HrFiEUPGjxSqhtwgpyS4LV4/TB8R1hPlIegRfq84RknSa
6plpH/oJVImeC3ORrL4BV9SvD/FV9VusdjsiX9hMmhpFltI9H2eVGLxV7HngdbTC5/eqJA1uLwox
p36UVXxVkuI1E0cQWEXn/du82yH8zEyvhuUCjm6EKK/em9HcuyJXHdU2vWl1YeRlXMiSHhgBE3UD
in8E6dmgUSBa6OV+aM00/x8Dv+HLzjSAbeqX2lfvlzWXjEp07w7A/RtEmnDBmFtQFlboDpGHoJE8
dGfhfNSFkapb7LS7Sn4cc7fyTsc9LyS7muNPYXHJhXncea3rskLzD0yzoonk7ePZ4Biv/SEgFtLI
3/rw4nvGy5mXDe8PUthq99NhMxjhfwEMDnHVKi4tmOAQ7R+GfCEwyLWXWvIF7TM29SoYqpyIxA4M
TG1uST+B9cRpIY8QuJriytwPIzPTShCY/ovvMflwiDs6xddYvcUI753EEjckvEPRGB57ivap/vP3
2lMqeOJDjc39eOyMLusoN0fVmgXotZVD/H45sWJ6s7c9t5eNsDuu5Bx1glnwaHjc0gz7Xj1l47/K
DrXbDQrtU0KKbNHDPrUmhadWqqtwctTemvgKYMJ4GCZ8xJLcd34Huu1wYn+S2YoQShcrJvSaT+J7
/EHyEFvDhXyWsTXqjkvMiJDF2Yhh5+i0IlF1MiUF8DOfupyt7l1Q+wXfprkhHEiKmEELtPDyYNY3
Xqd+xvjeOMOCgSO9vg+k4zMCYc8ct9QlVpW7hGio/fB/0zwR8GSK942JzkGRBvOqEg0kkee2MrW9
vOtP/WucC9PF6NSLvIQFh8gD4UHejYOhKp+qytjmNZeumiDqYa+Vn+7t2xXqBkqSbOt7tOTHtXM0
61gKNzv7uW0/3L+jix8/Ew3rBWZiu+B3rhZWwObGxbzIZZInl9a62fO8ymyFqnHdOM7xeQRwiG62
q7vhuMSwCmaaCTRi/mdF8HywQS4H7y6pushEulFuFCBVPzdROqf2v/xW2bHm3i0XoQ4azvYDwZjd
LeZdWuACvgKrXt/wthPlp2U+6iV6aBKQGUFkFUOQ6rTCkl5+WjMzRQkdHR9rBv0JuZ3olk0KHOkS
POHt1NOqKgfp/ZhUTEJ8WoCcLu0B3s13LGJCeKVzLH5j/4jpy6NS8Ls8j4DbEjQL3EaCR6pXl6N2
bN916iZZSD0Nm8Yr38ya6XUPMSFG2LqKseNSnhVu7612YF6RoXU60AgOeFXFod6pRVb0Ng7hvqTj
yQYQHFsTmktGULgUaye/rnOHgJZjF/ggVttMXKVu5NoPztnh7ne5jkr9pFeehjbbEfH2u4ZlnvMI
s4Pwvx/QyuXx5IgrwG2cyk9kssvMXaAHPphvzh9oufTb1f/qhilh1hTnR8KiJJ3m6ThqvXxrODI+
fshet59I4kN8+wvn5M/8Ib76pccZrgGzPUlwWLaS7sxySuaKpuugV1u+GrFn0mZtGtLbC+1lDTtd
TLhNXzufYLANsBMLA+vNmwhfaZImDn2xR3XW50NmkhGhu2IyaqaMntKlUjKm6aYbe6d0qjErfz6l
tbenGYxGvWT5apyeVfR6+q1I1pZij7o/B7Apsxnci+hdfQMp1QKpjmU24thvY4V9BoZYfpPoYzwv
y3hi3xAyW491vYkB7dk3ObPjwSS8FpKAKJze2pvXRRY9TZSq5BncjszT4/TBQ79g//fijm1QSCoT
cMONhL2XJOwegOgmlUHcWnrJG5YZcTbV87u9VXqWQVJlw1XkNKvcCa0IWtF+qj76b3TNpvqK0cSF
8IYKxYTs0Wv+bLorgbRg18GwFU2uTLsfI5gOkUbDVKlLnqkZRPNKYhr+5vViG2Q41+8xOyv3Fb34
VH0wREzXAzW62O76s4yOfv4sYJKUd32+12f4DAMmMkLWnK6La12gl6Uaho7lP9XoDmKqk5SnNfFy
ye34hIx7w7jUCmHijpSSJlubkwUVquChmRqJVCdFEiVZ2J7Dvj6lzM3UnmNFntv9rQcIrresXvW1
i1EmGn5Bau/C+SWpAnhrqehKXr5ndEfMljQynF5ZLiCR6/jzUwKYTh7Hr34JV1jmba8T5tjvlHyh
EuFZF1RX7YO3a18ep2VmQ3CrpLSf80kSQ5V3J9nt2QsiLIZUTabhhCnTAvm/nHz9DmxZS2hOM1fs
Bi4BwvgVr6GAK9VzzhVV/hVkfMUyHuCj1DuTpHez5n7qU3iYGnroxoAHUQS1HKI2KgYZYSaHCPqf
jh2gdd+EI78TKfids/B867eyTngbLrCitE0qpi1gyRlNg/82BDqV+xxR9u+oAb9LGFYI/8c6SLpU
No1nIj0i14BQkgewUEvodqSyGowIHZHGNFmvBFrUUZ0dFbzpOv5VopsrDtA1Ky6JoC/4UDtdiRXX
HjBUSUj/v1tcNqgo0iaFgG+/9B3Rfx65tMbFipArznJvGb40W4z6lPKgQJ4ERmI3fY45f+VELEGs
/CqZF+0KJYTmkQxGn4Ca06ECV/T7CVSq17X/Iwe7CW8Pg8XNPlQB/p7MN/+HhQ7pGH52TEnSkFFN
/WYxg/IINALpA0+Eu/M8RkgE5nMh19+I08Qtq06YsBAWa4WA+RXQwWaOCR+GfCeAQT7/mlZ3LSyi
WD0bxqsoOfG0EdLFqKp9Nx8ylsqN417zGEC46xMXQnGt4z4uqfEtQ6/tHI4eS5AXbyE1ZH0/QEGL
4YbFB/PxwsopbJgQVBwg+QZdOAOxoIcgkvAAAHalcuD0xMG6ccwRsoL116QD/7gb06oLvFn7YUSg
rkHnnCKiTm4ejh7KxAsr1YTwcwStW0udmWmQ1FsDMTWVybAqgq16TZJOnaLk0zDPZIRS/C4FPnPb
Z9X4avGA94bkWi2qykbC4o5yKf+9RvcfLBHSQxFtJblrRlcUxBir6JmkgYXXGRM1r/gv3sHx9C0Q
rWdS04DABvQ+zex5AmclNqOv7TZE9cbveusl7jdb7LNmqalJrS2ngz9Ub3bNZhC97cL+1izriCr8
faxXDb3nxL82L7pv5Llx7hZHCjzwUjWH8zh2yhnziG6C2iAe5tsMvsWltg7QGd1pj91OKbUsYHgx
TEmcCXXkHEAbQLtKyPPoNeYAUveM1rrHUsxjY/cw9haZUQPyNai166aWxnjMeUejD03IJAT5DK+C
JXjTW03e7Z9oJ3dKxAZhf/9vTKjdsfQs3JBlR/+R2ZPC3X6E1SD7Dz+46yi8lvAVPNZcSuOGoLks
Zry52U5oKs+HweQexEJaJYB6Ok7yJvViZQOLP0Z7STtKC6HA3fkH2lgA/E0ftSBkT974dNmizA/V
nqFNH7VVNPI32FyUeMiHL6IDcUEFxdZISZFK6I+zXKFPOxnjbu51f1Pm0gEZV/BFx+YKbeML7S4p
hnUJRCo8X/slYu3Bp8JYrflu0DJyR+BCco1xDgsI69wM//hW/DcBu1uwOD5MLCc4knJm96E73Nrk
ENxfgp2YQi1eXdhtXw4SJN9bZIoFZvFD/6nJ3q9043qQCREQr67ooiqiSdAdX15k3D1iQhjyDOiw
QQt5CgS86HTwO6ztM3g/EdM95l+Opkkl+zVK4YUVtoGIRuJWwiDZE4kBIqFdqYTHz5w5x0j3Ji4h
ikDUqriycS4xhTSIQuNwjuhrE6aq3R0oBwoLAVRTg7BgJ2HyRg7eYp3R6SBrJKgS+hg3E+4svJC9
wRlRJp1RhLjfttvYSGMm548BQVOAK2WaXSszI87bHkdVqLBqeueJC/z06/xGHgH7cuGCI2eZvman
8v8E/2VsRrRWjbvYaIaKAUg3y1ssVNzC497Jff6OKN8UIuD0ET4Ojq47QguLXOTt8LStvyuTUMSp
SNz/0Dj5fxid0U3DKyRFMTOvl7twKmWeK9zAQlVaPrYJ6vauy4XghkhElIlkVZqMv4UWtWjWBYG5
E5S8nY6Z0Q4a3mSPPpyxdWjW0DbfhAHLPniWU1FZtV2sreIiHaLbBEIt+KZtzUJVRmv0nEWJbdel
VGOH9dfCJMSIk1IghAs89VBOg5zLkx0ZfXiN8LyO8ZUTCeI8QZYlD2os8N5Qcq9w2vXMRFOxM2cq
/jZ6lLQzjFH19enbD94reisaBUxSwimNFP9MOVFvxDEYpAyJg1QDMU9BmloHJB71u7VU/FlCPReC
SaDncv57c0bXilk0KZHXGnV9t0DQGT5KBWijdvEr9ThV7WT9e9BOzGUMAP8I9ZfskVIrLSVc5jMC
xEVmOjTLVQjPDdxJJuxFdz/TeknBjUZikiWnIfeStZC1zIxV7rsg3hGAnYNGwGEXanjn99pAIE8P
VD1L6kTTDoiOGx8PA3s94aNvpPWVvXi2SaGjlfu0BZaP6UG2ZklqKqxn8vlZwDgm3qMBYHoHCv9l
1gEwxa4FcMDoXJin+Td3lJr9SsPlY2Zx23/y3oH7H+dzgMZou6ZghF9IMaNm/gFwALs7Wjcsg6LK
LP26yJQpNczCvN+8s+nZbpv5g7rpWbCnWcuYUq+Xql07Fgz2ckPzMITbgL7aTkRfxtxYPH6AxzFM
9ycRGoFqOGdMHviNW58EjqLcNptTaW54JLkKNkxHCwt9zWzvNBdwCXvqlc9Y1+GJkIssEvAGzaZS
q4HYmRmBHiB5l7IukNF2fbNESJy5buzWAmXVTbVzBBJ84p4fYxaKXaTgnQFuHxk9z/rBHpwXWi00
TZ2ZoG81b4DDzZF/HupKSb01ItxHhNHq/U24t5mNNjf9PCWtiV4TQCdah5+b9rNOlUcW/aQv8Bmq
Vc6NhE84cl/vlb2dsG/YUNuo/1Oh7OL8RTw6lkjmWCgbTkEe0alEH9RFhjt/kXHbWTIiAL2b9KqV
UhHD1HEvmvVUrjFex5RM2H2Bh3yF2qAxMTp9UHNcFrQGNjMn/QA6n/bjYjxXcib0/S3C20dNC0Z6
j5aEFlChub5uc/tDcRpdYmgVZm0AlJEYRQDprW6xMNW8FOkYOO5xcznCBMLdI9+n/js7V33TacDe
FP4K2+YzUdy0bR6SJQfT9hZKihsLuzW5QPzIITWDAxSMzOYHk8X13ODgK8IFYUkuXeKuzgVm3HW7
qk43TpEQIKh6vhqNf00//gJJrsSQslxuuzoVyWb9QuNYwj8UcKizky5eiaaZbvmxFK5/xDVPycVm
eglM2WgivEZoX2n+0/MNsoZZ+YcQHrKJOGh4g19dgwy/DsmbKoF31tWxlg9m9KaKmfkeeRznCh/C
fzRH41uzQgc1ldGNzMGOjwPAlibsksujTeOZFk+yYYjg9QFyPN85lIkBstUfERDsPLG3nC607zHS
2GT1rjASN7kKDYn8SCdtKYV1an4tzM4CLJlwIjvMLw7kwDGGuy8Jp103JiaHifDlOrFao7KrCykO
TwT4yLV5DJj5pmFWEUZqLeLtI+V0s6w4WCyyw1w3pEllmwoNkon7qJzfdIf0KFg5/LnlKJSv1kDG
F5FQaTG5alVYtAETimJcGGPVZaKIze6a8KG90bGb5cb8uRgkttmkkVcA9xTJikDAzfVoUBimvOs/
2pRPeCFBN7VAzkaS+bujRwQt5HYtvLwv90LA4xuuobYfKKSiy15xn8S+UTDj3Op/TCuaHL6oRy5V
uetyiwqKk8jM01mziFdq8qwotPz2avJBOzke+//AordC6y7r78uzWp9US/aw83RGTU2MmPXpkdKE
xkti7lv1ZQ9CKz7fLJtXsYCWQR9C7u3fmyrmdGCScH5RJGm9R7gwEb+njDn91UTSXbShGRptTJle
uWfPVth3xvBnz7gWpAM+STEs9gneb5VNp9avkkDjRveEII8Ll3aST3dMxkg4YKcy1DMozwnTCFir
TICZE+HHAMzT7opxPQDFlBJhXOstP2RctaOgwbaO9yd+yePlMqbOh+RQlKjXd4ZHB5bWclZ9jvNw
XU5PJEJZXSaKRuIMdCLrNKZTlZ7PFHWfcXNWHTyeZBfqYWacVS0BuwDAuB2uwq7LERZ/5XO1O08Q
Ju9UY/yEiKJKxMc0HbV/25CMveHGMhW8CaZz4YkA07e5oojFZX4CnxQB/KCQ/JGAF4YmpWaAIIaU
rPJ/sJm4uuuY6Xur/j1uVtX4YbOfPnUvi80TVKE8veDD3klwZFBbwZ2fjVgsLe9S7P6ZJvoPXc+X
J8rS5vC9yOLrjQpMewhZQiJ4usVIavOSeW3hwRt989FxJF8ms7DFPAqGcUjeB3AxdA5hK0whK3UJ
3v3dXz7mnyl+/tA9rlV2xYNlYLfNQyZqhd/EwRwKbr9GZnRUPUE8VP0w2XTQQTO5kL0y9u42TEeA
DnKhSHKO/KkakASTr0cWnHWIykDiwgsxHZf69XV7nYaOE5FQckuLdzIZ9/9M6zWOPra9Z+cJ0V+e
F8ZV9Npj0OBZ78mEPSN7RkCk8s1IMsvumXJwiTP+Nsk/BHWvPsKlhneLuyvSX9f+NSBKflNc5h1H
BMbV5RcQFQEJjWrWBwnCwdfZeu2CQMw+FsZ2RBzJt/H8FD43i84iskWy7FYIB8VLNHctV8FEkG68
Q4BJvFrfi1bn9eCZGGzISFXLbHWqS0LVPzzxGMw8Jc0gd3EY0HlEeXO8mfI0E5SeTfNIhhUo71fa
f06z8+ze7UzFEgjFpM+t5T/RHmsRz+vIHTUmGNpT3PKQaiZHluW58wasDi5psflVQ5e48lC4iit9
pXFB55WxZnt70q2BDyjdKvGNRZ+xG801QffsG5WCPYm80lqBdNa6fadilZ6ONl/oJfe8/xpIWIUL
XOx2B+/0HPAR4nTST4w+UWi6l3Yo45t4udRQEHVKfM7gP03Gbcj/+Bqh1P4mWzX9bmOM5XaZS+pf
lEanqFRYu3JVoyGhiQy0i4gfvF+1L/P3PZZJQAcFtwV97hETqh/VBA+iJkOoOYwQFyAlAgufyJW6
GM2joAqoNEE72zd8/9kuiW6dlEPoSOc1pdBPSCqYaXO46V0c4oFAzF/9c5NAFHHGnoUwe0JejtKE
bZYFhENSiV2FU6+ssD1fISe1xu2ANDxL6F76pRvTAmrA/lb2vg3x32eLnx07yNy9Aw0utjGtnUpC
T1httVra+5WJiv874yuHMx53lbSLGCmk5Z+Ga6dSk2yRMYXxuFs82yyWJGFj1L+5vvLcmbNa5QR6
+fPcqqtts22bXcf9OcY+z8HV6Hb9Uki0fAPjqmaSSYlyQeCYc/pqNzNWer7t36DKyWxzgxLINawW
petfHCmnCMA7JMaHJkXQR+W1H6BTmaama1Ob+w5dKgemmDoW0zyr4t5HeZO69Ry62iE1zB4RjjM7
TotnfI1h0/PfaFtGkCBIy5SNdtsNuWr6+fK7jcLCoHZXGkLW0ztLnhKIBvMYRvc4aOm8D9UIlyTw
bDFYSh+kzNZGBZR3mHMerOlU/PKyZF8+e6JINaOB3upNkO/TWvVTRdGoseSmOzcNV4aNvh0hBYBs
FfpCTgigINqtsPSDqpJXb+S+3zmyi5nhzmFHYZZQVQFZEcX9MKAskhTnjE7e6Z0gtZYsRRo8wokX
2HWPu3Rtcm21pkUz8k/aQIjhzKuEp0cnmNdVpwS2WZ+vntWyD7tdJTd59czaplQLk2xctZleGWdo
FT1f3Dq9bBABP/YuA6zls2FOpoN3VXmmU/oGd1Qt9t5RjGl+qUPEtWP+5XiO+Ka6EpHP5yvcKv5T
miP6cenHvByqLN2IQGti6bOlti07w3hqKlLRxz8cylF7eRDb+9tqG18ROuPLilRf8AfNA9trij+z
dhCjNMtxHp2ASOfkh/IDfzqRJkLxL315MG2YlLbb0rqYeauI9Ge1rl+nG9IpPHBqN9qHvTPXGVTE
qoaYYFJD3q3KcxjeK9ppJuaX81LzXvgDIJJ9GlmOdL6IZ9BzGxlhUKUrjN3fqbYPnYJoz/MzoTmK
1K2XXZ+p1HJ5+X+FT/Ag5IE6xtOiAW863fRSyp7f6qckMkK/RF6gjCWC/CfxNh5uNwPEAZejA6bg
or2Mg3wJxi07rECveUytbNf4C/dtcEmTRQz6SHytb9L1b44bn04DPGsRgIdMe/+5UzxOR451RTu6
3Jt1eFfsT9f/CcaOzb1E3XLcY7TrVabWAhoHz2eCy8pjXCs5b9Uukk3i5P7AstLlFTAvz1unhvd8
ZGfv77R6sPtmDFKQoaghR6N25fvHEHSGqSG5IV7lfTgcxeQWLu/rHma2gEKRiTDFjTreXc4AaFG+
5X30MgHrOq5jxPYsycYKO2134E+/KZ/enQkLX2eTmFPTj2ZpAhY75vWECuFuoM2wUYO0c4gOPmJS
nH6vCd66r7es7PgCVFrluAaWIZkaU5+MD7vPBa9iYRYZHMCncx4IiK9iGlZkxPqoDB6tD2Z9kN8j
CA1wj5nYS4hj9s8Su+RMF/EEBursUwaYkq6juGX38X93diX+sd1wv+Vz0YtWguHRsYONllohylCE
yPU7sySzTTyGRqXemPjNIOUtbBZ0FlIj2Bk6M02a9tf94URH+Q7SwiyMV82yhioUK9CM0m2yt9JI
+pEXHlmMcyfPlKU3XH+XcMBHby+K7eI/eROv9IkurYxiL5Sp43Eef/Eu+mPPXncGMbmbp4/+KF7b
NoXquJzc+F+aNRiB+twEUqCS7a/7b0ojR5FxJRql5gObxo7SU1kiaqB43+j9uGO6d0npthRYJPWy
/Qcxjf1SrIMIuSRiLopp5qHRD/b/1yVblkOrHhgDINkU7jDWPyvwyIBWtMtHHHWh28058Y5y667/
ctz6bU0z1M2i7oXZsoiL2vHsuidMcuWMmhpaAZsz0KI6/WfZ9j8XU9fzJE3iO1DBPwEBojuWmc4B
Xwqq1eaKINu3cFr1vbhJ2iyThRD/swE019Fm/Lc6fWPKXhl1qGTbt3Yqk+e8HkTDqWWUDBQ3byKc
dTS6vo7kQUVFmGgN7S8P4BHcKrjGW06HqtX7u9RbXOcuxppy7wdA3mqIaH9rhZnaoIBgrpAiGPyn
dH5h7XsJJ3P9L1Cb7S6fX1Orf9HlTyq2gib+KXMgHphJR0aRsDr9ZBY0MwCiYvCGfN3cFpgjq5a7
xtx1mstDIwJVA+/CgLcQ4ubCDlVBBHHWPxmrWErUJsMunIRf4C06AMFpQ8HtO2LsWeEQm5PG7pEe
d2SLYdpnGu5JFd/+slw0GYloCwY4I/wx857K1kBkAXEKLTSmvSvLuqRsHgS8XVBxg5in89S6lDOl
XboI44wMRGi8yQxkLJsDdX4Wywk4JC4N/SJt/Ilvfzc/Xaa69ozU9vU7t+bdov9pUAJCDA+C76Kb
c8srpYcODlARH10Mc0LYzPc+vzydpZdCt5kvIlw5U4J8ETT8sTenKdoL72zs7WE49v248yTQwouY
a1hmK5pKtxtpXU3DHgusyr9n+VDTyN95aebwaOQyvT6clgXKn5aafsmTZVnX4qWoEDhGmQpaMzV5
KBaueaDgo2khp5AYiwnPtGNIZfaMK1UTvhYIfD9REpT+bPa8bxyXEwKrqgysT40iEYmZg/5KoQD2
eC/oiuTwKSL1T5BraXN32LMN/7hwRS5ij9AD+hEZVVLRcSsOCmYVvw7YLQbtPd0ZJbI1qfsz3LMF
v3jWutUblN/2ogGlyOcHYoUKDVp7dpa0p0Ztn8cTrmEqzNX5VL9KqoeeZ7LTmOZWjeoi7zF/2cAP
iMXj1QmMVFZ1RGHif4VFTzMZMlkJe3nG+ljLeG7q/UgB5DnGbPTJbWGqzwKsAqwo6nh5SJNP4ZTd
I5Yi1JlEE4ZySrAVc+Lu68D8H5d/Ie3zVionbcdJz9DMTd6plb52rpCPHCUWq48bFbusQv2yB/i3
HO9wXG/DNxAA4IRuNOJi2WBd9LqcarcIIUMupCan7SBDpnUoZOMYuMjw+WTNz56W2cxFYEykmV1b
oJKJCtVXp2FSWBnreAsbNkmFaKuw8OFW/Ct2B4AseXI7S7KGl8xbazS94yzNWQ6cWbC7FimVYdbI
/PfCZbvNvTE0aDfAoPozBViBBzi/DbeyGzobu6CyL1yVc6gTy3WUj0Kdx0bM8uDTiiWHIC20vDii
N4u0Kv23XQBy4Dno8ihwAkFdYXIvHxfAwaCKW2jJ0cA2id4gvUwzn1AxxAm1PkC6sIHb7nCaC16T
aK9dgJTuowMioLxzguw0XCkg4YYBQWThYsUnhP1nPr4ksb3WoRBIwJou1dUdSyQ7BMePLYn/yDNG
Csr4vmLZXQEo+s0r0OIgxI4mA58Eg7MFK1d0SPN5gnkzwytYVvVSE/7jGkD+kuxaq3CIxBsTai8H
OtgFNTXZwW3p5wsr4MVLaD7hAva2JA3lNr7HQ+33VlCa6wWV6TcNFTYkkZK/9FDKmoB3VZBTyc+p
vI7joCtd7nXgdR4uDMgsozcC3vzMthqJGoAEC1EvX2tHrmJvcz+FE8+6jILgC9Y93UEbS/tPLZ0I
nk9MWxhfPYx18GIj8oDpRF9PQiLotiLyy1r+vhce7DkP90gXhyCgUrOVME+HlFOEIr0qzFz5bq8x
jFVUdANREJ3HVoJLPDW3cyT4WFmtkhqP+UuVOG6a/yVkuX0m8SyA6UmDKcUemKathaAPUz2qOHJM
AAVyNM1YGPwEd0Mz+hjC+mt45aJoExksF9xKb5vLeXHrXWDMDVHVw+IWfZNbQHUDyMhk7xQG10LU
SlIbdr9Dd00WQW2pkie95066igwYMRiWDfoHuT75oZSa/2q7z70i5z48cwHNALo5iy6r68QQEW18
NWCn1X77fMdJCEbdr6bB5ihUguqJf3JP5gbce6ls1OQlgGf4NXOyeuGHbDv91baG7Vx7FbZTdLEW
ySwFu/wMijmKk4bIjNYbLKmmqa3vf7IKEdYJvAgL3LZE4sXP5QNYjXfbWCIIOz3LnIosOKik2pKC
CK1MT1VxGc+AVz/dmVRucgZ9GTMF2VkLyOtZX51Hks0fyPfUttfKuCgJ3CcEpsG0j628IP2BcZd4
osfkTvgWnfbcHRcK+UY5kCDO/9ludJ7ZTtpEoL/XlFTqzSZD7NMR+5/nPjREEcgc/A1CuS+p9Kah
TInko42/QZg5EGfRUm0rZkDCHetZL0dD0JAFtdVhwGZWjpt4sPuEIP1Wlaw29oWWc1I2yhNDQvny
eOPa5OgslTPDe2PqAjYcR/STni4TUBOqBjerTj/etV8vvxSbccgO2nhSXfGXRUes+nb5nOa1fczU
/MX83zdYv1dmzAyvQ/ATyktsmwbVHiws/GmM6gXr9iUkNT95wg62m3sJ88nmVYwcQwU5D48u64ZA
4/+HRo90UU0Kk0g2OJbMmWJ+tKqYzenu8WcentILEmIEeA61nMNHqgzvaa5BilmT5zl3ENdVLjW9
I6d4i7w0wB8lK7IdwO8Bmi+OMwE9fPagsHrENkDFHwd3eYszUXHIC1w5w51cv6JMJf3K8olN4uFs
M+9B8LJd/igYGSt74qmqdD9vA0HJP62cn+Bs2IIGzIUcwXr5LfR+9Co6n6fZfl0m4HRbiP2MC+Ur
TvBknQKWgXS6Iw1sM2KFAnDLr9OrJwqMHdNu1uo/6Jad9I5okyyor8gcRKXvM+HRBEUAPx2uiSWf
T7uQHj6cqwCVB5ARG4n4r8zWqUu2LIuwIvIOHLWPl74jVvNPJPIsWlDCN8KpILYSvDW0pgmdf9D9
X4Q79N6hT4ZpbKUSagMmZTW8B+lc0FocodHpQQuabroQ8uUV+61BvnqhJ0UdYI6ov5szOktex0+m
DdONsnFsvKZBmfMiDwFlKiKhsLPh6nyu1JFwi8W9M3/n0HK/85TGpI3jdRbgg0Yor30kiEcrUJlv
TXOI5jh2bFWs4ZXWi3Wo0daHB1WmubFgBPd1ClSifFJJlp1sIdKHcTPCviPKcR/3D4llEKqbOnZK
Mvwll9jv1v5T/nl7FL1vhi/I7aTDoQYIi2o2g5RLNwncZ4lgf5RQcKkgT76qkIqSN2Ml7p2JUop7
TcAFwnXyU/8Vo8l1J3CP0yVhxA7RKwKT1SvrW9MxREnlpRk1BEl7+hxVS3ShslKnH7Asky/Q2I7W
vtBRg8gVdUk52wjERnhuSeSuqQFw9bjNXRuGZuN+s/h8XUSJO72rxo4VfaIMyTz15heBCi+afjdF
dWYUUXVj87SyxhpGDAy2g8GRxtaWF8rD9NkHWKRqnyvoJKKpmerH9nk+Uxj/tVBel3uAH3FqMrmT
G/OtSyUt6bLl3HaOpEiDj48Fb7T2jjvi/gbMJMDNHPkBiK9ZICBGb+xq4uN7+gNgVANoYFor5cSU
CKwzjluL59/JsxnPkMHLyARsxtCZXOrZQ5vKnAW/XZhqQw/YPwcJJ3ZgMRETOmaRcQbqHFEouc9e
+sdR3AkbLgXn5+iYFlu6eXHz6ERyqz0lecT06lwataqmsmRxz2IZj1Mfht7uZ+UXbbQxAjOIaUgp
p327dtJPtPbQbLyH/0Dg05EWCqdB6bcKBtmKXKxfgKfucPYIhCjSZdGte0u50Tihb2RId9RZPrb1
n64dH1PzaVOHgrCGhJUOlVRp3sfFGf4EUIfVI4fkW16QXrsB9S0txxcGC25YbAi3RacVFB81HCXf
8JtEHaxA1g3/XY358RsKzcC2dJ1qZfIOqR+CAgjv66mkg+St3iD4uv+E8Fk44NEpieD9N9lG5WUI
bGLZDxKk47SJAwRxW6HN5sHCcCMtvQf5jGIPwuKZc88/+DrUBgS/Ir/OuisEbvjglF1X5v7r0TOF
3pYAOOAVcasDraQEhJaxqfnLtX92mwNxT9kiSB1Y61f/OsxOQ06f5Rh0Moj9xp2Pql2d7KW1PAnI
3neI10y/zE3swgrRyZRo3079KZLKQh1W4uzzBeEfC+CHFa7SJwkhSzvcNkekHeA6279tAURYqzYv
jeAIKnUrwdPT3uufmt8zTMIQGc9hXnDWE5tQn+dTslbJiyVpymNNyszUv56JFNdSgTd248KhTZ+z
pDR4APLYAepWXQnIQJQ8FN8z0mYMttgdU5N6ssjyPuakNGJPJHmkrbzDDbrh9cYcRvs8aTFf8OyY
n8ExndZTzGbulQ3CtBCy0Fqri0+c2wm0G8xczHOc1323Lip07aGXT8NcTJ4/TFay6aJpAxLu1Sqa
2FkqDz7A/UNXhwOWxuAdpcGNyrRVaSPhndLfRw0VQRyDyIGUEFMfwsiEfZpVMvtoqn0j8/Rgp+Gv
ecTjeN9jEx2HPx+6jBf+5dtTPvQMY3Lj7yhyz82YWt33ul8FI8AmUrSw3ppOFN+lV8tqFkfsxHC6
IZH8vI4YZj2BkDAT1oHTOf9rIpvp+R0L9uDzGkzVJh4Pyv0GhWAqecjjJHX/+qeDGme31Deu0Q55
O8oS3F60Hs2WhVXAizZ0dGn+pJefk0f05d4ndVVhLSFIkxI0EpEm5HhU1HqLuWxBbLUKQaM/PPSy
9etiVYZ+tI2KgnuZwVq27yMLatfMxWRosQbobcscgfrWPsbNA3QSI86ctXk/JRZdRyckMupR7j1e
qyctwZtaLjt4S2mvcfyVfQQ1PbxKtoSz5DxKS3FoxBqYa7Srh0G9IL6M0drukNBuZQrOK65/r1Sc
vzIJyoWAQ0qtsDpC6U/jWJhjs3UzULfLAZmxw5s95/MYgsjfY8pd2QXvWkjNuhN0iVP8YYK07owb
O432GYcCHjgiPMin5c8OOZZNOOj9mAHW/22bNSgShp/z6bqGHtIR6G1ZXMR1MBhgnOQmWcMOm5xA
M97e5whRdxfZCcoIvX9VpB9CGrhBY+ylYqiPzs/Wm/7AOt1H8jM+3wG1CoeQVScwFO37fA/sQshj
LWbJjZlN3r04ugGux7Hry9E4orhUUIHgC5bSWa8R+YggnaLnLlrQYsbalE4sq4uas+bbe2UR1Tvt
mCyUb7BZYyc1cFFg3T+0Ye4TszlD3SxARl3kxnF4R/2f/eJcws6+ft9/OekOf9UhqGbKHJGY4YI0
aZXtqtRXTvyHOyzY6nHdryVtQnlUjOwjgxsuBELeXpCnHTiMIREGo5q1KawryG9huizjPkex/Uz0
GYqaMgLX0kMd6+k5AWJAo2+srJrizDkhAK9sqBUtgnV1jRhYYmjJawRrMtqq2aMKriDFM4OclMGy
+pSMl1W7HEygj6tJFrlbnYHeaBuFpaCz4vhmR8ptxEmfEad207vKbhMBoLSCnnehw/HGf8xy5WUi
PwOIi5+cL7QKxEKMKIcxHlCBlP051NC32SK3cWNn4Eq4Hr9MJFgSFARDnuWRtV9cZ1p5munpIAcu
3eZ/K+GcqIgLUzHCtA05tD55YVqxNfqwQtEd07UyZ6+Uq6Qjxuss10/D8rbq31rC1aYP5zf0JeOr
pqPoOt1MkWFoV4XkT22fRsEbx8yB43uFIHaud5QUjdD+AaUm7Pph1NnShZ3DPoJR4qTIVh8j8dOe
TY+P5JvDJM5koNVs/A7i8btzjGMO6kZDRxEESSQYQ+ZNvxDYEXKwceR4Ihh6h75VL5QAOzy+7EmW
Ht6tVewzuHYXhry0jtSqtMRO7QaO4HgcwQuwuOX7bIG2s97SQc4Yzn/OuUCIUMGOgoIkhGdAmVPj
Vd0q6bVuePH3n520BAo3HhfrDZt5QwQfJtS9Lcq5RBzBY3AxXouzAKJP+3XlPjvvTZTpk/LeT2sq
k+Is9SFmVYOZmf5Y52JlxXbzNi7H/XSvr4n6vAlysu/itKI/dxrULgqst3J/cczQBily2kqD9mrN
etsnveyrIUgT3OoutjwUiBEMn7PWq+sx+EaoLHD+rdhmIwsUo4WNJCcE62EuqSu6xM6XphKhMK71
/yGZGxww8SrdXg5ahzQTxyWq+cNWt+oyMRRfM/Wjk9yCqR0VNU+y/vfx45QPWnDa/a7X8L3gEkO+
clGJlyCehuSOLxt+KGLg7wPliRbtcDMT/0U3R2GCiwX0idLJTbWjNA3Bcxr7Q7PcANbMFcs/kXq+
IMY4uwKEM/pxKJ5xAgSVE4n5uUYDT8C/Rn8sOX9ns3QLYRr9BjuK2qegNdt7EqKjC9RC10fKH9S5
3A7QtiTbDGeiYFxLT98LXWlTRBJENJMXv0YT6MeFib2CfLr0NOKv33gcGuDy07CByVbpqpjgNsOh
SerJr4Sp7rVgfadHoEiKbEhAs7fQBdFWDucN25IzScuFXaIs1Y9gRwUG36vjdHP40651e7FlZK0E
pPNTysU3GsJKIIZU9OZn5J+EIm66ffvSWwpEdmQAz//fzAKna4bNAqPxDzuYYsULAwOL0cj9U1VV
3dXF875K9K1FI7PBbWNnmacXA6sb9TxP8dL8FPZDgZt7D7qSbGNw7j8QYN8TMJqEeM1NLz2c8/Hw
qfG/yjj/L/1N9RYGGLb5vHEG0upziXzUVqsF/uXO+oymRegv+3GZVhl7Uv1VV4ltffsoPaSqREf5
CHr66c5jot81CwUJO7FEf/Q9tYFu9GMF5vtzwKqpLPvd8C84woCmzmoo27atlIGldZYfC8RCIaXR
x48R3Gh0YBGk0GO8j8j/ltbjX45qfGrA1GEGSYAnaXh9BsKP4cKQs+noj0KKKaYGmHxWE5ZLSI/m
NDspbfC+MQO0MyPypHdGMWEW60lKR/FO1kK/zUAWRE4gMr/YC+5ufL9TZ36r1/Pi/m+C5iURVLDo
A4pVuxd8VIZvL5PPNvPUppP2Xuht0hLb9W8quwAann5dPqkZF6f5hogWS5NIcOiziwhNxCuB2v7h
x2biWfn+ASrM49U0sKRJ+kY9V0XlximxZGRV7kw0HgulNR2vailrLC3/2t4XP/Z5qB8ur8BRaN5X
iSMO+ZBwMDQ9zNlNLhfzUtTbP49nAc6sGT6xYrWxJaq2y6tJkNRy4tiXvWo4WPx2krvFv2Amm8a1
Ddd6hPAD3LSybhkD49iJhfEQ0QV1xPaLOYZj7Xaamf8SPzjLBCRDo0bI7mDMYbTeZD4l0fyGDP8q
y/vp8hIXAsu+cc7lggd4nM2kyvUxL/MCeLF1sgYDmy9fLDWeFIPMTD43snOPjrxjd0zVWWduEQgT
c0OVIbnBgMcJmXQLEZIcZZGpElm/NVL+UilOGSr86ai0z2Msqa+DTyX/IJPBxGHvu2CEOsC47P/2
5hbHEl4tORhPWrWmRLBbwQ8AbKR/tt0tcaF5v17VffxPk3mbN5a9DYIckc0JopdQq6WlRmU4M79h
04ZI+B/C6KZc8uL7DhKgiqM+nM2EGyqWdw6z5087SDc3jrJyRymMXEKEW6Zf9aZAQW3qeUYIfMGj
5Or4rPLQb7TYpA+0Jhlmmsr1OlPW1aeHGuyioDEjD35ofdbO2PCzUz8zt+/PaC36zTGNh/sbMlMD
WeQpI5lMBE/5bOISVqY95RdEnuhQIYoo3hS/m80UWmC5OklEeXv0EeUrFIJYYLR67vJPY4BhSC3k
RbY0yVFhsSLRrJL7KpAde4HalbRMGxAPb3M2V/OVQgmD2fFEJkEYkeJ6sslKAt8VX0hCNCLovza9
bO9PVDV+dbn1rE5UTqd5QhYgvzSZrny4eYmFosKHvtO2zUmmEHMFcR/qoSnViR76SmoRsqE8bLWy
zIpzJniOp8PrDj3aejLW94ERHaquLj4eKsXWxXCVL+Myxr9wt04R8HdcgoF78k5NCaFZsP5uNCIG
Pe5Y0oLzARHuf61Um83ZfDQNKpCOlkKrirnaLZtO2bTGdj0pfA8/uSqAQ6cudpgVAoTf4FpPpYhZ
0ETnQj9i6ak+JqDJYJuUeKXSdsF1GGfcO9ziDGjcvBrHkY+7vB7wDEJ7FqLi/FxjOY3osxPo39pd
VVsSt/fjX3o2XCz2iVCIpTMT+hcO7AW0UF9sbTQtzx3AdLM5LDtRbcuXTwsethYtAr2rGRX/ToSM
+K6o7ZECbHzwdpZXmFmWBqnZyuHnJQcM7qRwtAfeCHFmLCu2BNdqL2ZB4ZXjqaEd7KVGjbJaH7Df
hVu0kLxWTVkMBq5a1nmRXFAklYutcaNXMb87hdryd4hf5j3Iy8HRH9ODctn1PxlgnRD0cnyQ5sh3
LFsP/laxN1t/dsX34F1waI0wA7cDb3XQRiWRdySpb6RWTn9IlJPlsugM7pzVcdkXVvsGu6rYl4Vx
yL6kr0BsAHMQJ0rD0J1U9S/XiCFZgOylH1YAx64KeF6CfX+2RllIRTyEir9plPJ3r0/xu+EWWLqo
hd2KwrI9szincR80aELN9xbo3tDVLoL7BfQ274Bu95Jls+d8cwE2KWkVqEIJ1BiTgxb/UmeasdC6
7YDsEtnUEnNZy1ExJwC7fSCRU+sZhMRz1U46BB3Rp9Xy45ud34PIuY9KUkwsmqihMG5rTLPz99q9
oWm/pcH6uFkxoi8dNvz79pi4shQ50qQZUXssCierkdvgSQRSuPLS0MStsHAukpdgTw7Tyk54Kj/y
3znYUYemuMlP7QpWXpsZaWwiHPqzQtV42+suhH1+mmrNi3dXq8W8ur41L7Uzi4hZQ3SCLQ/ZNRfg
rJhN05szKdeyqtyNiBa7OSY8Ti3OYgf/tRfgHsmUfGhgkJ0oLkfJ0f0QQ3CxEm0pX8jTwClutyPv
n9bOR3m1dSF2Th7K0dzqf0ydkmnZt1iQhmT1Z12JKxEE8Ci21IXag9v5SzfUIHnQkwOitiTmVqhj
vRGjZclSA7dOcVmAs/9p4BaOi3DYsiAH8rsE4FqoLMoW3oShDKb93j1qxqDNTe96ljJ9se1sZoSr
f0h3ZB5yfTG4uA+VhQCnY7V8CGGWR9NtAZRlNK5mx1WYFpauBwRNKt2I6uTmMEroMU0JpFv9Jhma
y6KhnjxdTKoDqmFFErStNWmzNalL9ttJhbgPJN/lRNhToBF5avGC9H0j3ekLhEXhU/do7+O9hZhf
Od6B2xOqbc9rlbtcBD3xg/xCU595mHV3rlf0OkXvOIRY86fJqZ5B1Y8OXf6DgZDCJfNA1SEcrI0A
oYwM1k8nt508Csc7Y8DQvq6GxrtKsTf790V8fCdQ9qWhpDM8QXYBUx40zyc22nmJwNscPht3I1Lk
UrC1oRlg6YplJ1xJDAcwrCkEdy9UsuSuAzL1iWvM0Dhee6PCz+7lLwUSzK2FHbpAzrcPVyu456dF
/hFuG1Rp02VzwU/oyfVrSWK46UwYKBAyy34j6sjapFkjtrfvQZl0hTtvY9Ys2z/bwWXnx+wd8fEQ
niv6SLjnr+bpOG95qXMEzYIuvkOzsvMzoUIBF/y3F9nHW4I8zqFZXMN/kX5hEUtaGNMyJZ+JNNcI
kJc9Xf1sOBIjtOyo9M4qKzZAqztYyOzLMIqJrf/hmc0oibIsZORHf8Rz35JFiaEX9Tm4dX7AesxH
lRNiqw9B+L5yKgXi4LPf0dDI4o7Ren4/0WajyERg69G5S+6As+eerw8rxTbi4hWF9QM0dqnlZNsR
mYvwsz4uIdyvsbwqAZLMvdsMwjWarAH/o705ahUph0xrpqqpsOOYQQLV6I2ReCmyDb6eLeESNgi3
wyQ8dXJxtzbxu6P3zvoBw6YhC4NnhxMNtAzSRXuyX/VjH5EgUjcTVRscEgTX7GSKUvTqfloHWAdK
X8qm2WtTsQWNB2Bcg+b81J/2rjdHJdwUu1MwR0Nv3W5lFCktat4qw+IUF7l6cSIgEr3Nm6ixpSpM
0dB58K6Gjkq1p7PncI/GH8tItS8wiSKT8GTZM1flAjAufONx6lsCsS2sF2o64Kr4/ESThYlC/vaH
FyxCJ9TW3B4zs80VKmPExTBTlU5/wW7xIoFYQghPHtTMTw1jrWM90EVLkBTwqVEoclwzhWpDa03E
4EVpnlV1uqSOYMsGcaP7YMUg4Eqanw8jAIQeonSaBB+x4KnZvQjbOezggJSNvSLsMWIlluWwBNnl
tCurgGlFLUqr3jbrBU1E1mKo3KbWS8pFQ3s0gO41fMs8scOaXIHyvosmYBN0tQWoXrFWF5zoJNsZ
jDlMucsCVfoP62d1HVsmmOsKzO9hD/yTAb9YKyBwZNBXsSEChATeUEpOciywj7t3K8GIGn4RyECN
Z26GUV+JpQ4zYGkFeFCmpOwM7d9ql+UFsxS+G85qdBHU5Zxmw7eCx65/Ds6fdezTaQsPJa+sjuqa
M5glJBoMmkNcatQ1R/6NktXG3NrygjIDNO/W1wyyEXjb2jyzPINGnw0ED3KBiLQkzxzeQLTNc88f
a+TR3E5/U0x7//DBPWmBfVc17dYv5NI7+HeU+LkQkliujGx1+GWeaI3KyB87oGhylnXEsw2Osmke
9e0D18W0F/2qZ5p1Inj4YsFAg/ICEcFonbIJ95YTk2xIIxldfKxw5qEMDF/s+P7YwINXVCZywl+6
g9mMdjYlt7S4esXr0xwHk9X1vxwPUmIf1MUBkP/cNCV4DvJp83YkNWnmPSpXFbpMwlor7gbPqGCF
W2SCsUIQ9gNYeee2beR4On8RCFPft3qu9p4FgCpPGrsO3fwp+5ACQEgLE9EqD7DW7xzJWsewVVvq
lhrXRTz5R1Wv5MNyM9o5GDN46ELRXkX7GVJ8wd6C/MlF74JBsPZ7mkVZDKdkWdz+Hev/D7RI/on+
rOOSRJah9OV6rnto5jQNwyYfjZ1pSBTmzoa5yg++sttVL6SIjWhS9IWd41jZgeazE3QSDniQacJE
MusbyQZc+FuJT59hvhgJUmBBoYo3Er9AI2BZ1q8gn4MsHa8JjcW0f48Tn7wUAIMIwpe5njoqCbmU
eFfI9k1qQk2dOc09oLXzqGvfp0M2Jw1cpwGs6WktKwhJwEI0lJyAW3QUzhRqNwWVVfbHtnjkieJ6
66ELRtitl3mLOjPpNtHUW46sda4AFkph1NqGVmlXe6XMq4blzkZ4iAbn/XMcAE1XSS7tu9leB5NS
kuB+1rzXhJE5FCjOM0NTEV6g/ObQZgziN0TonOZQSgN12C2bsasG46tZYNbJ42Y4o/2tgQvqFACV
4Av65iUqPqdfFMC/9x0X03DhkCRkx8oGSYvnc4BkuKpK7axAztl3B+KMRJjgr/JRX7YOBNi6Tx11
86iP/KCrVT2FJjrdzuj9w3dJYj5EyH3WUTaTymKSt+tAYu7dVT8CJb52ogetToGMRRXv2Y3l7i35
iw8Y9pYf4v5cc0oSMv8ABTJfwuWz8kb19bHBwOj9h85mOwvH2LfMAF+NAG+GjH9volkfl2iSYqVB
/o+Vvetk/PV7CkXnaUa3Kmhkz6kbPTesYX/ZCiCMcXvqzD7oFcsXF31osqf7J7Sc+UdHeeSu+O2G
gotyROyqd+8FA5YeR/yq3Vv6GZX5cvjnDa5yFc/VEnrJv1z01zxxrqR3k1k/6Sw9lY6I9lN22KRY
43rvOZr0d9Zg/49zLQEivzI7JMNoZS/h7Q+i8jUZkgEGHL33646xK5XNFaWeoVBjQmreProPJ6Je
iS5lKlrZGhixBXGLdWEKpnXleVz/96CHVnubA99Fp6FX12JRtspeB8KiOW9g0OtwOGVOWwBmFxvE
4pFqcBTmi/GN5V8duw0t81/nDUEZbRIiY+rTN5WNXKoFbed0NAGRYrlfEyJyS0e6+9rgCpcohwpu
YCe06WDeaexFVZ+MMyBta/xTIKWvrKGUZQzgpY+5/YRblBrauIbLtwACE2p6s2oWdcfDx7QkHD9x
84M4rWrGs4vSUn6UTarT22jJLQNJ8aW2sIGJ5znA0UmupyjXJB1MftmcyaZz156yNUlOj/vtK606
mL78idTf4r8UQVzH0jIY2GQc0cIdP5jlB6eUkboFJKwbWI3ODhLbIZEWdTN7tutN/4rrQ0pPWkxX
P9hPSRkxWPQ6QaEFWz5+r5q+0g0yehiQi0SsBlrbVHqcyDWqt9yaKbhQGnq4cwuSi2BwfIPuvZxy
+SWPu2ysHA6nWub3RoFNpVF0TTLtftKuQ6DKqLixcy3ATGrK8uSrepA8uUQop5Q9lXRyEQUE78UZ
bKob46ZU6NYzc/zTEKhHDUg3gn5vhLsz3M3aBBaTrfqkMhFeihpWXpB8wn5VS0lNIplyZxViWKXu
RzgP1lV8eSLDwmM++YHEDi9eQGkcsWmAi718jKdZ60mPTaOqjDef4/ZmHJiDvqEbDhFA3Hppbzib
znfs7rRX0KL7XMANOVFG86qhPj8zyQdFgOuMmGzF4MjzpTLcQl7FEdRVrJoPLwoOEtKb+mCUVsDQ
QKDrVvsI9Rp6+7FeuiKZjgk6b7TWPWn2jWFEdZSOJkqelNjey9Gga9ENiynISL2AZh3moFbjGS6S
HE3BZZY3yrVERK1Y6Ygp3ZMpj3v709qw1cczj37Pmt2LiH0WcMbcFyjtgVh8YdLyay+JkryqK8QI
DIWkhwX/Ox0KCUqI7lFUtmAvvNk7szIAkWk/sJf/yiOtfJ+md5Xg0p6UPe3Yc/EvgVC2VdwlxWD7
1gv4aQTuyTRi4aseO1dCn9phyKnhgJtDBhZqUfY57ojrZisARCkBKD2IpuU/L+sOc9w6L7B6mDQP
pYzxWvFhu+yeMM3vgOetP0x3UOHAW26dCVTOzSwlM3JNbMBDvSkvnqDx2YS/dNHT1WVxFcDPB9cu
ozc8R88BAO2YL2bWY4siWvlSiwBkc49UpCt6roq9gB8oVlOvm4uwHTBzRaOwaT/vPZNvFQSnkQvR
N0OTzW+sonl84YuIXqa+SFqmMZhSAu1RIIwtCKhs6dg2xqcxcv6wQiwDZY6tUKvjFqrhjxJyxN03
XB1uUdhiXwUkxCT/Y7HXkytr8UvRyum01askyun75JJ6JhHJq/gpzp4h1SXwL4mKuxAVnlFdFyjX
Q45filCzDcL370X+kkC6ZnKjYWLeny+6rqSof+Fk49unemmDZ8VKdkOZ7IGEn2YFYcfRZRhCKYCh
719QVEbdGR8yvVplrtryY7dQx9XFtyL5U+lTWSxtaO/vLRRvZFZRk2MoKMKuRkawqhD3zeE/gzy5
Sh2MRDybtkD08Xhgmz8hIOdGYHNFQq9FBi2iHPM7fliuV/+T4mey7UDQ1jusBx5f647M/YzQdPAA
yD+8XB/wR3qPCcDRjd4JSOwojgymVYWIBAMyfgQZzqUghCYWfvjKwx/NkCaLHWdhnkfvkHl+VVwU
sMxv4VeKcXJsSJ397ODOFv3IDutPWCywQVD15ciPFZQIwFR4wFvgiPlL3f06bT9QBGtRsTQ5Wv5J
/QiFtssYZqTmYWc8Wbk03r+AdC2Z9Hz7bWlJslahZ8h1dVUcY/zio+zIn9bkXOxyzhmAIRQLlD35
Y49w4emd9n/RkJZCvfL19wRHbW3UOEbZaHsWam58Ppndq9UlfiM5lXad+5bb7axESIr8lhFofRKI
nT8dHHliHTbZXaWet+KnK+63x5jd2c4UaWWdYD7V8vaCecMhMQHUXBkIEMiQRmUkWVJLvMXCZINx
eKuKSZEonysFZx7e05U+04B0SQ+fCh62Bymei3B0ZxmMrmz8F0zWOTli8S5mtqDrn4AscKvu/IUM
u8NWoL+E/rHFbF23wLlQQZ27FpNRwLZr+ZCY4/3dq5LJmlEugF+UZ9UDvq3QvVgbLebg83wg8k+t
uAGgQldVEy0hKicvKfaTZmYVj8P9vIewoo5j26SGDbpPh1AwdCKf7v/ewPicJg+/dCaRgimtHmai
PlJQi/qxtqN70YdJRs9e/HX8ZE8w8Zmn2laESTXPEbTwVGSznHYDzCoTL9SVYkUWYZQ0wVxhRyaI
L5CHhO1YHAvPNtyUXzTYJf6LImU3UeYDfUjpD6zHU9XWvwbbkR1NoWgaqjoalWhtKQ+fz0hqXOqt
c78FMFe3O2235AeF5zoP29Akeuem7W42ufLCiYo/8tQU/pxGzUTnff7ksxuKBoNgO07LjCQcfG9b
NI6uFk8HVjPWaXfn5+W3jDitIuY0x1U+29ltqN9kvjp0j1Fwxy/OyZ/1jAKhvwQyYCYSOK4FOSAg
v2K3WbHadSYtleSUJsDawl+Lh5y1Thi94eK8B492RnbVPwZTOTiRnVP60JGh2UpmxjwGH/GMu1/5
BDGBshYiZRpZ5piOW0hmbbpDyaSC1WV8txt3bMSxORfBsKSbr2PrhngDo9qZdSqwNT08pFwDiMA1
pjZnyqyAB+fNepTpqU0A8boWAiAYHgcOpFQKP10OOOpEiMw+crRdawMI+Om2CZp6ZasiYnxvMsSu
X8FDjn+QwGbEoo73/daOjLrQHsMKSAU7lAnMZK+tx3idxUnrBp+SRr/JjYxM+6yNbuviZU1ykV2Q
AAsTnxn66YXqDGi6NRKc3tksf6GPQMnaDv4yCjsrtzTnBB1idMcBGQrVtkRUiR9cQl7+Ewd2A5Qq
C39iiASEjuc8/pn2fuAszAqtKiOdzDRt0os+M9lTgMlHeuVwX8Mx1/qTwNuxMKtKbVFYP06qSNXy
ukuPe99teWO58QjkrqkPMIp4JRJWzKW2NKDnyKhxvenTcAbqrnqdyHIiEZtq9ujGMoCpNZ2T8BG9
AJa3sibLHNpc+zoZI+YSde0olkI0nNreuceCsn+w7U0AFubGJxerH6PTNBdOQYDngY7mP76fdSLS
tPMZ/Jd7CJFzWPGbP7EhlXKMA6NSEYt1MzC0qt1CQwqTYt3xleGiQfZhmsxuJLAbh87kQiqbOBKC
IEMVMZNxD4jmV5+QL4Il0xVXbPyAkEaYNrNO9m99jwDdsVr15AQGVfxxqIDH1f06UrXgHrdHmrft
HMLXEd9r183l6bn+gw6z8MA8/ycIWWdHjK7ljKBq8I3nwJ11HTsJcBo2OojAppHYydexhg/Cztym
fmFpEneZosa7YqU5P7y3We9RBRxlBS3IWd3PtlKUkAos8mD1TN3uD6lTuuEXFI1Rw79bUR7ruZeE
pVQfsxlwbSDbvUXKRYu9ZezUY+Wq8aHYNdChozBYv64RgxbrbohXZeNA372Xzs3ToCpUFyNcBMJ4
4+XrvWdFP9TH5ganyjZLz82StzAFG0oDoRCc0JrxVM5DkR/EEtG+u7q0Rg7gHj1i7v6DFHwW5zmN
BKJ+UOO9pPXwKeWVPPnde/0va0G2075rUW9HoIrL7jOMmnpRA8xQmlUS0LCktsMsCvT9jl/dieL+
aXmcCstAK/nxL83sKsj8HotBiYsOWtJNobk9HYOPcLqYjfWpeqi/MWP2DQaSBsL9d6WTqkhU5wEQ
zf6h6U+2eDuh3XEE8ZIOsdFm8JgiTi1c2+ksqkyHVukogRPtTSaN7lnYYW0jvSPmVxRVNstIeDNK
HdiZBNVu4lV/IJiCDJ5Rxd4UBoUUV5FXH3ChkoC+psS3fyYQIjv1ITTArpIZ05iSHpS3eaOcX994
EIuZx1y846luGh7acKI7XY0gLER11OZUAWVzMrJgk63nZZ6KAFqTVQoFmKnMLUTJ5p2GPnrK5mVV
NxnQ6iJlVjh7V4d6fdJvaJhv0ih2RX2Z6V6Fmslp/rWSfQzP6Uoxg4WydSUwVx4ysRfB33ht+xcY
QLYV4C0JJvsE+iZPA0pL3C2Gcef+tLMj1v2vKeB3W5Iy4OrhBriHJ9y9P5+pxo1QjM2ZdJNkatpC
KqLhOnO1UD/IcxLdSihCHt2M0WlKRNG8//+KWaKsb9U3wmTuucK2NPbHjzwE8JTeEZoR972oBL4m
9BT/r2ipuBMa+qJ6rpm8AK5VB2YCu+eCIhia/2pztf5OzHLIkGwRnANVwB44WNnGjW35IGi3Y94y
6o/APFZHmKbwSMfR7mcW2cwJLAlwPLfy5mBBTCXLiEQApIxmhVvXcnGtWv1HamoL6Nd90o/0wPZJ
mjuH6CwqJ6M/P6AR1BV9na85ue4VEjEmHFHJlmXMIQbonB7Ho6kzvzoFPvha8/6KxnydRtSsYHjd
xdBkK46V27Tc/FPyNHnlJMdTnZIqPwegGcnKCEnR6mYQAxCNTxHCNf93LoWQoIfX+NllXAnD/DTX
2ukfpWgfQvdlKVTXmrPUSUtKJemnBwgSWY59YXv2ITvzAI2ZRGlZlLTP7M6NpowBVLodT9WAFtxs
Hyc+g9hc1DNP0TLXK/STZz69flU1ydpIN9X6NreNkQcbHa5Kbtts6nVhh559C0f0juI8d/hr1V5N
WpBvnIYton6QCzVQe2aFMr+P7H2cvMDdsXQm1FxbZdeSMYymkVCDsmHpLNYdqRTF6HOjsS77BcDY
6OdZcb0Sty8DFyO0e3H7javl8HGWC9pc9D08Ohx99w1/NPtbg7eaEP7FUnLyGjRK9naye2UHkhIC
JVVOFw4ksZd5LJhpeYyhW7uOmieyphVuWkggNYpIwyUooZE7434vunnVB9l6aOsMH/uD0Ru7Qu5C
SuSTYdIq4xtuG/5qJOeaJR+9BQf7QF9EyQRYmw/xHiOTyH1TkXp+AMOYs+wq9gnWJ8tc1rRcuu4f
f3/yu4Q0rny+jS7qPc+59dpdWP0iNIRANlvp8xa6M1AEgp8leL4LeH9s6IrxVvauWU6t44zYpOH+
iS/Dh9g8y5Iae7aJNT3g2d8DIYav8+tGs5Hq41L9udXaEqZpoELdsefPGzGPzX3VXTjRG4Te2rBK
wmuH+k86wGnpVrD4Uy9KRxjkiv4GMLfBFE+nXUjS+ViKmIKmjzckwhKXoZLVyHZ/sf/2/2jqwUBx
ch4MEj05YNyfxIYRSxu6W9aahX9JSDEwM7bbdgPpz6MlN3IpaHHEd80AE63z+Ooy6eQsJmfwJ6+b
K0NfAJmV3AYTjfi9ON6sWCZdGnsPWMT8yrZslaICdCjs7qavWFpZMwMyS8nX/p16TaGmk/kDcu0k
4rRTmo1tC4PzO3fXIyjOVXVyHMhy/7/NIfVz9rT+X3LnU7q7naTutWiEQ7zg4TxdTwcw47J+lGT9
N9bJh+kRYrLN/mRhlcan8Ge8/XAZ1dr27p8SUyMcPmexjxNlSbbsgMzLBQ3mDJVVBOjPttmuPJDa
JnRjqtwNkUvuKjxe++Nr+PciOKoeyCFouQdVDwJE87+PHSI1r1m/XBIqtfKySyQe1fC0WibEpv0m
CJGN4LCfU6fJ0rOnx8JVEqLvc5R+c3PVpc9bVadoCEWfJdg2cHmF1ZNwKz/uB2QNXK4k+vmZBxeh
i2ivcBZ4XxUxqQUVoNrR5F7FTgxXWPxbXX1w350XrCNhQ5PGmObSYoG4eTEZBpNqDWAhy/zSOW5X
5559zHCydVWIZOGWOsHfolltoGRSsXpwgJxRqJZYCvEvIX2j9vi/KGlrghybkMqhoWkHKqV3wr4E
4IdUvFMdSewmTtNs4JRgHJvXbIVtlDiKoo7hFZ3HMTOI15Y25zLjZuxB9lgD2ukr9zGSjsd+S9fl
c87eZDRZYpAiGfavpdvbQKd/USo8llUDz/OaC2YxI7lU7Rb4u4ougpHvnuiAf9rGMUzfg0D3Dye5
NTOjGNh0ffWHNrH5gMwLZzeRma0IiElE9vffCI0oC4aPN88IjZ19+3Qfuju4tyAWNOldhH1IPv0F
Qip5mNlp6Acu1V8/o74hWfaYcIAVRMZZoAjtoVHeXVB4aWtR6uHs7WsF1cRRD62hrDSU3L+Y9VN9
jFl7C2dbMcth1YmZIXA1tz2piHS0I3POMnvNOFzpjY120FTJ8rPPC6XDE6vHCgg81XR8dEgEeJpt
w8jOY1upgFHoSxckqc2b1hydd2DN9B0I8FnMIfiTi4X/XANK+TeklREtcq9bwojUBmOWCV7IXS2A
dq8RRqt9vci8fX2xqocV7vwXHX8nSR0/S/D9LTul37we6ftpRnEgOqYCS7DeAuM2uaHnG2X48jTv
akhjH2fPW6lRUfuMBlej8vD20d4menoU+q5fEt/47rWgAGv9EuQroHUMYwF+l3CFOngFwzs3aWBz
yM8tdQeqjFEsjHCFItH+zWFB2CP3kU2t8lLO86xvYpINyWqeuwL2B4MiZV+JSnHgrobrzhvEB1lc
ZQnWdon20BhvFJm9f1kpTnscQqLoGpMZviNDQ3sFSxfrn8h2G0bNM5XYMK/4UvTxt/iwLt/jEjX+
rEeKX8XyQw3BbU9gtuXtXvleWZW86NmLKRBlQC20CPZh4MgOKUOqrhxIHLwdvDohHAzZmZLIEcfy
fQI3QI5Ym6J7YNRk/KGNE5iNtBlxCxJhMorbp0ROTwFWo5GPS20bQSN6PoO0km3LmYuR6QaJ0gTo
kRUMn1jvd3x2fNxuMnujjAUpWgTVHzuF69VxjreE+4nQ28x2GQTusnSlA/05GNQ/ywOgfAqBxKK/
dbM1Qewk13MwmToQ2TUWieGeC3O9SB5rzUmtnw3XXPJoEe4u4kfdVyB0VSMtY5v0duPCBMkTxaWR
eSep4gnT2JL1qYAL2AtYGFcuB1lw9T1OUDyganqevF1jcstC5oqSUf/1wvbB48eR+0rqpHs/jSw6
ij+56YU6hbvqXBQ8OnmdyOD2rSizhTE7M52s7IxRz1XFUGG5sfRdiOiPSKA1V/QNCBGIguctf5HI
rdi78lnBjs5kcHXhHIxdGlt+2a6DgFhAePAZzQM6pr/NidJdPNaZvtC+fQkPL2YeuvdSBsB5Mh4y
8/ypgVGjpm+ZPhXW+Kn2Iwl89FL0ueEroUPp2rQifCXMbbZADYnrptIGbKhXMHFe/8ZYyYYK9A/Y
0FPGqqtK7n2WazvtE+diJcyy4ooVi0f7PyeaxvI7fIBb/bk2x1iWJQYrCf95FVOgWRkWDnGWfs7s
lHgT0p3MRp3dE6aw2XD6ma35E9k9G0YVE3W1sTK+NBBYn2jzcnB9b9qcnOqErf5a++pHRl+aCjW+
2LOhH0C2wd4YyZ57g9h08r+6wwq6FCC0kve0z0USAuoJcbzpI53VGnytQQTy6C6N4Avr6WCHmL8R
pId023lfXPUoG8MTh9oCgxF3kym8Zre+MW+efMMuU0y3TPjyMLSa8yfnmiUf9Vvelp9wyeSxYPHW
teNxciKxGUBc0huum3V+B3JKNcKzGdMm1yyPeHGascATsBNzFhw/TbAUIRLCF8szO0opz34wETHM
59Zm1FNsSU/oTTq3ekuHmFjW4aXl7rts/nPjQniYtWn3aGkVZsLvC4JgGYAVoVayx+yftdNqZAgs
s4IyizJfERtfTyeH9hN04O7ONaYZD5x9qkfdxOvyO/oa7SwX50T1UC8Z52NAzTrRJV8VCKpc6S3e
F/8B1l27gamAKoOsoD2SkOmMonSFWdfVXrMWaI2j3m48JrLQedDIxgt4tN6j/ssKxeB1BlsLqlaQ
N6LeKDEvIy7acOdX8cG9oG91DNJK+yeeAsL4mYyelAdYrc2LhaxY1pf26370PGTOJ9NBQt0GzWVh
U71xPWH6z4ZFdAUw8j4N0AYubaTDCJ4TcIXjOq21/rXSDlBGf5VyWLWrPFqvQUOXystCmSCLYQzW
5iSrTVrHbj4qodk+isfRHDZfJUrGMkZ84Pzcniova1F5U1t7RHpdbFOj2zg/X/hjcDAvuEq5WhMR
5jz87zsDfIs5HKn0SD47cvgiZUmnsv4GaBliT7Unx43UlLDfWn6TkbqnH3co8xYiFEO4vtuKeiLn
R5VoAPe5dqXk10ZMDRCdQ75V/uCyk+4DzAxrQL7juauViNUDa4mrPd2rBEInrUZECVkCz9+WINV/
s90eZgoIPDEXtrUleWIFD+ac55Rf0oiqq3bmbGmgAYo1Akn1dGwYNGJrbKi027sL4JeSZqCHNdjh
raPGrdvjftZ2leY0WIv20i18VOoOL5EpQAjESfb8IYguDbLcbpuRl+Tlq332z+EfBtVctJZgZs93
3QxYo9UfYAlgIoIsoskTBEjk82skD6ndpt3t83upB/9LubJO3oWK7GgBPxCmwuNTKEJ0RfA9gqXs
IGIVldpovchWAQnfIDe5wiOSxi2v4IA/0m58jhwO044jrFmXQXU6EbeOk7ZZHL639GDWfASSFr7b
rNJfThFjYiepTg1PCVEUwA2K5VYWMRNv+jXKSn0rzcn+kwLFMX5wRO/wuvvt7M8Dw5wXADl0JchZ
Bxy/S0vPscmMQTUPgZjmsBS631GP/ShKW32Q34t57xoRfR4c1KXyHpDEqjAgI0Sg7nd20vXuaYqD
SHY4wE/EHujfr2uTjcjVE+w28Oi58oB0hfXys5UI0iK3MWqep+9F0IWPmsbbGzpH+zKrPZBgG8gH
A5LuS6asS0QfbSlXR1krmMFLeSatl7dELUVGb4Y1QqbCtGBqQDd79KzoUh8RiP6OIuf3SwaNZ7SB
85VKNqACW3GpCqCvEyGTY5AorC2PZ3wFZUpk39TamN8KIPwNm0BBwUgrkqn2ZNNyji2lDEGGlUdj
kzfiQTVTf8r0vg1eXzw5Xo61mfdQ2Vzb5GbaF4Pq76XzSdLe4gjlQJe+6UiVDlQmJl45fQVBUTBA
RG7IKwokSN162XwOKzBFM0OF4h098TB5M6zDcPpbLBzd4jkAgBaJdd8VKzzYZHWorX8PNjzXRd98
1TAQbJu9m/9oUXBkgv+Gi4Ud/4/wD1QkEjJ/PYylFA6T+5aDBPcQKprgvLa3s4jlwwGcnbV2/yC3
tPIGMSrbztTMfRK4ttkHj1hCLofaLIYzXuYRXp+BbYv/TKF/8xWgFBWmW0MbA8tV8EgQYrmqUnsF
w7NJhYca9PyP6Yk5wrwpfKfNSgl9radBCoCox85j92RtcU8mxvgEWDiL0cdb6kDor7bAUjfZ8n47
sxxFwWxySMoApXo5Ao0Sg66rPepXQBeg30qZ2cdD0z2+2ffMDz4SuKqZKnAERx3494Gtw2Kc9phh
7L0vztR14UD8wbna7qCfpkNWpKj9SBFu0U9Pq2Ww97g45S14ESJcueAG1X+mLONnpQYv+KJLPtoZ
RkyCqnmWYpHmr5Hx4xOvibxLTL1otYNw0qqKHkn9g3ipgnZ2aed2SANpQcu6JM6n/olxiED0uuda
c5C35XGSl70iB97keZ4T5VNV6Sr4Qb6omqA45hspFCXvWBQ2hVlFTCtAW/hr9+GbduJJgnAE4v2i
bisMidVq69rrdN1kPq+/JGUS5dX2MdA5e9X/7e0xAcbzw/9tB5wOaEyOrzM9OvKrCv+95CxE0mfq
N2Q9ndOJ03n2un2EeQYLni2fRM5ZXVHswG3iXyoC2Zoo6IlGWulHmG7qmOegSY9WdxbSKzRmXvIB
cswBwvgmHGhfGD5N2dye69cY/BLLFwd/FQJL1PvPt6PsanAGZSHTMKF1VqNv16rMQ6FYJ9N8KHjw
3Ol1C94wIpFUlIX9qxhqqPcHEInB37ZzCyywpVWq99s4fExCKF0oumsos66Vy/B5z5/iLsmvAAPM
mcFhgT+bQxbn2CwXGk6L176OMuObcfrjOoEWtfZG0pAI1SupOSg0lgAOjiqS2j6oiDJw8WIduQgF
C6GXT/Qz65ZmHGh8ag6lbkSjb2FJpWnvFL3EyaVzfZq0R3MoUTABeJCnndCOmDb/QtrJTgYQnJtp
bsXTYv83EkuFr1DZsQxpuHJyb+Pyx2KMn0VMUEFCJUn8k3jOTxfpIMfBfZAqk3RImEu1TK3FCqYr
gNZl1QelEZzIoKEWWwHKXIpx7oxqLK4sPVYmk3p9Ni7gKWdaB8xBUDm+p8SYFjMNhOhvbDatZUOe
rxMq2kirM4gL/U6APkdw9VbdcqIObFeN/C7uSo/p5DY7fUKSQslSOuMCOVvf2dzmI0LEpUIRDhr0
OXhqT+fz6EPIIkidUWIJVf26IPHzAQjBEgeqr9dEgKQpKbWRtX7a/Xb0s1LgZ8lj1j7R4/6EUh8A
JupJbYGqQ0go5sMqDZV9XvfxleJwafRWVR8sqpn8PshoxbczrcpgJZ8jvFeDJYDXuo5Afos/Mt8w
xXat3gHS+klRj3Y/J5qZ1/NaMHOfkDAPa3HpXC0apzFWDjUPoRSg0kuYB03KPc14jxo1qe44DhbI
/XVPsrpUQXURuiLAGW7guZAVtRnhhmxDSOcuvYKH9bCNrbeAER+xf5XksfBBgHjCgcVyYp3uTMhe
SnOGW6XYCiL+c+adxBytpiaMMuTs8Js03jVrYRKRIQx6jYEvCrIDpbHOxLhz/zaGFZK4zTPeJgWF
h1nPVJbp5VliKkwAdJA5bVnagy6QhcXMsZkk9JGheEhurHTL+trBHSo3KW1DiMeRCypRojOnMtcm
DPlmlESnKjIDcoOC7liV0r15LYvIJxd/g8WQ6i6mtWV1KbPKj9QR81gxQwkhmvLWUoB7Yf4Ngkwv
zzMCEXtxu1URF9hwENWRUY5PkWKF2btzb/tj1nTrDKL1XNx4H/isalAm0WfuJkn2Yn0to5uvQNkZ
2cma+AiHK6IYu8k6ao8O6HOL1TWm8ZIGxqqruxlT9a1CcUUQu9IQts05d/77QC38ZQzCdOsEDXIq
7dQf/MSYD0cFwQefhQFJ+yCoX27OPvTAFP6RISG+GKr/FglOtpgsnOW+S/eWx7G3G0cMbg5ZlzKk
ctv9BsGt4NKHRCdih8z3eBMBBxt1pYwHxdX/Fs4YT1YqOuumjMJVuznsrMCCBFQTcN1tcYvcWDGq
GM9QFNBeHZPyahZfFIL3A8ZYM3yoH1f8CvbvYCIwLAce0BYn7/LWk6kKj6v9VuYYnerecX4N0R5v
vt3XmbRtOpm52Nn2pXgZNC55Ytb6E0DQ1WbrR1JpaqIeimuGYyBN8M/W6Cf+45aXImb6tnRcNKun
uh9Brl2tiIhJdniPsGXynjqDCVj1CAs2utCDkDpGOp8iRR7G8BvAJTn84/MQxXamO3ANyuKpfx4x
oVacl/BX5hzbqTc3v6bZ1NOPKz2dA4aPiNb5C3FQq0Hby63YwIWXaRQIF+xlAmW5PKKKh0md2uyS
LpEP9ZpVMnJvo6yt08PdB1xOaLQ/xrqFzgRjARRQyaFHYyEW67FilP/SL2wqxsdrNcbAGkhmxDfI
JSQOQGyFghfNY/9l1Um3vqRpuEWM2mNj4M7soiBjEpxUtXqcj8Lx+DGQtx8UQCT2rv2aX0VbPCaB
2ckpfosMShmUgRKkCsIKn1bTC7m2Ev40lNimTvnLQzaDupaxwQbagc2DiWpv/0J9vvz0WHb+1wuU
QjX1eDJs1NspM1+dvGMnI3GrwZwetnFqgBaAjt3ON8Yy2Jy21gYLx6WKcjoobTMZrOlhmhOnSt4O
qb8lDiLmdzRISLCx0mn0fdywLjAVTCQQi4A9FX/uwCBbD01Oc9DqXha4bdsV7RHURAAF8y25DJCn
ed5rJ7f+05W18hOhJx0JsKJr5kZ6jf4OpNayQbMfFmRtt3SGpTBHAWqgQaoSGqmJH1+IeSIi65cd
EJLW17+85j9Nmxfxtck7J6zuyp88lbbIQFuU/UN7IHZ1fgT6pWMq2BwobtfAqzVfyalqSprUWHwR
dBLnVL8huXIA38CEcFps6KztY3PTXL6FDtmzTRigQT1BoVpLX9kCo4lnRAZST3YD+LXmOwadJEc8
9Rq6eJJNiJnW7vvo6NGEBTAnma4vHOv4LqRea+fw5ZZF8u0dd3lIAgyJ1MMtIpQbYcoc668yd7Sy
LtrsVUpyZRtsTHKEreRCXQvnGzd7si+bBtjxpFp/Kp2ACOA/0wx2kdqfRitZAkGi3DQfM/87CPET
JSkEm7TDufXZpfMjlTmYwIXyW0+ooM+P+nqySjfu1VRbccoF1NGYXZdEqYD+oIYqim1uV26ed8da
/9hKIOtN0csgtZ4znF0Up2bUscXpppkpe1naI/6QUUqUV3ZxzDfw67Pbny1bU1UcFJfU6E2NgGz9
ijLd1vIe2QagZMzI3wP2v2BNQwmcYBRn/ZYIO2xV58Re0LkUJLnJfNV2TTSHeu5BiqeNxskcGzw1
yeqi41NUcuxsdVvZQhnx4pflYcLmROPbSitf/HVAdF4P8ElBA6l+9aPAPi+X/Cpi98L0AKUR5+Jf
xyfXW0Gzr6XI+4AigRJJvyWTOxO2opko7/d2UrVA13EZN5L6eCqCc9QPm93Yx5RyhsMU5Vxp9eMs
HtD0eG3/fuj4Xw/s5jmIENeBwRUZ04nr30X/zYs2KMF3XW6YmJSkLtq5+ElV84/UX8tGEXbFrfwy
BDrlXUPUhRRC9kAKMZDCZzLGsmLKAezaGKe6DZGIx9tLytY3AxHeW5dCvfzlyoMj7e8q5g0Ecvz2
MhgoGqTm9LPCRpF1tD2yNQ6kHngvumQ9Xyj7rs2ydH2ohsAUjuhlCbEBIxtvM3g1hazoH4+JUG0I
oTyBh5QdzwI7W+/wJnr/ddDOB2P4K5IE0z+Av3dAbiQecTaISAwcRoF7nqVBcsp8lZ9SqtSwuPIZ
QQCG/uSEXUh3C0gW+fURMEgRwFJ23r899oxLwmz3xFRzACPMPeWWAGEstEtp5kvkSJoNKaMjzFhK
cTDuAnUwNtP+BtvgEv0GT1ZCTxSWNOJGQ3LIg/SQJl1h+bWIq9ea4m5e0NGrehuV/uOqq1CH8XvD
jQn0fPyR+8JrUYJmxiKeoUdDaMjitF8S7k24nrfNSpQJjprMi2hKiai4bmxino9Iv4e+CGuY7iNF
yQO3JvDjvuaHIQff7dVNrbFEYrMBpa6L4OvC5k8WRxRfJ6LGli4t8JLqF6J6r90Ke++220KBrZ1X
Dn5r9v/Tj8oowl+331kpr0QuJ4bYMoYd4C1XGvhVCgFkx2nGNFZ8ZBsZzOOvlziccMaSQxmCDERR
8POZYyNFqJnOEUd52cSLpnitxhCjfT71THKbgzeuGjk7JXVhWKgPBx68WiDvdme+xoqmnhO8Mk/H
FGjBifFIRi/G4LYHEBe+KIYbFwpshfEO+K13EhxOJcexy8A+Zytd0jg72SiXYyiBmS+q40AF5Z+v
WL7/2nD04vID9i0tzjmZpvde6NuFghWDvkY69RXqBmbCph2MGY85cdBPC0UaXnOGSkpqDlDIpX6J
g4APTI843T7YxnOQVgGB27FPm1cb3X4Ym7jfFkHZActHLRAK4T/039+JvNhgH5BwACTzMNWA1oGy
L+1OktNL6XAztH6ltkMi9igaxpUDontxpLTfMz4rvGDjUovU8ZL92lZ4G9F/pukuEuNFLcAFBxCX
PbXDyrcVbAp4C76214LBpwLZHaVPplcz4WSf4Teal2m2yrZDtB4LUo5rTLJpSGBq9mKJQ2tHkFBZ
4qwakFDnKZSKC8MXcdyCKJujlPjj/m7+C5dkpApeyRyD7x/28WK+Iu8uHdlfQLT9Qf5GvI2GXT7l
VYdUpNWYW0c8YyMy5NnBdldOczk5NiwX4TeCy4R93YpIMJIdarqxQR6GTtlS692Hl1h52DA+vSAH
7q2/PJC4l4OGY7PxS7ZXxgXpAAGM/Pq0wl0aTpRfIxJDUoEm2KXMdjchssgRIzso1FRa2ju46xqo
z4qZeZMG8mBNEoKyGc6/g7tgliHlyAaO6SKcECRRsuI8ie79BEtxuP0FQAtH05CRXQSuyJzT2NRg
+Xt/CbFuKomFFALRsF0Cmrx8Pxtw3Gg2ywLdkpLU4bLkVI6apGExAbSx4zfOGM00IRaSXVb8Q2WY
VhkhubcsUaOmEa2l0rXgAry/39iY0T/eh5ssWtCkrP7cU9GAg7w3T2heJciHYVhe4YVd4NH1Tn3h
jI7nzOLKBaALnwx3rxqWbcOZvqdOkwGeUXPKgxvpfV9glZ8PAuAszOa5UcG3ff4FX5KtpnTi9aBy
j5hhBKkiZXdJmJDvd0PKcEr3VSQ9WzIjrhTVIWnZZ+/L7E215zgKW/JYVhsZd44Jfngb7Zc8PPDR
SoT3GZxlvz8F/meMKRy9uPgTUvzMwuV6UPKJZAUQXF/4sByvNg/iWZyZ1ztRIgzuQzIPcU3ryebj
JlcVa2zNxwVb7daK4GEMqFWjFCqaXudWQn/duc5FT64pptE603J0oikOLFrPHR7Jh1TTxlTtIGyw
yOYTfOLouclQyyc5C3AezLMm6VatmaQoDMkU09NASo3omwKQWF8tkAPFwQUY7ZrHwxOh54x6pIyw
OwU9TD1wwDiWi6enYFIE0icXnVcUVGpeC9ICbaGFc6zZ4ntwwYhqDkPgLFLsRP7cRpvv+6CCb2ap
7PdElExGZS3bHJjm8Uu8w2BDVCTQvg8jYsUaeCgTt32cT07IyltxaBR9W7Y1zRUPXCWV5sqRO3eX
tfEQsk+T+7XEIbCRZWT7rnyAczL2aWEHoBV+rXKwis465p9zYrfH0u9QMQ+E+cKkaXko7cpcn/of
iSYyL3tCBE6FSa9DROFznLBM18/jzvOCwNcErkv+nBgQAbqxftg/8LpjT8lxV87dlDsSJr26ri18
kCQ6iRgsKavEANcTEoRS4RWcDr7keba318sknWhIkRPaDdTAC2ISh2mBdtsJ7ewNi6rzXawO5b+Y
aG8lihb610LVqrhGentFbZ9DoOmvN+iZauTwSEL5YozNRFV0pVsHoHJAy7s7O7nqFKJM+6kupdR6
Lr1ykyJunZg1z31UqK8rgT8Ea6iETyD8U2ImX6iYWIpKJbNS97yMjtOnjUXZSTLBruaelfLpqWhe
lwcpxpgbCH2G+VtxBQXacwRzZlpe/J4jJO6YMRJFaGZDO4lw6TlhWAqYF8bj0rMgUOQINNMc5Kty
knx8ICkAuNlFC8TS/7Da65BeeHgbh7+WDngFioNdorORbw7a71WYFZeTkNitaZx/DWk26EnLW2Be
WAiCviKD+HJo4n6VdtnSvZwvqvYjBCi0cH2DU2TlfvWgwWnNcQy0I6ByRvtsIR8aZdnRKQUfvjrV
pejRS8UZ3TQZqfMGI31cCakT30ZIdu0+jiNyZzjhHYyWJA9NhBkzkubEA9DQT9Y9Ts1BhlihX+UA
1y+OWtE/RFjXZzlxUDwURosoLsOjwADd65DH+O5LbFNLzB7sZ4oTu1F5SJhOIvPlhwjpirb+xe0Y
xy53C1MmI9MFwmHOa5hLTzQPAKoGU0VggR0gI9Zei1ZwnfSWQ35aRmZPQQatdS2hGDeCpg5UOEDc
8ptFL9jgeXUn7jJqrkLCtnOaZfygqPSXzuz1tQzgfwVgW65i3n8ZUyNBzD0y67aZIoMXsQG0jA7Z
decsTIwnv1tee8DUqzjwQQsGzba/NirRWP/1XE3GlaWLxnhZAf6lQh/iYg/sEaq0s4xOJAgihhW4
GYE2VxF3qHMCyCigsRbqCSGlS9Ve3XCNq4fCetL25HjU7xU+F5mTyLYvutskMwXrMcIPTagm4p3g
1NnBc7jx9+O4J+c1uzhk9jXu8aabbGGi+1pPMb1jKdgA43dcqZoSeXR9bUPJny1sawGv3rNqj/uD
Rbh19DwByDpvJinOfQy/H98UzzLE9kiKLwGFm+UzN7bRYS1MC6UopM7uSDSEVxc318SRXhgutaGv
Q4P0WJkaS5Or39OiX4f/NQ4YHR4YgDJ5ONGTiZTJVt+Ni/WxiMSXM5SxbPPbxIhSQygM4AaXdGvn
6Y1heAJ5SoYTdTT7w/e7x48DRH87m3eCJn4KTy2fqxF/E6plfTH5mKQ4kYTwl8JSkYZpV0bH06h6
tYAdolLWiV2drrysXo2nlzfQZTi/sSXClN4uC7C9FgWfEE4D47twK6lCmcFCxEtX8U46u0WGd3s+
pgeigkfBWsuHnBMBH0bHOKu51GtrYMhcNnCMRIvFDEogxEXXJ7IRBk5DmrgRwwUH2KWHohrBfm26
WKitzNsTSkK7SNzhd1SHrd0hCS80OPq319MNBxOrTUST1knaIzn9L3YnOYDjT19Y84CnFpRIamdH
N+Z3ixaM+kpbL68IqzyMbSSIueRKbL8vqRpOyHDVMmvWC8+hyI2/Aigphbnwix9XSPaqZBhOtM0N
qWs8XNCkyDh4EjhXgnn6LjjVu/HVPk0jgMsyOIbA6z8jn0h6U5CV3gRyS3xH2O2LCx6TbXa+Abyn
h4QQnkjSWD6KN/to8OFWYVsqUxApxe/FmgJ9JIEh6GGO2q7sbkve1wwu9E5br/QbhKQWav9L+BRr
CsiYgbZdFU4vl+8J+kAphc3uMx5qesK7h4qgHU2fUZNmU7xWqEKANqffsLQEuxEWm0+Slmltl1Ao
98f7U+DacytRmW8Rm09YInnyW+Ao1iElnrrhyrqm7LrS5fgNqH0EpSz4MoH/7kh5KZp6op5i03yg
MWb1iZnGbxL0BxkJDrMGL+mQjEnTdOk9y6AlBD6jrEuucC/S8hBWGETFAsx4g8vbuwwDaXXyiuZN
iFhES9YcMzE3EtjCSc7ZUOpFeREJvUtD5JeImCMyKJPbR3UCyBp+5aCsvwdFmiYyYVDcj50NkelM
NocpvVOIH8yiw7mzN37hAEA+ioZdcP9DPC7uLxzJ22lmuVm/ioWW8wHt8oeO9maJOhFf6xQo/gGs
IbL7EpXpYQONdP0MvMrjMaA8RgKD32VGGZrtZtdL1FbtbOKpv4tDdkLdfXGTp0cgbu0fTCejbI00
uJvEv+R6cbm8MfkWOB2eG1kGKbp95T5rhtWUJYlTfnTevCWstqhITUjcdcbWtkUsNPWvKKwHlJ0N
Lfs2CdD60g7r/yh1UgQO3tkm3gYzl9EnaKLXKhXQ9p0EmoFW7NlpnFw3dRa/lIYKCDiH1NRtr7yG
Bithg6vrZOtfZIp2SvqcR5Z865lUsWhXO20S1q5u9G5n0pGl2CofQo7K4UZW4zP9JngQATn0g/NQ
KkrDXnSN4szzSeBr3u2T6t6wlCF1yYfShYCO03ytGp1sjyjJ2gzRLRFbq3w3tuEw7v7bp1EPPPm3
vxzwEnzlH8QeZmOHJWcy+UEdQxenYHtvQRG2N+TLQZvwFiWqGaKXIx1x/Trw1gQEWZ3sLDA0WFVO
rSfMvpJVDD3sI9/6WLIJmJYLaIFId6vKoAxm2g+l3DB06BRev/sGczErroAFjs5RkjccqybeiPeB
ok+T8ztim6A7OHRCrRxsyNRNZp0ql7LToUWh6C2VCmNaZAvYsINYd/UjQsz5kCsK0E1LweHipYta
LVE82fIc83775tTVu+1v13LLgkxcJPbxRUd8gA69aUh/HIqy9Y0WvK2ZtrbmWx9tuytO/WOKTWgi
fIpJLNT3HWWepqfrnOUaAnroZcZ3alwn/yDuKDVO6Lp1wp1pLReGUl1A4QK784gzAogTDsdW5MlJ
aAWouZ7Bi/x8dCmV8BGWQemVMiGkQ0Vn2Jw8boRar4JBNz2SM3S393wThR2ZH+2qDONvfeHBmhn7
RKcOFxZmaU6ZhRlp5g9fqrbcAmBNOxM9FddVqkjYyuysDmlfVZN+32wN2zhJ9On05/LyKHG+c0xS
qm/20d/FQG/RNh6Ya4+WR4KbNTPC8ueNioR1AaibTO4bStsSYb/oK5VjIkuRbBN3Bh4zgZ8K9UZy
+uDtHjdkiLpPnLK9pj272nCEw48PluuhEkfd1Onr+DenaI9qN1ZyULaeC81IVCkKYv/aagvNkDbt
98qIbC96tmhOKbZCD8jKLQt/Rq6UZgfCmQW/PSPvRPhkgnZJd/a2u5Ta0c8ds4mS36t8wfKH3xaB
aOh59fmzWbBaykKcWU9agNRcbL8KOK6n3hBn2oWkOeTpJex971RCnBipevFpnvBYD8+/+JKgUVps
EPtvB0HtDkU0O5PX3+mkIDg20Gfgrtj8b2IkeHIs4WHt+C1ByOp7M9tUNFY8kUYEFOSubqhbmQq/
rc73CaGt/doLJicVbmvFKzHi2u5iNdUHKPmaPTTBbbfpxL6uEsj+AtIuLscAoDM//jdbfTfhqdAt
EkAUXCl7xdBhLTsWHVp8Mavsyl//pP6J9s+k+xHCcELKvancIwgSvgLdO3S9AjIelneA4GGbbSFY
yyL6vuATYEwaxdV+8jwifoQZSbySzwHCAt9XTfixPPlrYrLysggMTcW49jnVUvBdss66oRc4f6r7
6OblB+BCEzO3vO2I9Y+Hb/QruHXm0ObbjPrHuVnP37dNQvPA0A/Z/yA5R7RSctFzBt3DA7oWQ9E/
rAEHPUTw3SmPVFvF30fvzkqMgPs7JVE8bsc0o0ff/rsvf4x/3dzhW7DbjkSXuZI6a1KkOODwx0Ep
x7q6J527NlBP8OKI2FTE7I65kJT74zDtdGNqBQY0v0MteRSSWOgqvC5i876YlJMgBgWs3YHfwcBS
yq7Z2mlvoS/Dl/iuZUfUjozjcFcXMfM9HsdqVGKhxEhSWt72NXK7aDEDovBXjXozwBL/FSJJHCmL
D7PJ9Fujd1aofqmM9LmwgFGay5vajN9cl4HkX7VXbAj+wHUweLk9ILsdKycwClOCwcESb5q1Etz+
RWpioH9ie6yGOsurG1dVc7yC+iQTIV5IdPWGlMDyWAjxgPMQgIuV7Wn9a/a/i9HhPY3iJTb/BTwE
Rfr62T7Vonu6SMTAEU1zG1N3ZmyLJ34FFweweLb+LEnqKcLDfAorX+IZvLrLNB9H+Lw6RlGeI5p9
G2iTvs42Wrc8ZpMfnQdY7/8/YFw0KPOYFpSdlIidxRi3rS2Sf2JNyvT0Ajc2hgy+7FVSssC3mfYz
QI3iIvpMq74F6ZcO57RCPr75oCFG7ekjtnjsCFXb6h0k0K8rx5B2lJD4cbhlBuovwhJysmeoG60G
3o4MuDOioNTqp/IuuEyODGSoP/Sf4tJX7/ISnZnJBMxJwiFP9riACI9goZ9i0he3ro8otJrI90cP
3b5ObVyNB2EE44mgDhQbxx95YR1zC1gggwosBvLHX56HRIpi5uMR2hKjS3NZkzLw+IzMeNcKeCmS
wL/lWazCPogLpAxQclt76qCFRCKa9o3mrQXD0RmoPKEd0PPUT8lUEDhdv0nRz2v+I0CXHhBaJwld
+DafiykYJBXpoZhuoV/ALWk8hM9ss6LvNheZ80L3S2L1sXrndgjlA7NyG0hLXeJPWD+JZh5R9pC5
afMrQqjciWRfoQ+fG1pN8JxNZUCQZa6du4kQhy5TQ7/k3gN9RFSTsQW0Avah36LiLzuX6pGLkr5Z
k6tCPswzcZXEK81ej2UVq/f+QhruBeBkaHWNKYIIt2KYXO59n4hdzUHpZ+0P28XR40PlMr0NTR8+
rVkr/OmyR1bVNSaNy6OKcbg/u0aM5G0lGRaT7f6aGNqnRQC11Vp1mqjazZsNRnOW3fD1qO5ZTGg8
N7LmDbokaFm+L3csjad+mAMu8+iAW6FzGWum3dQCLOcDMIkXuhnJQZEnF7Tmjt9voNu4vQt0cUm4
KUW+5TbALPOKDHNw6u1eDu5Cdr0hniojjtpAO/vzzE+7VFlMu+1LGyuwujoUhA2LleuLQX7Q3zWs
xXXDHcwLNJtDzf40qVn5pD7PCyJTtIeZYwEEVEaWctw1l7NVTYKrZJO4aQ8hi6wYzbjzYEtWHBBS
JBwFN9G6phOMqWvJ6ptmvTD8sasHtcbyNlLxeo7a6sz2AqMYBb9mnms9QWhv/Eigevta421uJOVP
PFsbKmvbmZPkTahfVMP6AsUZv9QzPtFpZk/KktlWyAfrzDpMh8R6K9AF3vl/xevaoEXM+SgXNncS
8zhsg+OPL69Fa8nmKJFEiO7eaAASpoSxXLDNyXbOmNpFyxd8dIN17BqL+Cxc3plZudSJU3HjSmjR
gDpUJybbf/kpRoqT4uDgQqIW38t44C68oOJljLkf8JWi0HKbHzmiDJTLReRHCAz/U6gy/6i4kzFA
tTqXFGq5surYF9zvs86NKloOd+uSeul/XxfvjXKMZUK7SNR2oFK95CBu80Z+dsEOTyG28N96vLyN
t+dONeY3qOqkABScicx30mxFW/4VzDNQN/zoHU7S4PK60bUUyMDIxTmYt8FtBKwDPSsvlrE1Xafa
9Ey1qrvD/MUBaX8CwSUtJs4bcTMAFRz8pv8LWJxl0RC7dKcUJxjBs553EHWZyHhMuHJzt1sQzBwM
0cGiv8BUrVbJlpecQxYqCQW6D9992RuicX2njHfv0jIHDcJ3YfhwOXApxp8ogFXEvMkmnGn6Wekh
7cFErU0qytbcnouZprBycwGOXtwoU23j57rtAIjbfsicv26LG6vJcGEtnITK5vKJx1DoH9TPAFyr
1gQgU6TbAVIZPAkeh7NVlzLHPJNYKQ0LGr1TvHSfRKFXx16hjdv6/0lzkZ4QGoGyqrMC31ypjNU3
Ak5vvC56UUA66WWnkmYD2CjGCkhMobDHkG2xp0fwBzfvril81Cpjz7xF7Ic4t7Rso7GVKp1ERxpN
t0AWsradGwFu8h/IIgCPmcELh8gKVdSxLvF6Xxkk5+gKTCrOtJsAweedSNSUoPBzuEyyPhsiA/81
9X1XvD1Ka9AeXYrwlyzQnYGKLtSpH3LXrUbOij5n9LxeZ4jL+q0H3oNqDLUJ18YiAkY3GOx6xDNH
AB4J7sm83jAyB6oKXkiqBZGKC3nWfJyC2qcuNd6GO9RtwHpJWodiq+d7aTei7o5yVsJuDbF1X42f
vK8uooWY/6zk01iaIuht9xu0B41fhOOcU+SD6CYoX5NNBLLlzobTryXvTx2CYfAjIJNbrJhMYfEB
vUCzgvZYDzEavE0qnUUfDpd31MWkmAWUtrzvK+Tr3E/cFcI0U5otTbvdTMU4iF4C71zz7p61KzFH
K/24DmmfLLjumwfJIP2b2avUjOEH/xFCI1lCAxhpmuI4DMYy5hXcYUtrUqUKEDUu7ITFUiyXA+8h
UqPEY/YtA9ghoPjJ/Tf5jVZ+R6CxXgOcQfXCmhTukWxSCeipHq6CImf5jqt9M4lvizWfk1I0CwZa
fKrnJIT5qU2jpJTadTngRGjRbx2Fa4Oa3ftfqi3qYja5K/Z8DGVxMUPbX+iPM9T66eJemCtbOPkb
KSM8uGEEbdw1Uu+FTWIx7E1z9dsKR6MFLOR1FwaCwBuyoX1Dgox/C1xHiyeyM8DSi71wArOSOwNd
EwDIRE8BpNwA5F7yetLm+Dyw0TrIiu27ORlGGNzb9H6c2DPSIywWFhPkSfU9D1KFcqxoI57sos1D
C8iYwqRXNmkboZDPb2PILGAK7OdlqcPu6fh3tq4+qq4sL80jo/+Y4Lheq/ERQou8TcHf4y13f2mC
/5ESrf11rwPgCuLIukxsPICVw7WAfebq63Ggra+5fv4vi1Hn0klouBpVgHMfa1Of6SF8Mvn8Sh/d
KM5e5stdqshzXHyGPW1xVIqGBLHqWyRzIuCa5TuhMArR6xarxvsvkUAwvR4+UAYBlcueRX8y7YBN
ek67OsfZBSmWY2bkvm+U8YAogddRpdwAxlgPVlxaia9Ut9PgqQAhNqveVPOWuusjVJalh5Pp/jEO
3Cfh0BNOBq7sc58OiMbgrn3l15sXIcO7PEvnbgBNAHHZEgAlZ6r7fcrfKSP1v3/rXE9fAxJDXuvl
IwHNKqACrltrwxhN07CpWd6gDo9IQFq8sVP42BEfIdFgu3ylLHNIf9sDmY37j6zWsJsQVTEwqMoI
F0/gsibg6EG0jsPt1stgEFOU7WL2T/p1iu0LAe8Mm6Aj7i413nVwRc2LHwKg5JaOp8BGZLs9VPqI
bmMJWF8CpluXwtz+vYjJ10alzOnZeTA38JG5m1F4d09ZlcSaRWhP4EC8OkKqGAFcY1bQkwnBxoLp
8MNpcwP/zyGbuDkTzwV5YhC9nWDSjiSWwqMvL1PK/8AspSDBYZ693gaHpXbsFwKYdX4c+T0pLuPQ
T2YSmJu5xdfnFn+pJ0LexKuv26kaeuPWpycQ1i9ygkbcvQQ7RHfcyKViz6bK7aoce79BstSeeRvQ
9jRUEhNkk2uh1R6MPnetgEyYHf79SbyEB2wzVJ8c03yrbKN0X6m9ch4mhMdJ7uqnuf8iaHgyFNiK
HSyhqweMR4YFzHZDknw+AvmEtjD1OmUIbwI6xqPN52go+TyaETy40xupCTDfgVxKYcpJk37q4VKx
oPu7nhhu/7c3sCphYkNHFLlDOu2Pcnca3KX6sQDaftUn0DGW3e/zBMFEB0IxpKsb+3O3lc8hCzw6
zelRQuUQS9qgapop/FOCWOtPzKVU5+S/rguDVCQy4oJryiCzGCuzPO1v4nrO8WJZcKU17gMhKYaA
B4CMdoKkySo97h3gwXCyFYoB5AO5CDstFoiTNkdUDNgDz+3tLF3ybLy+r88PWfVdbUEaYJZCtcfE
JjwVI4B71wjPUcIfo0f1JRqvcjkdgjQ74EfFonYSfkIvaS9Hym38SLWva+3tmmB8srIiYOp73kVp
tP0d3X8HttvlpvWGQ6rGwS1PtXm9DrxY/sWg4Fv7CCWcV/yfKDRdZKGWUE6co5xE1GLoAp9JoRz/
V4T1v0MLWLUroanp9inSocQp3sjuvmrPyo/RD8mEcub88iE1CfO87Mp20/8W2BtSeJ8qnUMoVrF/
L9J+DDRnvyL14LthKpPkZTcp+lVq0CF+0MRxIjX/aKofGvPoxKBqT5bK+VeR6nOfdXLbmA01fmIh
fv3GCqiqgNCWRzkRBilzHKnFVe+3aOHq87FfNprsVx082QEHEpaO6LfuZARE0GHpQhsE/bR8n5OX
XiEv+AT62pmT+kR4T3WW0xJU6q0nhHV4/KacObpuNZUFd9XXdZ2rr6Avk5O4ciha7FsY6vXwEInw
D7MUw5+LXcVHA7kpul8/aMXUY0i1lUXYOkf86Dpw09+deTyDqHIbP0uPnlvVNP8Ljug75JPtZouO
uvgT5HuHzuldzQcMRCXZopMpZXAyY/k/c43ww13LEUtm597KfNz1qHj1HukFmpNob67kcRYmtZwi
gjenrmuJeettaC+6lPcUG9uI9VAg30gYpp16hdtA6kS0XY8nkoaK1wdAxtrJry+QM4sOT4seAp6F
8GTH7wsloEYrN6zoCFjxNtckynYrigT1gp6uqWCAmSEneXOIQ2o6SD30yKc+jtoDZI0jyUb+8dlb
YdbJ12lVDvkawkaOiBNr3uy5kif6xfgLd+rCvMz99aBVdjjpXVjJTCcYHA3dYIv835TNkgp8O56x
iO9oajsIVioaBdm1typbudzZkYLT6+dVito7JwEfFEP9+oGXakZHbn0suJRsjWa8avCk4KSvmeHm
LDqUYYVCSC9UGJqim5UDau5hLQmoeeM3OtumNkM4r55u1+ObJrXJseIBsAtFohXnHUFXW9yTMwBP
v82TUOoS9JqXzueSeQ8t948+v+Ptb8JlHRVrwc6lueoYaUHmofKi+kGiUcRAAXX3wab3hMfXxI0b
vLXmqzD7/R49Cec7hQ2bCZAqQKOIPhJEcKLrDdNhuXaKWPHDiV+gy377S8XQqnE7QOcELc/utADi
mz+v+8hqJyRdaDEMYDqkiZzBLRGME6CKVQQ3aV7FrCVWsNwhcThqcl3NelmwASl853ZV76ONnX6m
3acBqmFiVizBxPNH6JEsTZ52k/SLY2p1NkNNf0UkSTspbaWlWcFbzIwF/2ddAm5c2HQWIme2GkHW
e1g/pFrEhvitFBv0AQ1SnFLxEhErowowAKyriGTEMpFbjnqaYw/R7eQSpZnPj8y/fEIT0pkNutip
709a7mJmRARMcIGUoTgz726UVlfNVZ8CYeRVLGXpzJumpwfa5gqSKnCeXPNcGudI2il2fhMcv9Wd
d0zqhQI9hXG+UNdNKvBcfhgvq/3Ae/abQame7nEWRIrbXsOgmKXqC1+zf9azNIqW5yu9LBM6JM0H
dXA6m5FAnJwm0j6Tw/dku/PIGbgLKp4JMXVfnxadjM6pSxra/QNce7bGaBOeGAizEULzFIQhE+xv
ula92cTDVsU7HbRg1l7toQMEfZ2LtdXE7BcIPCnuRRDHbKkebxTvhyeuIqa69mSrltlE0yyFQX0b
Y381KI8kQz28KclkKVl//J/XbvviP6AoagmI/zOX248rHXSE9FZ3OjGqgpGG1t1iib9FZ00yF4O6
p5nyD/GTuFPWEyHZ8oZm0odEAdeEOI2FJGM8VaGx022s6AyhpZlVsWOcBDngTXtVxWD8U0G5idOB
gA+pBihSTqmd75m2+XWxrL+3VOyQun11rzDOKCLXWEW6i6PbcQBopTeJioQIMRTnxE+/i+RVmn6q
rSd5x1tAiSzR57D4WlM2vOBY7XKIkWAH40mrmZaeMsYusfhM+2/PyX7y7yEJqRpbjYecJ24CqeQl
DaaiJfXLfEOgC8G9kQt9enzhUIR1fvM49VmX9/LrWxQRvTlN9OXGSrdK2cT3WwrSXLBbMnSW8Q1F
qYJ/aR6eVfnddxHI5CgXlHjrJC1j9OKtKZiYUJbxPom2T2FHgH1C7fSQjns+DdpWN0c5qGiav8O+
gn1Vk3DGgQr3WzonhKgjM4duGk76xqQNwQ8a3tvMt/EEEPL6/6mKynLAP3033xLxUW8znhMmciGp
ylj1IB601rNe5Enc7LwA28lJYJ5C0E6+Qoyx3AiHUPDh+m8v+5enmkk5WN8uBlyTTBf6RPEU5Z86
P7u2NnklN0jD1yDDHehsZHQMj/P3dtrcmOG8nX/IAf4nJnVvZES1UGaWq+tM4r9+YeLHRZw30LMk
C7P4ki5R1mf0I5YBp0d31QU0VLF1earcorcBNLW0A2sYX8N7kbxggwzOei0locjXgbKQNOcNqJBS
dH/EMeZIyqY8VjuI7OAvuGZZneTkIHU7HhoQiYD7DpUtxionrj59PPvkLjn0D9cc00+3R66OZur/
BihB2eVAIUGASfqDQ8XZRoz+9yToYf4jI3RRqGaTRYtoUkIMruiBZPAy9jlapkovhrHBIwGd87u8
7M9McZA8Pfq9e0fpFcFq/2GcNIXRpKN+2aC/QHFN/0GU786JQ/pouhr1smJj0wxTsKVZuk9mzTzc
r3PiEUfoS2mZYpXh38lwjpFxyMXtNt1t5fliafW/Q7Q5nKSZG2wj14oHmrNvFbs6O2sjD0kZN7yB
IXVQ0bX2Iat9/wHRopjq3FcGQ2X6Jd+fv30fYWyEapLL11+NmdkQQ9gwfvCp2G+MQuZRilfxSPPu
eG3IZBM2bqfQYsCcLZdNYeYQQMHPSCW9s3gjRO9TMbErGQl93ZDcSIo6P+3R8PG17i7hEiKtkNHZ
YN+gr1q2GG8YIcdrRrFkRRRpuWoZW0MuBMQpgu5q9PYH7SGRn9ykNKVGam4DsbisaqsW0p96ZBhH
ute9v8XfC/lFqs34KaLVzlK/c6ofll6Nv71o2jRKDXutBlYjh9ahz6FDstDHb83T0g3Dl8fB5FLL
XyJEUigPSUmVjrCRbx9dj6p+BLkAIkhNeeSpK9hPw0lo6tkzlq5lzVRh2E290b5drJDQ8I1nA/Id
3bSsZOEfJPcAOVQYvJUHqyLmIyan8aGDidHj5JsRqYUBg4SwgYeoPFrADmGcu4TNefa4Lb6xe8zB
2cvR2EduleQl903e5hWPdmyNsvxLU4yvdBuRaM/pj8pRyYNu68ifBAIndN7YzN+7DqJIesGTGTic
y/aDFZnoKMnkyrkUf/97H5jEsUfosRqGjsXcbiXedyVjj2TWXxY1bcSJgO+AbZgmgaw6I9gHQyNk
feti9V5j/3ytLWTYOxts02AfyEmiYTMCIDlXYVxvJO5BWJmzPMeq2dZ7hXPuGSgnAuLjWBwhonbi
4O9uVSbtPNKtIXx7FbrO6o+tah6vc+Tr3hkuhWFVv7q/XUEgkzfc9ztzpwgUVMlocs2EKMGPN87C
NcBSK/IqQ6qxzS4Jyk8tzvRCfs/PGSUWpB82IAPWV0MSEhjKECH2ojowhjPDK57hjYEnx4GFrfDm
RM8K0LHCzIxAPI7XJhOH5pQo+b8tqRpBI2O6lhWeke22e7djLQVDWokL0Gr4UiwvzCvnr5l4Rv8D
GWv0fxyQBDhsG+qAX215JWEpOel6UI0Hh1/eYKukD6Vwk8PKymmhCpK5IFoSJ8clt6B7ds6eecQ5
cKtpSx340PWUvZtCnuGMITlk14FPTuw1dITRY1AlK20kbFKhgQ5wqKEoCApty5OnxNCeyqQkjnuD
WZ2e5MFetyrKWHv7wQY7tlSJqTvU2X4baCQ5OgJEGtwd0KASvPX6HvhVS8y/Ie02Hs0Qdi5BYksh
tTzqory5d3u1HKwN1rZsUYU1vQr3WX6pLHH51v9kPc9pYYaKMC1mgroQu0CvtKeoEO5YWCislQi8
31DykcKz1g9kAUmmeY+epAnGxFzD2UVwcTol1kN8BY8+P9LwHUrCYDrXMBdVreJtmlGWhNx21T7x
r5hIJfFRyiMWvp4+HDidiBCdiUvME0B1NCsX1vrSQub4gZhqR3Yll8mwnyWW5PcFYfOT0xnpV/i3
iTJuq6SHibv4SyAZbC5Y+3apH/dhdisoqMA/qdRivDelApqGEAAV72yTZqehoX+HtgzGvEJM+KX8
iTdQp567GGg/Se0zvimaN7PAQ/0xCz34S4LBtopfxrqzPn2gmCy73jFwyhATTMCxQz/1qsb2vXCS
8P+XkkkmMPn2gzQgmJNKCP09vgPWKEKn6lt2voMwaILEm4AXHnHuuyECfxsdq7eBSdjn1+XA/6w6
HDmKqSkoSPpVlZBumgjwQvePvUgyp8/VR3gd5ObG6dmdhCIWyeu0LkrMiwIDvsCVhyyvZeVFqIbe
4vsTXsB5UImq6KFal2g9RpZ5082ZTmTWzDyz5dTxLGsqGit7Xr/NYWVTzLKCg7Y2InEqMpTQ/DPN
cg2cXKRyTFiRpx0HGHM4IccVMhLuTVUFv7/4HxO5TwEC2VD6snxU+Lu1REcS+HI6/xlAdTtj/REb
TrH+sLiA/TrDjxmgaMgCw1UYFhzCerXua21VrCcleIcoprXsY+uXr22NgxU0R8ZZn/YlwwabJ/be
ZN38MpX7XOlxz0DEbb2w7gDRGw+qWFx06mjSCRRxxCPp2BfdlBxJhJ+QCbLOc3Ob7siVm/8GyVzU
zIweywsc0Wbbu1pWV5r2D3mFMvXHGtZa49XShCFcF2eZdQwhns2NXkLlIqKabjkEpJTExNr4J2bu
Y0bPk396OGk84ZcUCvBeM4sQeZzVrVbSyJjj/73IjLqkqVpTcSVsugYzWAlTAYwXAF1uwT3Wx2nu
lN/WVdu+S5N/wuctV8Rf+xIfFA5SPBQ4Vc69OFV3YB+P6eJNOIllFfWKg5IV7V+mCoH1xXNxlIQC
AhRrplkeC0A4s98aYKBJh1fEa7qqwMTl/pZxJ+KpMqomZFkTejvjBDo5AA5bA96Dwj1Hyph2JgG0
VaWeYkZXMNUb/i5g9OsqaLs7a4fZwhz7gepcyD387nN1azDXlex/Vl9QIx2tDHIPWjNbmlissijk
iH+gtJx5SdZLQ77PHN0bIDSArcP0bPW8MKSfz22LEjlNaTujXa3b0S4kjhUFibux7alRNx4FVxPN
fKeFdDC/foJWRMCBzQ84W473hErdxLvXK8Z7JE8+SwHWGGaWwOO5TnKozMKcm7td9dDXmABVQTpm
hLLtHaXfhrRXBxkyS5muOhn3r8DHtSG12HfEsLc9s8L9xMKIHWPKkQBJBKCHoZOQkI4cobxIYag4
B49UTbhi7/1j6Rvfial7qhrIBGNnATy9WqZZsp9qGRTJkl0B/uqvvIyhRbZI6+71nNUtimR5OibT
tIfkB4RIm2wbdPXiu0JUKw18BWnQwOwJUHxAnT3qAJRvBBKQDkEAGoIGkjLKD2ozGNIs8kb0orSm
fDNl90qL3H2BR9Kx3NrJHzskQGsFOhq/1zN8XDG2FXxsu4DrqO79lcAX0qSmIzUB+aicDGh2IutJ
g7uadwKFT1e+tfbjY+tOviaxsPi1TanwzL1KJCyVejp10Ic4D8gyxHfUP7yTxgmD/pOdvLN/6ENp
mQ1w0Ca2jGTIAEJ3MvNaCXd0FXwK4l459Zvv2yHPOBxFyQTwor8wiPIVeWntzDsia+IJxjii6AY+
lzROV3RfQr9tFJyvmair5yqXto4RjQQeuxov65ZEzlG65YqHE4rHsmyXPBnf3tgB+LLGHTR4RXJQ
Xe0Bs7hciRjCuP+UyPeO/ffWd4QS5HjqYtDyesktU1M0OH1BeeelTxbllGnJUZvMYTUsTHymPr7f
8KvtZXO5gthRzEkNovClz6sZfJh/xERpJ16G2EcOBZJEmHRrTSskw0Y1poSqu19Tk3OyM/nvj7Ns
in0L0D2uxX89QBn5MAXlafL/y/RposRkZnUh9YhnLjXZKnb3aBHRJp+v4SJk1fuTTKpSQezLlA/v
8xErDlwzuKGUXm68L6DlfRHuxnXbQyS6OIAgm57v6CPFX9JgPWxteBZp+1ERQi39YMwqIx7XXr3H
YtpLblGu56bKfw4zw4/pvdbmUcPgF4dqneWxfCOUpIPhXtI5Xaeb5hHuoCWmBKcaF+k+oijcRTN7
GioSLOrVy+BqqvmdCdFIJ3SC3QiKrniEozJisPN3TKO8C/+MaTgotDrLN69PNaG0ORanqV649Vwi
Nco8XK1TXo+A2nUtEG++u5Oo8GVegSyUku1ugiHuJUMnieJCiEkLGjTiOUBRD+G9ldrAr1yl8b24
mOfV5Gfn59YA/H6MRWLKZDWW4PnAP2xhYnBnY5X6Ox/Muo5aOyQVGz1BbZrCemxXI6Jd9q7bnS05
5gkbrOH5aXRJS31zdr18dhGvaCR6jrL+E40a/B893iv12x7kXtBd2WdxhOfQSrrrroTyDWUYEv4s
2pmDKU2xnUgFJtQIoaoEOpwyXfMhoKx/pprihgqM0NGXU+xWETFTKvYT4Yz4xavRtGyvkgAnE3cC
mxNG07Iug6TbdKpohC8q6POX1qaoMjOBFc0Du+D7oFCTAj6pKoy3oZ56q0Xtzts5GTCvvCEVA19M
Bu4wdU+XiWBO3wuN2yl3K4RxWcLeunYwh/DLB1rHlVy9dIAVJn3npF8hl0M8gqMGIdS/CRA4U1cG
03TosSZCVeSSs0Fnz8Klx5DBkUX4Qk8pi9hv5XQJIjxruImxuOlLUQ2O5bzQwA0VOBldZqsVWqx8
gYdZ35/SuPB956IUp44tIiokwoNB8Yx941uz+FS2aqxBGlGusJHgWnxFSaDr5OJow/C3N+NvL11p
JgoSniBAYWOhj++aeP2avkqBay2Sy8xPFClVhlXZ3BDvSTptRaAkWclb/f5xpx7AypASJRN4A3mc
Z9m1SZ5Je08S09a1mEXnZHKQX+7SsKTTo7l0GFLrZ4AiR2fmoJ73n/Qh84D1E18mjswkPpfthHzI
wIdUesFTxTI2WFej+yPbdU0a4FNlnrI5vhPXrppP6DWSjuW5IOMNYf+sRHh0IZ1yylJw0CWGM6dx
Zs6LCYEq7EmYYHhetl+5pK9HcAO6x4y2UQH8XHRruis8U9gZpHkrdFe70i7HbX2+hZF6sTQQXRm9
NMbu0FPakwqWxA6O8j4gsiz/pJem2+/6nFMHTdDv6KkgR1GcQwvK9iOBdZRdRMsL9SYzxRkFBmf6
fWnPXhJKDpmIfd0iSZJPR3tF843j8TFR41qWdj7M+JMetP1DKMDA6ZRKC2Y0zIJFJ6g0wON2mXKr
vy9rs4oc8jVUjFjmviTIyZl0YX2ilbKwVfbvMcBH27vjGoBgJINZ/4pHnMaICiESJkgz9D1qGeGq
QLUobqLWy5/SX6h+ckWZ9J752rZI71tKGKSC8/P3VT4gzFjVZqOBA6S3uDC9I+MeGaSuCtazBdgu
SMmZhGtq5hM0J7kzPJjEEhaku//4W8htchPpxI7WbcRsn2WLL1lg56FRLb58K9uXeLq8OEy9XsSw
R57XC5pVq/pLv2i80A1RitQBlRwCXIE/TCegoVtpEXIFLI2uEUwB8l1e6hSj8/MYYBa6qLYeInA7
iz+bq8icf1Grb984GGkQsb2LTIYUt6pd6cPpzsCI4of4DDOKDClVFONR4I1DbA9y2ZUgoK1y4utE
tMOuLOMnwz28OYih704tjxfYQk6j/d0NtagRRJ4EVOqPIhJ+dzUaVKIf9d7w21QcNBpp1Pv0afxE
Lqn72AlSga9+84+TnvM/rI/bhVNtsSniZ7oxGUkbuV8c4kUMEX5qd1AfMS5fHxSfv3DjsM9PbZQ+
PFveAVypF8FnmXyRsyTT9sVFl1X8pNhqqIfRhubXxt82iFQu0cfOXULqlyt1CJH23kFISrAZDH8g
WJR8pUqFhV0syk570ROD5+pljNUAMkC9ciW5pG8z8ByrentRtRDuJwoGJDrDw+JhuCrShRRy7SCd
/r3jXxBLHrSHMkYbb2ESAIpCvu6OgSRs3R5Z8T5OxT//wGf88yPwGnA0D1v7aI2rWxOV6NH+aOfI
4YlH5lcv/0al/etd7m/jvuF6vAA7RUcJg0Rv1RoUfb6FrYFR/WVOaO2GLzH00wvJpPdzu7bjs5mg
SAX3jZT2clysgJrjKyxxlAInlOKn0V9lR/f2svBfHFGxybC3wdpBJ2P39UYZ9uQ2W86BaFisJVK7
AKOvGL9SCz0vkBfC2p8A5NBtG/WHPYseeQ/l3tD4HQHm0WWQpCTniUJ6sgOLbCSZIfk10ibvD/4v
q2fsNgdA8AoJXAYXAOZgpUN1GwS7tV2apC8wel7r+y40NjNL9BOPRcROpLCjme9bId2gAMZ0jypc
Se8EE4TvxgvO12QQK+s1R9syhqp1AhLI/Otle6KMPNg9ktEElGgCbT/CRKtC8Kuu0PLm2jeY2iLN
eI/nEHJ81CjCMkSW7WsSzHpmdOzlZ5ULJ1ertMdZ2MwL1dDOiJEnbGkJnAA9cqsHqwzr7CoLioQR
JW1slXjGhABHOCchzvPkOrYeuM59ZD+UjTsAz0vOnAKUxI11CurcBN63mnejDwZhNJ3TvWSkevkg
i2R4HjXqUnFy47eVixkcTkefuFYIgI4Lshp9dcLlQm1mVFtoFreHQHVlNdsFhVW5IETxZ90TRNe6
VrtkB7eznhdxxpS2dv9XrSuFjUbWKgC7h+2rbDta13ruRKywtdpdtzfTEM78VlnbM3OsrXySa27d
TEgKs8bcnxjS+LZwX0v5f1+RJf02GrI7ey2Jxd3uvGMxXQsvULasVoJ1j3zSBHvafI7D6z5R+Bo1
mxBnAuoDX75cC97CC08nwJXZ2hZeJUvfhPTU27Aa8tfzJzqdOlqqlvHE7lyOkEzjUqhuMUy2Ps34
W3tvTAkZpHkXZs7ijk+nDDvjqPK+rY0CJnWEQcpOjEBhBIi4ztFSLbI7oy7GqACxGZhWS3sbumx1
CiVmvO7cEcHb2o6zVui2ZlP10/jIF4bpVI7eMGofCVCr845juTxc8vIRCzRCjlA5/2d1Rh3sb7Sy
SDNY8kZwNmZfgi8mOlu3hj/5aL4FCb3WU0tES+jRFbajJNc40y3Bpf65mXqXvdBgZKhVLgJhECHQ
bW0cU+0UeD8GR+lujgkfEd9v9oUuh8/n92lFCP7fhiqCpOvCWr7nFVHtLVU9uOLbap3sdQXC0FhG
U4vA2xZscSu38/dPvBl8aBkepisKJWfHeLh4X418EYMl0baKrbPtE0TQm/p9PePK4BUwDBOQR9yW
HdnUEvrOVQOttkg8Dr36VRJxial0i5dmPXwYjji1DvPysxG65kMKsag4jPzM+2VLu9DkXM//bebY
vFb+kfW8MJq61hYi91pBLSXvDz7SYR3O5ur2OT2o0BpoAgw0GaCBnciyEwPfXeea97zmoqtAsKeC
HnUyRzhmkxPqRib9S7YwnMg4xaloOVYhJoVQepHqKpgN1oTFRCW1y71YhQ1qs+KgtuXk1vvplF2b
MEF4g3BdZY8PiR5C1o8Kh5ItNyAhs7NuSWqEFxNr49fLU6zg+GqfRvKZKOerfwWogoUcTFacZ2Ki
CDR1hyMeZTtiEnHTFg/B/C/5pDyl6MmRjS4HAY4W5kWEFG8jkR5Nuz0m+nkrJgBqKWwhtoQ0mO+u
oW61D3ZN+u/cJdUT/IL6nqz41D2JRsyc7DX7yOtp5dEwN1hACzvtpJDKRJHden4wdnNyMGvzZ0ve
TxmkFRa/7/KrMmzYdSeB6IBeKP1y+hwCKHvj4e08QJbO31XqIWD/sI/Rv3eaBHklnDrxp5Dp1006
KrnDeTJ6t7zShZEUgHWhUo3h1x9boerOa+cLF3T5o7BxPfHGLWrg9TTqDnuFY/njn7h55kOIhcsQ
qHHJqU0G6ujBWQLpyam/NPIuPs6j7s+domYtIQl1dGmglWhwiRZ5nME3Mc+FBukQitRlibCMu1+I
ZGaXPhQUmqUDvaeBYL0fEuHDNeQCWnRM7+Wks2W5oq6yAWd1+BHpstXx9S0qESZUgD/JBLkxgeGL
TLGpSOx78tZsmUtizUbIII3/k+yYz1Yjkp3Mww5xC16yHPsImlCk+FwMjdpSGlPsnos1WgazHGEH
/awDZpda/k3A/ixl4OVCIbtv8CFNTZvYIGUNNc50+c1agH0B8dY32yyYTMs1hPQfdVddUYtLXNjP
pIh3EU1NXSM9ahLjZBgScx3YPv5k0W8BRz5dNNYVuNMekK3tdu6AdEw36HYASNPWlNTnYdOmo8IB
P+vov4wGAfh+Z2KF6ih8ifXybSAfGIww+dHUD5CIk698+JUI6Ia48kfJVHEKZ6+QjZuj5KbEo8K0
1JxVoq22c0Tj5mHbMqYJ+NMEKzjZyg7Cum6vWbVuXw5UtH0GTamOtXNrvK6WB5cbPz3odKjqZpeE
oNfQvapnjckv2Of1uJAaiYct+mfRvFaARXIAfc9Nz3HAiCBESqxcjVHTzNJsGOGOGcMTDqPqf01C
E8y7lqtqLsv95jScJBi/eUK6rcXz+HzFnnmyrj8CjKB5FrFxlkGyYez7pEqVm5CjT/qxoSs2hzjp
IgxWQfDD3oLiuHs3gc3deGFhQpT2M6ZydYXlMdgiEVWLIT5YgbDgDTue0suOzBJseNVOwvXq78yb
NOBlIylx3QbingBfhW7cGqb2RloC1ABgy4YTYwJAlVZfRVLcAdt1BfZoL9tv1iR281BaO64FGPic
wt9gqjMUAmNGxnrHimaOAjqkSbXVaYB9Phz32TTklyY8+VnqH/tbZoZfKW51RvSVvq22McJN6JLZ
BHNoVqQNQefG25cEwN9QN0nCWJuJY4USYIfCIO70ildmA5kdoVHVaIwfNOLgYkE01ANDhvhpFFcd
Guoq7SDUvDOl2V2sfkqjPF9Y6Va2HBOA/LzvrYLO1+xZyt4ew2aXhDuYGaFLwcK5xQ+ngZGjz8iG
jzhteDKJENazhyJdYuCaczkXyi4ec0c3EkEaJrKBYunMROkmlQ7TZ38wetgx9DaQoDnfHFV/8noC
BOQj8KfmNHKvuG+VWcVn6iuyhmt4AaHr5lZnJXESWH9Bw2bassIT80PnzvMV4KK/fupZWZWmfigY
/+StjGn/7YzU2gXZBpRd6spyJBTs81ux9ry+gHrYEJvsaLsJJNM1nz/tK+aPZ+VO5EB34w8JHT22
2zLthGAABKJWT/Pjcgu3F4k9QiWTEsZ2CZJifHrLuBVgebmHU90+vOYy9F83JK8o8btjH4yIM8V7
RufyLf208H66VpDxLa+EhNtXQJwj4Kd4vdT5+XizO5BODw/+jBFuOkHc875z3/l/2GCHnzMvY7Vi
6mQzAP1jLgr87eptqaU6BShrj+NDan3G2G6cp18ZniYH9JllFrgUnlyWQ8/9Ac9jonLLcIaTTlV5
C7v8LeRKvctBPw9qjbItHBzsUC6fAGDCSvt3aTIle9UfleSbxM4yxBJGjS6CzRgHTVxtwwZOzPzz
gAqXvcGWgwtORAWV2YGmgXJDwlPH5FmRh7wOpLOxpq3ALszfC4HS+9xQlhNrwymJ0sobMURPBqx5
PET2bf+DHOlNCXEADiDp4CVviYuc3lqG+n3EgP8IJMi9dfREMUVLajznMAGGBSRLu2HC3OMyIZfb
Mj+gRMkMagJDeHYA9PnojAOdHoB+dA/UWXPVZMNfh4F7cjYjVRm+nJZUJS3NKxtw/HryFgXKXaN9
DOlFN9CQqDi6OqdJjY7FhoyhZ510FXQ67Vy1HENLzv8JotnA6dinJhgMXuMWHW/JUjre5Ln5DaLc
YGpHtA8AML+ROqFOW4NozLcP4BPQ8UNnAdsjIkTS3cwHStCAFoWhmsDXAYBh8kFDyv5TkqXA58iM
B2PhHnPSWAftPw/CZ6DtU8jBYC6pO74L0SQc+AZs5lOiQ3pBs77aM64oNsfJbCQRJ6V6C5X1pz2D
tPmqqn7N0KlyLeil6U4nt9zxs0S8ZbX24/2pjsvy5H8EGnoEqgRy5GxZqgDUoNiTaEa68SCrx3EN
LcklXwGSoIHJaFhkrs9L4TTBD53kg6CyAfi0ENdKRlQNY0dJYdxN6oJzIph9ubTmTcIr6BtuQc+x
+8xcOJrX0wPpFa/E+33+GOlx7fjuhyXr0pBfdivfPtouQFdPt2CoD6EGNU77zIcABl/w78Gk/yb9
5CLOGMs2pC7x26f5/e/HP8qlKYdUSkdG89Bye9eHumtSWLLbMhaZXYZrC+ZXH0ZB3Jf/79b7gse8
Wb572W974fr+JMVcGMpHvQqRC57AY4iFNwVMumegSk86dhMWeKfOD9HLpemwqiZkpkX4MtgLcL9T
7NOtZb714+9b8Sg0cGwBCsTqADe9elwJO8/Fi+2s2PFhcaCT7z4bno6MQYkdtwjMSW1PI8qEByc+
vmEFNb1xEsaeR9YIbpr0xPvm92nj5i2Trf4OnihUUgeUGBigmYPKXVsm2c7hSkog+XDX9MQYwJ2n
OuAUKfZZvWzc/nfGxGUAhD8oFVwjdj1hgs502qoZuVXnmYkolWaF7aaIpExZXFbLpLLDPJgVPVo6
u7rDCqxavVZIbL4bPoF8NODjyvYl9z6/ZykpY/Gv/OKCYTNeuaYlUi4mJj+o0yv7efR4vkc9uf43
S4CqLMz6HmWwxk5aNT8s6AStc+HnCzWCO6gvx+ofYZy3HoSdiXxOGU0X90IUXmt1zS7k1rsFmYwn
h61d+Fjnr4CR+C704U8WA5w8T4xcNioTMqcOLpp84Kvvq32uRyXd8X2TPB6KBhBAOkib8UbOukV8
rMFeroS9ySds++LVCdBP5xi51NSWvGAdGiTTNz0i4P+S7315TARf94r6eM3KDPGiPIAxT/OZjwqS
87amYECgx8BkVubsEV76EVk0eEQ6BMitufvOlQZNOtL+KYKaLJPXr4xTsW6ADaYKm6Gy5o/ec5/f
MDLKOCOj22a5GFgjSP+WHI5uk5BvRc0fC0SnRqtWNOsev2jzJB61FTq60z58dTZas194/dq1p6jO
IdloFLdli31wu9YfqtOkHA+EyvMI+8ObzWk+uTyU5hBLtzslIp09d3Jxh0aBT9qQltV1l9XACvim
phXMi4K+0Tk25DnssgA2WnFROyXZeL0uNZrG3oz4znVmbvCMk09isTS0cDB2sOzlzn/oLYB8e0HA
alik/PszQtZBEf12CgMpKn10WPj0Q8GC1rFkSyL4b4pDa1lqgXFeVASf99xWvmrAo60h50+Kwuge
xNDAc/OmnzUq1OtdMpHQYyJyCMugy9xm9swXU+SdRtDEk2TyMCwVlN1Pq6lEellBeYpcU9dRL/Mc
ucToGez0+BfFS2Zb8/tmDqLLI5gK3ZDh6Qdbg65nUR2H4thl98yKP18jYeE/tm8F/XSz6n76g/oz
zXsIJn64Fnec5MxBVgQ1i1ul1WxZ7BxNv+oVcnJuua/IHK7cfRXYYCP0jSnVN1oiGcC+gfLFdU2G
0lZWgTB406oTvkQ5aoCHoQz/wDrZgpBKfRBzn0ojZHtf9S2SPLeCyqZv5wknh3xhwy7/S2QpAc68
sxiFGg/0M/gK+pbtdr6+VYhqO7ctjLpiMd70d8ebhAwKWZLvnpfKIDGUe4jm7V/VR0L4vZmMsaZF
hgDWVMuyM+uRw543Uv9IIr0nIqZV2/xgLlZFv1U3m+sC2Ttm5pHE8GLVdhbwQyBlApkzgGO+Uqbm
CiRiwImsAoFE3nMRgR0VwHXoB2jru6quB+ed3vq3km70pHCAq5Jp6q9MVjqQgATCorvyMwWFwnPx
5iXqpXSjmJvlWl8zGnzGWw+IYyuqkPo5QPEE9cTLOOzz3xc8z4h5getI9snWEkMMfZ2H70MGhsks
EVO8SxAv8QybCwMg9LOMEGID/AOG9qt9D6wWSZt87/NlrXNzmlA49ZSNQpXcxmAUpaDhm5j0i4X3
5ggIya6ZoFR/ZngPXyUM/1C4BrpMuIk1Wrxf2S7m8gTFRmMqkUC/B+em/OpvoLKsPX1baKPxeXBN
7Zr3UAPFpee53YOLhQ7MAHmZY2NwO4IyfmZP1hGk5TKpNzhJ5iv2pNWuvgkPJAG63sN5PlfSFrh9
4GTEz9k3owS3CxI4oofn4BXxWPnZQ/9sFoA5DUohB++rnE/mqwYTd24DAybvbVpuoSJ8/8SJKSAw
wv+Qujyv6JPIYZ8gHwQZl1sk4muWm6BCiG3eQ6w16KRhLTIGHL33bAzee8PVHOm920faDrDXZZ5m
jphOwiIYWNQ4tz3/EtJK0mwryC6HuPHsQoasrNiASTkdNHgHRCobsm1mO5dsZTHiudsUjNX0eHEJ
gBYVRPT7ESyrlNjOu0zFVDlWA2uS9RUKkFBOxa1milRmx2O7GyDpdo60IM2AMMfYn1h/ECUZKUdf
OCW/ng+vTwnFWiXof3tkPbatZjugo0WKKyHIssFbf6UO3AW89fz50b4PFhh8zFKXH701SOYYTxju
DcAB0/piRKHkIoTIkPKN4ewefgDAzfQK9Stebrx+cmHNCz2n8j3lqqYQjyjUDPok0zLsOu9+6N8+
KlO00oZpwqEEc2z2V5ZnB1IVF9dilDm2jXzyXBjrCiv7jwfi59MbNNY7YzTTmYjdwY5MUhbCRbJc
2YMBmBLnF+4FsLcwU6Y49p5HAQtMZuEty92I/DJjzrooBcYVXFEaoXMokvy5SL/47M9Myq8BZX3z
ciYSpGSZz8G4LHYYOqKICevSg+iLNfy/OF0cu4QedPUHmGvVFdon2ZXiYdX1N09ArZF/Y7+Oorhf
XLqrKTbQNg2vP3c8HDxYsfon9ZTgIccAIFNTTtQN0R7xOwNlSSfh7pGKTWyz8S6bEWyzrvIVMW04
185q/LwdvLkZcoo3NuNJzaXjuC8O2i5pb0rKjfBWh6dp8nGqw9a0VFDyrkZPK6o41X1aN+eNpk2O
CChGkR4x2+u/Ogc2BOTqC8BeRJectmgAe46CEqTjdRlg4cxJn+F+E1PcXSnbsbAv/lsy+lcdT39p
KKFptMSaHF18bznXGgEpXl12VPciwAzTBztgoWNyG8zWjsHw7pqDACtOy37YW0jX1bzuC1aorbPh
Ux3anPi2bfXYtfPUEPhGRlF0UxFaaudcXi1LqaFxS4u6+PaFwSN5fi17Viac4UUDCZfe0ZTsEb7y
m0M1kFjph1aQFMZbMr3BRWFxU2W6I7HHBX+uA9fVyk5dl8/FTKUkaPuyCqnWEkO2kbuk8lSkI6/1
FF5VDmBRM4VelnGQrWHMaJ2fufI2x8PTcITzvAtpqIhAPqbSVY9i/giEwPawWvnGlglzhdHGg+UH
/w4yxd72t38EaCaJlqlQ/xjrqc6a10eD6B+K5iLwCT5LljefKyiTBDjYDNmJy+wnyqzWY1GR/aMF
O87Bb8l8P9RUtHA4AKpoUF85JK0YhtooxYvdIRHH7+fMJr/ylRkjW4RYnhdC7HPO4OeIxZMB5avO
ZDjbgmqqISB/hpVpefcmj2gQj01e0B8BqH7O7zUyVp293L8vn7p+SPOYWsuRc0MNq1RfqGDwKq77
rg0fXkUD/yhEMfR8EQtXGNqGp8RnxlwQyri75ULdQw4pDtI3ifql8ATyRg2TK6RIp2xJ5k4AJ81b
rUnxk7o91fy6W2r+HdY+df6yqKcNL/TVGxNZ/zwm4wjdU6VoN4pEMnVWz0PvczR6IUI4NQeRFWA8
SuCTAIvcrffXbvYdRPX8bHGp4ZeEchiuCQgzi9Pwv5nNCJLUSDVX1nNMwCT8gRPGejZyRO7oOn0F
R1oVFYUtOP8X7FrWKH7qi5uc2lLegtqIkpOd+QrEM3CmDbeblL1oPqlRk2OB3+T3EPII5OxxF4sr
Vc7OOTBn9FdY4gK7l0I/ARcXAJRk2Pns/TEAM7WM9sI05S35Nt+nIUiY6w3aMV/iUXIM4QmosbGY
h47g91tmEHLO0/f3m0hrPOTye1dwtW7Dr++1EhOfdTcz2wKFq0OHNVxqXOtkF+yctqT9iw6SCmEQ
ziFe8AET/OS/gE+/SrX6GYFX9zlJU/7Dp1hD/33u9KTpHEVf3lzOjElJ9fX/RbVlo0Ge7ETT5F0R
Qjmfo4Jlh+YhNbF0+kl1b7+fcyFP2vuyi/0t9OmWj2Npcv0wet42qlHV0VDw9ecAUDmXplE5+xS0
xNxF+tulD6uX4Rpyt7vsaXQd0rtiH40h3m9OtdyP6xFx0E6VZFQVfUimjUnkHQYsTMNYGYarMQJu
yf604Rd7ly1SaP4uOELfugWYqVQYeol2Cz/gjlnViRJ5yXtgMWo2pa9Rh6fatsm9pgXfRD8oigER
3krv/p7Qh0Cl84nlEp4lU3QxKcUzaFsOItC8QXcdjFgWGIt4FH725gIuEcOuLREpUAAYQyICV/Pf
yrxVQ6BB17sLihw+RM9KbahZvgHyvQfk8805Dot/oUG5dMCswVW+Xxd+9pd+CIYJ3EseKgekmHyt
Q7nlEXhTSPE6dRqHAcompFuhCgN1vulo84LyTBY/kvYdBxpkMT/g/gGkAlMegA58WBJvgXxHVlBO
puECPSJdONupWAQQ7WVkvMImSpMCl+1E3eswLWMA9etjY9UrBd/uqYnSZ0RFiJ9upk+eQdR4F8pt
ubRnGX3o30U9lVTAF+pegSva+LteFp+//3FjU17e8WSDzqvG7Ti0n73nvoulTkhx2+Cb09dJkY2g
TvsFz4B7b7bbYOkMYhD1qxOUC096e9+IPuky7G565zG7sU3yt7Z3p3LvR8CSiDI6pdlXA0+zjJJT
Yu7BVlbWzSHAagwhyY347uB9VFcyE/B+UQPwP9jFCArV/r2lEiHSZd9CpxgOh00unjwJf4+vOuXL
pdmSM4H73pj8ACj2o6FYKfTVETr5VhF3Nu7ZIXXvmjIrkm0Sj0jVOTERYqLsCUiA4nbSRzkbvEbT
bl3p1w/1XEslVj+YObkvEQ4fOtedDcogPG8olCo09k1mJknLlYX1Uzct7Lm9Ks4N7xRubJJmJOtC
+sifYOd2UkIH9un1Vj/jvfu3eoiblcrShd+xPja+xph/pzhmBDr2EcV5kg6JMQ14g/jDCqOHFcrR
6W7nwC4csryL4iwTnkrYeIZ/DtfntucMZvvv9P3fSkv41T5NknDUwr2InhdNdKh0Wpqaz1Y7UnST
kVD6ruWAvxB+D6h19BcllhoXKfuL5RJmJNEka7zYjlafs+uifz8kFZuPgWH1USIP5W/1RhpxpeJO
r0W//PojAzKpk0DjkVuyFLeKoJsw44dszcSnE0UXSK941t9HJEU3WBn1MLSRBvMKeazgp9jot2X1
u1z5tGYWJ8gj/a+ctGXQQnl9t8bOHuBeDh0wBvrY8nyxqEzA90wC6T5jui9oEZvFc5UW2CzCEd9/
LcJOJ+/KLBpMUyumQWlwW9lrYONBlVOblGWXdehgnPT6p16qET9JS9JhLPXdzRQ9OapNFIcJtEbS
UVfWO4xIlL23XyHZcW0g/8vWzHQ1c/iCGyDFq6y9eTiZYTL9CQmTYaU5s/U+mJK1IpUQscd85eg2
kT8l8qsXXvt9lqPTonDDFGStYI9GedaBzlWHloqkwXjZF90oaw1Up7fTypHGeXqWSmHqbzCPF7z+
BSHfprXtQiRA6Qg17W+Zfo0gJI7puGF+RXD1DYy2KXiwfsNX/Wl17k7JxWblJUITLlOZWHmSVIUu
tz0jlzDhWEJbIVgiLiPMqmQtkQv2VsWznN+iTAuoPHIQ2hk1nTTktx2D4huGKUrzOPPNm/tnRvXL
2rN7UOiN04JZVefzX/SaYoybMRMhLsD4C4M+0SYwho6Emgnpyv9ARbJCoeG66KrN0OMOeMsYl2UF
XQWiHtfMu6qYSiBw7NFf9Ae18ULAdX2vsLpw2c3PgEvxPcxNCPTiHcizqQ+sdwaab7RO3IiNx7wQ
EvxOJrbGBhpxayr8lKjLLMT/X4VnKAGDobUKdXJn2cO4B/TxsZs34zWytLo2p9nAL7DDsz0eDB/u
raUrGy58JeNRXwz9tLx7+TwQx+uBdS52UD6MV0U21HdgPdKsccDZplxStpk13/UUSjxaDjvt+aJR
vhYSQTTyT9BwdODSfC6DNeoRO1u1veORZp6/6UFyDzRUF1Y5fYTd5Hhc1o1SvHQ8tSwMvLSyzsZN
uXPqbtn7tMhvOw6mI1d6kOLLpe232tUaRcVp6QmzTsc//T/ahQsOrKxDQOZllPgfiyjMofwotNe7
sb4rs2g+Y1wExfqI9vBvfdTfDTCvbhjGgsIk2u0DPy8SkFRsV9sSyEMHOUSIeG3ZIvkXSWSktSHP
9+j6qdiyDxuU+Sy4zb7ZLvzSsbQnzJDq2xQWv2WKcblGkP9NR2fQSvobhI/j52d3ogyOt7iflku7
AwxG/3FpRXiinZPO5t/bEby11NxXSbmDxOdXIMEqoROYCQFXqqFX0Jfk4IIlGLd/Ux2ZWcEzOOUa
9GYOL2xDjbKH3JOQX9XnxcBYB3E+2YEzUc+V4lcpLSJCdUmZHMxhTYPkgCvJBYUpLP0HP+FnIioq
n/YWU5+EkcBck001LU6ffkV0cwROShdiZYToNvmR2L0zhlbkS9wJfG/b1FxKacAIa+yzETh2/svn
CPrriW9ICRIxe1UUhXQd/M3toKoEOvb/RPvJB3MSL1gAHkc4PRqrCSFsUysFArI+edrfahE7Hra9
WjWlAfgWNPCY1te8EanCQRXfk5aIB5leXX4v1Wliyi1Kgavrfx/xM+qoB5Uhja2KHloxqOACFWEK
yFcLuQ4YSHZ31HrNwFhPAp9bppQT88S+9AVs9yVM/kinsE/fgYTtJtadfVtYFiOFG+zTuiNY1iDt
szsW3UrovK6uBC35PiRRuml4Ca4foAW/7Qhg4IMJ/5wj89BtY/9BR9kpJQl6v5fbH5jBPlCAAeVM
UEMQP4kY3hGBmG04irKpFyPui+p2Qm2wsIMMBE1QXkiddYu9B/5h3nbedW7remYDJ2m3vDF/Rttm
QIPU9mVJLrvsmvcLayO6/sAZEoWTRU7JtMK0j2TmMsGGYrUHkV8n02a3V98u7sip8Nr8LRWE4dCl
QtbdG+hq8k2j832pwPn+nUdX9RTjruUzmScqhQOYxNPwX9Rt8nc2O3IB34535Szi8eAypBlu92kj
JD6u4+ytVUQ2JacC/aoFyacjpSVR/TbUJcZtnVOMBLcvly14booTmHS7Ur+O8lLRhlIVI459AnwI
KvT8zeddLfTi/JiYHr7gPcKu0Ggi1sZfqLHRU8RHf7+SHBTrPzJwzMWFveaoBg06KNjXqzq0laeF
szvdGsMwnai2w/OAub63JAIM9zM2uzPpUSr96BfAcj1gm08PcfJbVIsoAREao39pvxTyzr0hyjH1
tfUOFkgaWNOLHBnMOyDPpKm/PoVK6B0WCPtrX7wfsGP/n2KHir8/wdWI861pC5tANZP7E5aWibBV
AxgZKGxkLAlob1Wr+Cp5ra03wfQyWIB6loNN/28caW2RmbB7lo1xa66abWsJKaJJXUjhSAXM6Iit
ibMgab93rgcLG5qsNReHLNvuZnot+AxrNJaytmUO4AZEtDidRrpaKYkd+GKgI4tOb8Kx4VaLRyyl
sEyN2FHd9d/she6djj9Yg1W7mWxMeVwUbxeXb1XTKWz0hCOH+aiHbHkIt9K62aNweXeb/YTaUzwy
NWzJqU1l0XVzXobGN69S6xQwndA8K0XJ16ad4PDxB2cyVgeTsn1GZhOKYqdy5xuBY5Slwa74bt6+
3hGEA3pv0IEad0Ptiku1+N7xtUFKYJNz0PquKxxotNRZN53TVQ92w0BKF0p/Ez30wbZja1VzfyD6
YV8ZSIusmYw4xSx9AtZNhOAxHYf42P84duOhd9h21RVDmIzv2QHJDAjhYhDOkZuZkGSVh2oftTtj
IEtDIFlY/Wndo46pfc+LBS5ixB0as9GlnFn33djEE4KDiP7xKCyLrc18qJKsJZAPNrJfCVS7USr9
o3ZRTRxUAUm4qUC0uG0UOcgNuZ6zqEJox5HyImB5yqNlsow5fNt85UzpDbGDtHAEn15Mfr8A9qPA
oAce0X3dzv61GEIfGtzRTyLTPz5bXMIAW978vBuiKmJclLtmEnM0kIsRULVCq7UP06b4USIu7W77
PNWfiJmTK8g6ZxHGm2KyaXhMpbRjdH628HSD4Hwr67/qlqoO5z1UK23bMW91W1UI2QuX6pXj6XmF
QQNxyUEiu6gXV6IiFFLkeQSnYaEsvvNQ/VROKZKWfLoNNGX784FrGjeiUUzrDzLbMKqmllHG3o6h
roIhv3DIw0W4JyRSlGyYmU0CBCIrnNMVgDoma4uTgU8C+GHtDZHoSvmoXAySIyOosM5okr8TMmkE
ijaDZ+1D+GLpyBMCPOwfCRQ6M6PuyLMp8V+6OT4QPxkfWZhH711OD6//QZHjcjAULRII3z8wU6vL
AXkpRAhf7qeBdkbRjw2BHW6PaeYRau5Jd/ga2SQk0+7x0DJ8q32f2xxwQBaI/9RfCH1wjYfPdFER
3bHa376OQO6tU+UvCjhdAHeh29K25+6jwG+8rB+QIdyKLe/1d/kuKdN0RZ3OrT4USVK87wwf2CTQ
yQvym+V994yRaxUlETvlpTcAbrSxR//SG+atn94pslbwf9DWl4Ib7EtLlmK+XiT4V8c4YaemReSy
V74pdfLWqK448UYT4Tzv5fUS9vLsVIXElqw88JD019jaGRhW1/U3oZ+8ygvCUsEZ3lt24iPf6gJW
omausiCwi2KBHAtWMswBrFC40HgiCXaTyYCPOc7A/rub0+r6tDnbF3BizYa4tmGHhAvBPCcpf2ao
KXuA0zr1MMDpqhWe8fDIPF+x9gsMsNCBoqe/ixS1IMjN4KO2KaPh2KgXXw0sZSkbVqqIbLGbFGxW
l778ewlewQpKJiFQxREYyW7JpA4QNQB4qjvq9ujtjRiPMK1f3mCaOPDQISahzoh8D4Ss/F/qAEaZ
rawhZUnhYlpog8wv8mK2jRHbxYCOLygIy+3F/LjfDHbWo8BP0r4qD7Tu8mfJtxkpGjOHqA560lJT
6too82jwdZmrF0N3dQQhsGwmUH4nDX/vwcNpSSoCyqeurG/VFfKfDsMCa7VD0gEj4nq7gOfeNKoN
AARtAv7J9bOxd2kWHR1euFj3a/XoOTenyRcdF8inInTmY6J2z98g3PVpNPdJ4x7FpK2zKGtrfJrd
xj1jsUhCkqiJ4pxJiDKZ8r3a7oPOchSQuauiiwDl9hgCBFy+bJJy0+awh6+iHuJKnxMEScTL4meV
4ccTvCPodCVXyOsRzWE1ZdkPYnDGL9HdhJqE0ISAPEmK2Ut2BL8ZgPvEkJJmpdste/9SsnZ+GA5m
tr/AkIFkGXtL0Q8j4eY1vimLPWA7p/4uXRUsiFgctAwcICrBnJT67LeKF45QwJvFo6UuT02pygyW
qwaOgmtNVip+UB5tUxnsbkJhaP/SD5GSPhcYahG3yAIQfrDII2eq2RgdKqx2HfU5/VjfPFJuL3R8
x4GDnpAGdw7L+61mr6qO8OcsyjZWAhOf2jcB9AzM63OCwc7+n0pRC3QZRhhdQVP70MABaWzHLqm0
OUAPRj0nQF8gsnUFLdLFeHHaVOQB5IhOBYd8Hy5XIVNV/asOdU5Npm+NV1mBPK8lk9vprD/rrDBg
qsPkO+/sEaXwyxOnaJ1BawerDnhfrkMmwOIrI1tr5NXzMtd2x34yVZ+lBqCZHI/ybxKdLiDH+QKo
6jQRcbmgkZlp1X5RPCz/gBRXiLPUvc6+BGUDsWEGlJuDNwb4h57F9Xg/HtExnbBdgYGjH3TmVrZ+
tMf5uoIhRD2KgMBmcww1arO1VYfs9peje5C4SbW0Bi7FbJ3MscN12FA1GaVSzb422OGvxRJ/AV/3
EkCHHF+kGNpY/LCnomIiIfa1sNqZvFSPsg+OpS+jM5LsBW1/Q5Tw5iUGm4ltjwT0LklP93YSHGB4
laAIKHWmONBASbZU6oq4HnO2GnwZZtC9HolQU21+iXcJZNvwcd6ATDqtnO+pQbhSfKpGyMn1iRQE
8wIIXb09uR9r076wWU4tEXgdjud7yi4Gd9DoIiLMrOK9HubLZAfC86V4EmSE2ImFy4bGxI7M9QQc
NtisBsg8etRL8jJozlUpbpRvRMWXu6QgvfutZbTQQXOQ2Ug+TI2HQML2C3PAITKS7nIVwDqlSSLh
Pu83SSKGiU4WazspQ7ljLgG2bkFpiyO+QeKklcVUqP2wzuJ0l1aW3pXIvaxwP3CQc9USFWtNliTj
/zMNxXlRFuUbEL+uXoPzFL60snXmxOC5IVKvlMXAyJxApCbzd20aOGN39r99rOyqlu1JFOzYjelb
iAcmJgyGmk9b0ximocVgQRlqtBqHlHPot9ukl3uYvDEswgF4eiZumxPPOqvXFLLtujm9D9sADgF0
JWqtPC8HO78HTrmQzgYIMxYESh2X28eNAKjNR4fGtb9LUb2tDdOlkPsRM8xWGsBfr+g/OgyZ2Jb0
F+Kl4fXXLDN+efS8snTvvn4kFQ58OHZ2b/+qdH7bjdt/GswlVVN5SWIVMQicuVBKg5Hs/gClBIlK
B1qV/TbQvV3+nfSI8N3OZmvCa0dWHdtj7wowwGxPT1BRmMDZcga2QbeeYCVkFgSOYIOKfGD5dfob
Ww2aj7tUKj7Ko4TM1dMKXmNUIYtck82Uc3e2e82xp8JIjpoeuxjWIF1O9xl+039Krn75dHsCfC55
2MHhdb6Nw0MIjE9pHLuooU9MmwWVM0grNv2P7PTtgiIpPmZHcd4AcgUhezf9kze+l3J1YzK9+tDA
xV+/801bZJTH8LfQsVqNCtkWtq1mXdvoRmqHZLA2exCU8ttNGU7WdnrhUSQoBHSx/gJNuKeFlhyY
SF5dZzhdICSu/StGUXZCxANVd/UAk1aL5zh89ebaHY+QILxIX4S4nN6ZG1W9Th8ip4XLa5LxRhGH
ghT0kWo5HunXiWpBA74O1tYzqZQSz9Q00MB1Jms0m+ra/giCrGvyQKOgZAq0afFwAK4hZOAcg41Q
tXA3I7WJnlyIUAmtObb8mDN4kn4OzFLugGnbNVwAn3NimhE7PR/NyK+x1w042CV2ELIEb/L3Mxfx
JfDi2yMkGFdmLxawcmYXjWQGC+hfqGpkOULWnexv5AESD7Nd+CnqEh1fD+baE9fqug424y6iylpQ
EW6xFQRb4/HqWGuwICq2zuPwLp3wLI6RmcKXxc78pZrdE14Nxbgf45tUr2i455VRDHz4ZT05wQZQ
dEG/1ebe0rZOby2g/tF7Dagxvka3/4xPDE+t49wo6b8EhhSMyrm0INp7xlgML3X/ZEqbTW6ah16f
ylK1SZJfoY6beeDPjcOXg/k0UQRd26CPfEmxhzqxuGe48UYHYVv9Y+B4vZnliK9WJyP8rLiqlPm7
M28S1BYNEpL/pXIB6NTUYsLg3pV+m1PDQ+FZdBBj++GjFcRhu9Yi7Xbe0hjyJSi0giatQsNkWYuu
btvGu2/5uH9aHnYMvUAIhrSmfD/m1j/EZRABjb0A/R8yZsdJSZJ+VPJUzsvGUnlok4WGD5PxthnI
E8rQYhkMb6qkUcs1Te1hM81d+rQuh0ASokM9U+pzGiSgF1MKLDvb74cybFFoyxVc+Da48R3EjCYX
YVHMNE2+wZ375+vYkA72ej2kJp4RI07SnKsJftKMqJVO8ugjOGtp0gJb6sFSSp0piogQXk7l5z6w
E+dAR4kEO5UWGDZsNYuNweDortZQnAa0pFHi8dQZM2BzKflIaKVA2fl5K8UY2DGU5gitS8eiIeK0
w+7NzXSg7BNS6ExCqyRCWoaBIt0IiHL99ezbHg10C4ID9QUJw0Hg9dGWgNZHiKrMdZNlN/kPt8p0
4rqLCL9plqMM39t1RVJKPGX8ZnqjRHn6pN64qaUfKVfjUOAzyG2aLDUcAD03k9bBGv5g9jziOIbI
JY19gKYxl9QHz/G8w6RfkmCArvWUNAqBvPGhEAjGPhxaj5M77WFWh6fsqV0VOIcRThbr2v5jK+MJ
WUxQQE3aPx/O9+K/hD7L7pjIDWP+k9ay9blu3DalYakCFljZK4MwPGGhAsgGdiER1xwl5GaNGVLU
dRTZ8dT6Ed5BLPDkz8sOb/anPh1KGmPfzYD+Jws/6gphsYQ/OOAzljdG2SAMUb3sjx7kKmo2d/8z
P1KbTtzeibnqDugCNwATxNSHwEol3mcCuILjCzSGUQHX6UPZOoDvDADZvRBNP7/9zSGS8OGZcmwv
BYBE/TNaTMq3EEU5Aw8f2FGWn8b0hDZaxhGwKaxfNFkgcv2iy7ZN11s8C0w2ouSXWRF/gz+xXJd+
jTfntkkIPsJoetIQkQ3pcnx5eOGaMG1Csdyo37+0xay70h/cj+fitEcTQ1IUCMeleqGX5sA1rOnx
Tqm4caa4t5CGYK6b3nhj1Iw0mwqE44spkiHJzVVCX+0WhCRS+wxwO+r3Jc/xslbHEqhrwboy6ZOY
KJUyjjl8a4YWiS2urPK1hC+4AUMITu0sW6gFZTAg/Z8ptyPbd+sAjzjRAQY79MVfoLLG+wFDlEpd
CjivhkPY7GcBNO8ktRO3jypKqlttWwS0W5bPdXJzQHyf5TU6oApAoaRbBNuZ2bWKde6RUjHKCl+R
Y63M1GOoRocY9LPf84OrlieOUaTmSZt9wzWgXOYAEA81GGYIGTh6opNsIU4PmNdn1P+RHGyxFl7f
fUdcQhb6t7pUPhTMdAhTmUEnzMEikimqCON3QtzHoVSQjtqFP/Z8d08149PNMjhqiNLbrbK+IPQy
ZRFxVXDWQY8EA9GDtfPoOyR9diCqAA5xyyJCPTt/b2pfM80hM7e0PffUhX2dn8Euv+nAfbQw12ZL
ZcqfzGasw2gKSMtIG5MSb+fbFEadplLd+NwvG5YPc/lNHze9KqJLNnFFw0SO2OTDPDD2+4QMxxI8
qMg65pjXOe/I6sk2rcnOsV6zR8n1c8upr5xNup9rQx1j7j5W8V6a61n1MeN31/+11lgE48AbZrTN
ll0RnVWhYzWMKcAQOC5R0Y5JAFGO7/YnXINDvI859tzG7Fsj6bpce3Z/dV9bCJb2uUugxCVLUNJv
BmcH6XElPrFgDFQKR0eD+QDPM6O02zbR++DHehcvq7kYImb26288brgEvNBs6KD52Q496mPMrWeI
fPRqk5jZX3TRYZeOOSKR2Kfjj3bvEPpRcKmC/T+xLNL4FIccEQye687Q6CtKi2KNvYg3LCNAXwRc
yf1NFY6rwns/x5WOg+eCeYV6z5x2QbcNNxJUENJy3HTGFA5m9TYFFmxrk72+YXJj9eRtnJZsufGq
6OBRs9WPbU3W/8iFZk/OB0nmp0yFLf5iqsGj1A0NeTbI3PYQJipSiMYqluTrTEfm0/2w1sl+rzAI
swXSOglwK9roytuvww7JzVeor76R5hQ7Vyt2iFcOfiTB1FTcoAAKEyyyUrDq0X0E+zdC3+jH5yJn
ALwod28saGM0C7lqoIkDcN4Atu9JmqlGR28gGS7eBc9A24YENtuRUXPFFWVHDS98WxRGd40a2QKd
siZo5GWgvHMUrczo/QFdjd7lWmEXqdLXjrkcHdu/g1Idthxc52fmHGS0uXlPOZZt0iUQCmZ0cvep
jANHuqPMJd/N0OmSDWThpBK1IfsooYJOcJu2ODvb+fzaD9ZJrwgVRQuLtKU9C7PKcEjIO/CLAzDX
rgILUXW8KFjYGl3fyWcQ3WgfXmJsWUxMhMYyfBcRFpaW9GpDLnCM9TVrVjUll14w17JFAk4vdLMG
paSgu3BiXLhp+zypvoKBSeZ+eCSqyDJ0zwe0hi4bCAbQk+gJ/nh5AMSpuztlvSuyGbSwz3hD+OIG
hWn4WHYkCt15STupb+Q2f8gm2NdtfZTOpYz+WHhuwdcc29Tmxs2i8IOrzaTkuqxrGraAJcOOp57m
J8pU78g017h05mrsE0FAFmhsXeTTNkz8rjkfHGibVSULJtNs5WK3Pu+6b1AYlTUn8pkEh+SC/jME
mAjZoA0eTiW63yEr0ITGguxRuOIEYz4LKzxBOkj276gS2uYR4jM0ryg5Z9kqU7hLznUM5hvTl1p2
geR9jW5LdgwAlTWoTnxvVW2lWL0/GnEyuI6Ygx2/3nZG+VTrzrJcKHOGWoCj0AmsNHFSCgOhunhd
VxqhlVUANig2Y8LnNJTOrsAu3tdV6KiGbAGm7tIuRiqmvLU22MJcnKoo00pfgzxQTCYLc2+vOGgJ
WP5S2pEgwZ20cQA0D2/OzXdNnGlZZAOJOq4mHFWo/gasTrIHYyKTs9oMA2uIDlHywahC/p1BSphc
lPGLCKtrF2Kwj7Dq3kbCk5gXfwn081ly+cYE4Dusea+Pu1KH0pFixJmqucNuIXNONdtG6Z4OWial
vto+85ynkFUYsxM4GOWG4YQjEv+zauNS29/9FVcHICPkgNe1ckfEK1UMJNmCKKBgOfw2eTNE48dD
TTVuOn5eddiqSYkm9qn/gH3z/la1GOxYb+0URrCdJM/GWkAeOCZ4kwBFn/6a0zDoriBdqq5FIXG8
ykiG7o8Py/cKUUvYQgVNg7Ebf4Ib9VIOz3Giq/8n+9vpLvM2/RN5L8y4EIREJjdVCwYFZ1a83wPC
rxIfGRE1ZTHqTwQTjTWWlVljgiGAOl8vEkYPloHt5TuB+ceru+Nz2jtK6wciPxksyDaNiGYfSij/
Ps4MunAB+yJNPrIssu6FnYiMtK1/IooQ59Uo/AvSX9qEw742+IaSauftFMNomn0peRn/PQvOu1Dl
0k9o3lbLFcCjZ51pu6scT2GzHZEswhhFf5lYxRkywrfDta958I9eqGDkM/EUnO7Cb0BxS2jewTki
iuyCfNC3djSkTz3xmu+hdVRKm6BONH53NoKg8a2pQ/ucgu1tjYnmuqEGagQ7fmc7FOYteqZ+itVn
nFcxFC73gqF7xed37MtymmGD96OZ0DxYLKti5NHaOUFrmfNtkQsvR6xHtTRtYHwk5r7y1zrnQOrZ
MLJcM8tcAnzNPErohieI+qmKclRUklVbF5rrM73n7eYv9gy/nRKAARyhXx1+RFvbiVvTXclKcVdN
wJxh94MaaalFh6HJPtvrblMU0FTpd4kPbf8tjnrrmzDq8yL39N7KI+qs/ih8EKoZVVh7cVQs/stm
mq4Rbjdbqgu+kgUYsGeW83zt2XZVntdEtDogZL7MyAJ0P476qtgaM854OBmz+pDcVzifPJKgjj7z
vGmHwaaLfupmTjxk4bG5mUdXOQ9jv88308HOfEzQo3YGNU27bha3fiDRnl8KyviB2JGPI54/SyAI
pMPv8ji1NiQGffG6X8hot3pwsUomrU/fS44dJgfFbqhZ+F6PeyG2UQ2aKD57jcCFdFhmkJjBDsjx
jYqfOb+aPQPKS+exMr9EKofbFf+3XCvJUiD5z6yIINderuijYEoQ2A7wp613rOsqPQX8KDU+fsQR
u0th2eTm5hpcvGGvbWq6j5SM+5uL4zNlj/Ge+ugwscT4KaHe+OI3eoawyAmu5/ix1QBm5XbkTMLW
UQD/WhhTl/HIkrBHTD6113STCz54aIGDVF0/sQWJTXBSiPk96SOZejwhS19o/HzymJs9smYYKYOt
Chtze//4W7pKkeG31odRmcuf6RdoN0Gr+BkqHH3+yCSA8jNr/YseSqAU9ABB0K6kM5SxKLKfYEP9
P9GGYPhp6veUfgm48id1DJwxVDrdRR29PCVik7igcKFcnDAnoCMB8zM8VFt8CC8fGGonRU844ML5
idhs/xc/xdkTV8u+9kmm27sS+WTTNdckHAaPtbeKSZvN+uzNbPr66DZ3W0JrlDEIdd2dUkL8UBAY
N5ndImqCVJ9lc9Xs9QQFUZNS8Knu/4t4Qr55GegkPSmHaBies1OkFGIdgjKCEj0vj3bRaIv/Ug3u
4zT4aGnKnEACsrbShO0DzqQhnbYQCAwV5h9+ZyybdL5XD2y7wij8dSa0G/KKwE4rX/kbT6o24Zhm
f9w+nV4GwFcwKfqzsi/uwA8IWC5U43XFjRseguFEf8eFBJKl1e5ZsrgFYlshQurBbHG8Ypl/+Rj8
vFiaUQqkj2BuyaFXSZoeTnmTQCsatCegP1ZNM6edo7KfcThJpQ0O+i5+YvEql4kp7SY2i2CIT8ag
fmCTVMGA1EF55sHOdrEvR8uOqUJW6bcWGLZ3GQ+sSPON0gxpb4N3EX8lQF8BLQ/enTooE33L74zE
tuy68+VQWoguXfIkRfVLl8q58nmmdCT+zi7FiM3Gjl7BRtuMez/SaeDRFnWgMqC+9BgFoV5CdI6z
WilSgNSrm1ZdNvR5NMTCBx0JkxfO/sqVaB3YhVdEbxhC5/+hZ6d3XkM9KYzPV0IT8RCb7+4t2aop
GnS0XCD5gT3GGqWU/KDk93EycRldaAC8/qemQa21K3UXDOMwujx2SwM79u46VFucwAwo0GDryKYt
sEsvNE+nopJEVDVfQYClgKwkDsCYURQBNZ+T9CZpoA/woB9Vmrh2Piy1ObeZpbV8b3GN06T2Hei5
2/qm+xAWoAmWM64+JCO04Xa5GuINZPXkao9upXWlfY/qaYUL7YADQ4ATYA67xhhyNe7z1e7A/IOT
R/lF4lRHHKco92AAmCnde/YXovWpoHWiurhAM+H5BOd8XRhDr3WvvYk9+nI29ptDwb8Xl3/CD8Bw
bUlW6eGf9Rb8ypWpCq+B71H34pc6gXfJ2kvE3/90sN+SiHK4ZgSG8JU0giC/z5e2aRYELBn51q6V
kQk0ps4LD3c0NEBsFoTHFjUdToIasQoZHFnvXBxjRJ5d+J1vnmr4EjPZq+P4mCE0i7jACmypIARS
qD2MgKxXoKpC4iXMhs0X01X4vZyarhQcX7U0qjbysc7Utb/PGPFetpZwDO42Jq37tcUWqPDVcnru
K9AtThklYB1it0ezB1fKkJFIbb2EedNnZkH8nPFp1s6MrlZFy1rl5Fqy3dtznhH4TQa2PvcFcdqJ
sZt2I3FwpJy7d9gnvVImt+GJvjrKt2cDllWWTh2FGxQ6poPe3fhFIeKi0wHoA8VLD09jJGLWSTkh
A8mZo+9kNXnPcWacXkjo68WG2F7p8W9Z05NFQXYNHD375Z/q5IYbpUUq/ZU18OuTfhJyfAylBjlH
oLbDyiw/jrr/WwgaU80rt3Y0TzIhaIc3UEbQ6OAFSZ9VbDpdmCzyYsT8B+zArZmdkXr7CCEg6dno
LG2GIU6Tjh0iTqBWkmFVL7VeUaZirV4PCybJo0E8v7Aez3V+eGKeZ9n+kbCah+BFwxQUH9xQRQqG
QQyulyzYfAfAk/Td34ow/h9p60FRqDGWeYNYjRXXslf/K1d9ROEXs//eFA5UVQNN5TKYkWgyoAEw
SKG4J2+uK3mXbC3MCjXA7Ek5MYldUQw/icxx6hXjK3N7rk/rIUkta9sTObkVhxlutGW1ob04aZB8
iFeaWdRPGpagKdecv7rpd3pWzyNkZ1JAbj4/4xQcnx2sz9N9psXyr89qb32hANYjuBAJUTsk2rJK
w2u0uzlfdOKMQGck/XJiMfkP2HfVTRpetMBojPqGL7EGviHzyTq/PxurKpnHJO1/HJAggUphj9YX
bSju/aZkhUyN0a+Jv3ZAGtU+sVEQk7+nRTrjS86nt5qHSFBFHsbxoH04ofA174ilVRJaNFgUsci3
WE2BvRgOxnTKHgiD6Iz+tBT2AER74igcR5ZBAupU9+zqsAGgAOKuXP8TVZAMAUUaTNZXIrRz8b+e
bQu9BqDw1LOZTuklZDtpSwGiV7iA3VVP9TuhhOYSvYaLFaiTAMGFYjKEYRZbDSuxhsu+tMdkjtYF
yzmBaAogIBSW8qwsaSMeNm++hqeHBBPrQaijn4IJVGprV+8c95/6Rz//BnfNJVdOkeLEysqu0wYr
4Jfe0WFddY2KwjTHTfeqw0cWkhfusBdlQn1uSOoE8rnQ0heR/u5CfzcFWuF2iq5oJkt4PJ/+kMiL
8AzK+0eu8V/nGd6bFd+7FrKXJWHrvar0KSWOe9iB8PIrQalAWIrPXhN1NmUsKs70yZ4JnMg4APn6
pCw/6fV8pbf146dt/regxlH+wDgzMq5jQCppHeQVPYQHZPU66AYQYXOT256sB9V8SfzffsEdy0PO
A02MRwsbAsUi5N1GtoWRXnA7s6dP2OQk3ECW8SFCcMhe0gl/mCmcjmgna36ShSAwmFPYf8rLKSDW
Jd3yGz1K7zuIceqyCjJPAgOg4X46If1fptvJ6CqZyoWIzmDoCjaPnEJGhi3L6d55VR8Y2Q+rquZN
nHvi3CSXQOxnIB0axzxEJTbClWA/osrrt33UrD4PlUJuUnLE9aVOZCRBDcz9MFv+QT3JN9959gRD
w/lg/Bafpc+yYp3lvccop+nlUeqo4vsl8meGbP+Mddom1sxMt2wzyZjPKCZ9ztOWLE6v5W39dcNf
YEPyNkGAPpxej5wdGMJfccyCsb107vQcN9A6zD979ptDQ6vOY/DDAgIv9Es69+/wSRVrimVDqB6T
gJ/jJGmdcWWAVgIhd12d9zcIfXKC3+QSd7I6FPMHEF3Bb3uao3Wzh6kVgsDWACaB7tPpDX3Fds62
zBF5P6g0RM2fBEnsuDGOjDFpCH8jelTLCxoXe6xmzF/3o4WLLrbs+muDCEeNozG0tauX7gdR1u/w
O4oNDFzGPxAhlJTTwNO/6ggpY1HWxBIwpcK/VTwoWyvknoY/P+54kOHk4NbNC2SUxJw/ZpE8t60Y
oJ8WERCmcusxhjbgR/a/3VLoWqkXvZWvbHAt8aTINaK77zGW6S2x9bvvz/oAPYiBNzlol3QwVMuW
z0Ij3IX/GBwY5H2EARw/oIdBgGFWXZTILd5vNhMHGbLidaG1omAtpqVuWiosXIOnLKJblpnTyYYb
FCOXhDglDq5+oCsiV+hjaN2blMce1fJBwlIFZAoQotTErobeMiok2g/x9FMIJy2OeMUb/gPPX3pE
qXRvPYPra0aiF5v0PGpecQHlDXkS/0ueB+Zmj8Ot6o38rBxzIWP21DhnVG35EX4vOYR3dJdGHvMg
xTZ+UYqfjH7L3fhyxHE7T6At2RoEyI+9PihC2wf70Ui4o0C8eKxrfH1Pz9m4HYSQZHU/ELUSI1jw
SgOKjHUNrBf0R35DuC/REid/AebEKBKdv30sWUVM0Hi9/OSjWGzC+R/yLd0T21E/IUMcu86cq84I
7gGv2zdTw8lxzRqY30leMoup58eK7PtYeMMOjKWp1+8jJmCw7bryNgI9VeRArSVDi9jcevaZ1SeA
gtJB06rg3bJ5K966cfNuM8SwS0zZ6VClLfbdtKBJp9qBlINwJr/YoNFmn8MzOXbn8NYeS/5Gh/8o
55VLOuSlaig7gY2FlCXCJGcbGY2UIXSx3ds6lmjYpcF8S34cUiEtxfiKGkYSVhDJ94Kbo6n4S9qA
YTIk35lJL/pkOf2AX37F5Zty/HAAahjhNut9OnaKvHAMg38t8P/7H53e/FpAEwZIU4naiVLveT/R
gOtg4VBXWFmxyItbThbma6TmYVXLXTmNQL9mw7zHMq69MAVQIlGNPWNKfu8zEc6EyHqnFHgoHCzy
BTZXDyKr//iP27/ERPjVHjcEpysH0dLQzmxPNTK7ve4sH7m0R21jaeCkS+LdDOPARSMQuxpGKYi7
84TjfOvzV1JkOgFLbmIpSUBGQSApwHT5Yzx+IA3+noOdDDOQzvukfe8uOOI1TLT3rJfjtGPvm8M/
BDYJW7ppKJtxN0HJbfHPlu+msNIsZioQYKJMNLY6AwnEOP/J1T6CPvs24q6Wb6AQbRKXIfFVBpZD
d8riW2sykoG8Fsax4Scd2uIfi8BP2NQY78EXY+LHxKFzUZBRhORMf7LZzeQbD5G727aTjyigVMfb
o/jSd1rk+/xGe6YMourOoqokvcH73Drhp4s8SnhdSZ5a6PZr9aQ5pi2RfMNh02b24OPfA9lHmFcr
EUAsKyqIOdlE0a38ylKC/ZvXYR3vLz0UrE8jCVB7h1kvuJXI0ZpymBy1ZvJHKIwUJRZydi5RIqkr
FgfuPvAq0A0FWTamyKLkIhTdCjQJdgtOY9D65CIPZot0bfiW/mnZ1kMJEipLOjYdDqHmXTlZZBOL
zWHNJmWOTl/XDvgpaDQnt2w+n1pkuZUSiTvc18Fcn2hqEzdDMPgVwovASHpsfFHGzIjoQJ4pIOFK
ZT+zytiqJuUTakkAfWTdsd15hKbVSDacrtP332fLTneEP/JXBSaxpqFdBZKCw1lvZyUbAA+eCQ0N
2JgNDbtB5IiwXzUlSGzqZ6kkN2K+atH0KMhUlBXy+7d/vguZcdLyAYNvDC7W0lELnklZEkmWU/vk
MVwMXuBUK9s8I7Eu6kQNBgrwue7cv0TrRr16uy2lhw2HFYUnvrJ6+JCZdQsuuUpfvXgZaq+JrgtU
GNpyFDd+m5jTU2K9udza9uhrllVZIbjY5T+f5jOCM/YM191+iK0kkqPIM99cPij3wViLUo5NaxLO
QjL7mXadD07IaSbmNeOpybM43wRAR80+IKV/6zmF7a/9/+Mb4TyDS9hJ65Qq1c9ObYsGs4yGD48t
FcAb66J2jzbSqqatwF7MspDJtb+WgQUCcF3J/y+RYeXIJj/Gg3bppOf4pisGFU+5rcxnE+truF2/
huheSfdXWE7slxNaHILm1D4RvOAADvhFi54/ZVY2gUrY34Zu48vOG3DyE/u0HcPsAh/zC9Axj0lB
+3XgHU7pZYE0e4ly4rxyoJiJlw7C/zE3Reqwbf7GYNHXYDYviuToXwQKmAhx8GVrjtJy0XqBbl0T
EE5iQI09Zf/8dUjDrZgteVSg509nUiQPzJ315572dKZqrmYY6KB5wHBhEXMtbLhokRGjrk3A0Vba
jAtgBOj970WvxPtdaYLDil2/qMr4csrbnPSzh1wC/dcj+0Nee71fPMzJzmIqA3IGGnyCRhipAOw1
nz2bnfpnkk7zzq7r5On+JwEnSdoKDxss/k7nTpWBfont70VQWpXpYB41wR1tJjn51YhScarFxOvJ
TqizH/9WkXMlzEq1+P6bYDjsHUAnC8MjR/4z6ZXvwjuWtFXINdh8AEYuWW/G/ue267ifIwQufuEi
Gac4sDtzrZfXFdgwyJgpPaaUYO/u8AYBb3xqbhhhEVKlmuQIe5Zuw4nT0ByXi64qLdXijgnEkiYm
sQ0wznGFfWACgX9DpuUFDI+Teul6nBSUvPupgAqXF464apHIg9ejW+TON6ewEKcaAOuiJavDHKc0
Ec4bfonhWH08G7y7Suf2NPJ6ksSTxeUCB/zHCKjYnaeKjx+89lD3NNMB4d6KEBi28Ef2JcW7MuCJ
ixnHYctRNfdKGKtO11F1i7Yi8YeqQ0+/9KSVD5sCHh7korKhsArt+UTifKS7wzzLY+vmhU6EmErh
n7fpIsBiTg08NfWUdYlPmycIKAgnHc98ip4cHXFh6yV9jtLsl6ivaRegV+N9MfTll1zcIIGpywrh
rYd/pMml32dgvBkaMFSASh5j3Og9b8u7t25zvXVCE6vdOaUZz7CvpBlIA2UajbpWrqIlyZkK0zML
A+9kG1wysyuHOh3p3ImtzEJqOKanhLRRJnhfPwqFZG0q0JQrUpZ/6SsflOuOHNPnDmcBJdzC1a5l
jDRPlDq6GTvqx8fkJB4xQ9yKC7A8I4tazwToOLrmzBvzkSSoYVUGG8u3BE+rpsEThdlhURy2RnD0
qbq4KsWRzrjHqysXgRbqQ6QTkw+do029+xUNiQQvm1sUQlHPrn2IRU3ZmFcpp5wcC8MfQskrfrYu
+Rc2JNUwYiQui9F5BRczTrxqL6OVuOl/NumynjtCNHDqVIvdGFC1kNLIZfq6qbbSgwodvqMMsJMT
r6e17JJRZbJbGgmELYHb7WCYOvjouA14WqnnmKe7vtACplhpYyruE2N3VsTCm2DNyP3W4KBPnj7B
/8GWWI3pUk4JqjDOQvXYT/iU80HFTbxgUi5Sc3XaN9ViBcYP5wOa2rXTrxVlWLO85TdFFvRMkg6x
gapZ10Hg3/6y45H6Wx4qhCu4eAWJAhTXOhKuiCc9LNS2pZ60mCeD9uJWI+plDhDStweoaH5uqqDh
9oW0TSNRGOhyOhucwU0kNwWoiJco2Odw4e0lurvT5+389zeZz2OOgwc51d2Yjct/aC6WXXJ/2mNl
ryXywlpBdjfUSq4GJaxvgq2fU6wWHPW0M7uNfA3csORcMfF6Ooh8CNAHoXGPzxtSW8Hrn1v8ijFU
NWkvL9iDgV/F3+UTj/GgNdhHNGXotT27nzxghmDeJwcTWltddRJMNrBKLdgSjVRKc/jIToTYJ5mu
tPclh2TqbWskWIYqe4Ocxwg0LMzGwWh4JI32EqioesRaugbrxI8aegCT/WkZRkRtuOic4tS22EFf
7ceQleEDR+xHslwvAqU6rohLlGwI2w1kBgvzhuDSfHnovTTuZ/xdO4c3ucQ0b3yQGorlZPy7F1Ad
oOS/x4F3fiyFWQz2Vs7OgmePt15tLG2gYs3xrUZKi1l+8ssC19NBuVM1mgBXuV0plIZwUIOjdCiO
wuxy9D7Wfwx5uTnt39wMt9Dn2PzBmbIf/wHiNR3zk3oxvaBUrYYfPb8XQhIXKX9crhOdBIvXK/6W
eEwk+ZlSsaBvNvo6K3xFrAv800d2OJJeywsxUAre/PVgvJcOUDAbEQqnuftMA210OOEpERUqBoeA
sG4VcXWZeDR6V0YpOprCzSrgtxfR5VFZ6UdtThsSEhyqgwW+G8AqgJ+eVTg0bgRofmLW8zp0uHGi
Du6BCSRO3jPZq35B4nQ+BHtXUGILb+ygtbKTdjbbgjw7Mk+MTzD8KwVoHz5CxJjNsyRnzMjA8T6a
gicR5zD40lZX4Zw0Uaf+WCmUrWJQOPxkMb0eRuOTeqV49xZTmjwqGzobtXIBLngk/7LzS73a/wan
9GTq+6oumwMcHqthonV9HNwwTSVDBYPI+Hmmcf5vfsS7swh/wCUspJRRj1ZDaGtUppVUufA+Kjb8
8ZFFM2QGIYdpVz2JKFfdmcboqgATCIqOLPz7K0bJnsVP/zxuCMhwTQiD/sTkrKtpS/oKCOM5R720
qgoJxkpohZvyFa0mGfOhQUA24+whlW9vzusKRlcnKQRBtxYTlAg+n+LO/UOqvw2h+SrIo5ZzX5Tc
zOUHFrw0TKJg4TF8jhfTc5kr4CBh59dLTjION0nnopeQFS66x3uqjiSI1pEy2guEzHX2ELm7XZWS
hLQ0onpKTZ1sNRQskbJ+uf26Axi50s9qJ0XXP0iTk7xGRFc9ja6K6nnfN+sy0B4tR9pRVrOkFENb
oKL9I+1WbQAoOJtwxFPs/XHYKWnkE2saolOpNMvisQF4jtqplOV0LLA4Su1nNKO1/CpEXH/D4rgb
e7VI7aRGnTW2KHij3Z31IV7eBXV9rtC5vZLDw723PCaUs7C5Jp3eflK7jqCM9RER2a4MmmKBg9GN
iGjB2d0pL4N3MbyIr5Left4oSlqcRGg85R8wOJ/TSzc0cnElM0WVnCmA7ALZWGpabw4uvqpi73CS
Tw7rQCPeBYMKr753VJ/shEFQ6nSUiExZcEq/rehwN+col+XdvK37Fe4qMsMGSgWaa+gwOr843M7C
YQQiBjMbeBJXxo94qnzVtERp101K2Mvtpbwel/Paf07ocFtdVCH7b/leyXuVsbdi4t6jlNE8ygQD
agbMG5E2B74DMl1NSXn3NjVHz/uhHSSvTHDbZrkgXe5jyMhb7J/WFR3l0W//ielxjRDdq4Uacd7w
AuuB8ovuyR8dSdPqbtOl13FCGWbFBsf+0i+7rJmcg8VphneJacbpPSOEm7tPzzum4GH4K4dv91Fh
s5rR0NTZZLN2+BHNdyZm4wkPSVZDDb963OYpqy3pG2d64rVh8icvM7WCSnJ1NZ0I2pGrWclQHjap
YpYpL1Gf5knwZzJvUBE2sFNVjNg3541eigHU+Y6VYXVcl4MsRlxJQ4Ctwej/N2nZQ2j8+wnLZDFs
ltv6iaz4aiUvYrRldtnYdgh5KOpzT4mJ+Xl1bZkHZWGPlnviTJ9t16uYbZkFrbV2l26eT/o9M4rr
/AYAcZKRXWNTw8zkVK5S2RSFPIwaoL9+LuTrNAaUf/9qyd/nj+plV39Idkc9CkTkuzyTH5bPvTWQ
iJIbb8xXHf3211Kbt28sS606lQRym1eG0OFSN2UsgNlRfnogOwyXPWyttcepPoOzzFARJn4oM9ot
oZi/P7j6O8VdYW2wa/STSuZ9+OfASO6vW91haEmIWw2GrT5NFLj44jPrFSVFEZUe3YQYzffLW9I8
OOUPSq4scvDOXPQJNcdYhevxH45kGvuO7YCFNK/RPnIJwKi/okEacJLyJh+BNl//cUqMbjU2ANOS
Gu8VV2zXyJGYKVKa8q4Aft0oco09JfFNcOLR4gWCbjTiYlMDwaze5ZuGYwkm7Nqy8SZWALq1EIh2
Q7dIbvr13eJJkDlfMl+nJUA3sOH2tohQZn+LeUkW3tYXi+Aw9GTBUA0X9VkMlu9AVn7UmlpQGukH
9vfXmLcPuU4FoqbPjU0BKsJoVbO2Ga0XT+r1AcldgsWxTDwWicPbYFkFOZ+9mc9pW3kCk+k/Qdwx
0A0FB8yTGjYjvcxGtt5oxk65NKBrN3Ba7oAdM19ZDE7M6+6MHVLsJ95UMQc5DX1mKxN+qzOGMbGd
claVl0uUjpAVW9eFF8bI2+HlI4xgMbEqRvzip+0GpyjNG7GHP+7MBhBbSJ7vhz2PbDo7rNMkhpkg
+lEzBhEx8yoBObRjkjrHATTXPo5beYBUk79T7Rq/xgxcufLiaNBnWCpYs47qQhW9umX22gt3Ix6x
y60iF4fphHgH7LiSU/Ymf4RKDqk6FuYx8cZTML92hT0Aan4Obsue6Z2nY8NU3jaiMhS4/xVy7y0e
wmMFcwhmA2FVfvFt3+XPpDgWvNxsTlFWoDud3TMQDXvkCG+4JurJZ/zTFACJzLE4VhEDRqwS21hW
hBrf/71LoJn6u42ZKWUAD8oOQogDsEw/EZEYQ8k3DMZtOQsnPI5OOkRxcom4p6174sldCCPIoTzd
2LRYOPs7PuXIAp4qdiPsxFwEZYmG0mvK6QtVMzhG9bp46YAJ53lEWyYV0hOchWmK/RK5pfvktFvs
iWi17GG7FPhzwp64IClFhB0Z2HUp2xbhEnL9GgeDRR9+h8Mdybz7pDXtuUGmyPqQXqyhR16qptB4
BIirA8WWzA30ssU0vkvPMJDcgSoE4iBc1PJETdR+XO4fLv0tknWYt9UvkPMFHcyybBjXLtZbK7zV
mI6tZGMuWo6hv1D3tjNNth7z6phpUmQgrkX1FKu0CbfnLLFCxqvBY4OGZM2v2pg/epjgTip8n5Rz
6Nv50RB/KFIScf29LOuDMgMyvJ8Uihk5Hfx5VJ9Jo97qssSZwIxBO/SZ3ZD/xgvrzgrluk2ygSxN
GKOe/zkilTGpBIWKE0e3R1yHmEyKQWIiveZ7g/conEr/CY799xowkNAq/z+Q0k1WB3BxY37V+8YR
ph5Y67zyfEzi2taNedZcbDe0dqJyGookFpvsnf+UGbtDQ84RHwTiRFehNSew+JvW8/tz/2JyUoFh
gqdQfzCRPHS+IjymQyylbYe2EsDEeNUaSqfmWjkg5KogySV1/4nslET3jJzaePnxnc/MUcDPlRRA
xZOnt6jND2vb58vdf3SGxiDm16sGZTpDhuuBwLS8TtwT2w3ye2xNvfjKtoTO5tVc0IgfSRM8N6kd
M1gZoFBw3uyPE9eGqj4qpcQddszTuM86y0J1CLZiIQPhyujtvRBTQUSGbazvDQS5iycbRWEbJ4Hk
shouRWlcM5Svg2k/ltYCcPvGfSODUmMZCla0+YuqBSGfozFLtyJk5cOzbPcQwn5ftgYEh32SOHlm
dgfBPx3wT2dpeoOJjVi+9Av2Z08rkbB2rVaKgo3yOSpLpWF93KUcMIxJIZKFNeRlxxts4zN5GRSO
Q1sxkWz7I7wGQRUgGib+WUigSPJFGRVTCrbjaGz4yfvcIAD3AI/B2OEvStr4Cn5XjRK+jSjzGhbV
uhax2+zZq3KBc3sHRgG9OxrW+PUYOAUzmWTw8Niu3wiDyefOhrk3GvLovOV0h5pea5XGHjjzIBRy
GgzkdfUKr5kAOsRPgobaeo21dVHozTs6kYFeR8Utgz3L2nO59eIpZsoqwfwAcnbH4M/Yj8qqfOgd
SqxXhkklEngmFMN5dviCILHQNuI96CQyLuKanSxBwCz2FWqXVrlIfxg2teHRCdhqabp+NbHtJizs
VNPXgWs9QHYDKgKe3MpNN1zzpkszq+7eiq3EqNYKBk0g9B6xWS9dtmcHMIaVhE8DSUNFgsSTEd3/
27q5i1QDsof3Qn0Hms2uPRZeyl2xjwHXkUhw6iExi5vlzqwv3a9jM9jzcnpKXBCLFV1UOh7xz5YX
aWFEwbgR4bClbHEmZP2bLgOcJPEv7Y13bvTuzQ7QrIKcD/hri5WhHWy8ih4E05GhxDM+OnSAHIcL
Wqm3DLnuhHXKzQZPmk5XXQL64dUiC13kmR6508Pj5Qg40gv883Ee8NDg1SP1f+hyJ9vU5/AwsehB
nW9voj1GWHlu3JgHR2U+SBjna4h8QZFsZLK7nDqyRw5Ka+9yGo2yegtNAquwvD+IUyi1ymHVrTJ8
Z3iCkkI3MlNv51opoJaLSWphMzZbKQk+VFZt/wtIz32fqLFBvg8AdnSLumodw2bbF+X0K1UrEEKQ
6ZKXZDjYtvomZzqCmG57J0QMTeJYA2yywdRYuFW+VeSw6ks2XZM4uMbRJgOkkTTcHAB0bce/lsPg
si8Toyse56PZuEojiSRWbkhJWT5vX0P8/DWSCP9+4Gwu3wI+Hx6r5JmeRYeHdupQooaDyraeOm+j
YzCIV/OztERIdpS+4nvWq+2MtS5b0bgpW5T4konZlC/IEKRi2eFSk0P+eGa3KfB20yYK7nWrS69E
pOczYRYbyyww+w0OQXT2qEySRRkkGgHTna6RZ6S/Z5BB/V6PkQkwN2HchXRBR6QA8jQFI6EuGdX8
omz2Ptv4EyQLNWL2rhxeVXGNlke5Rk6jD4C4KvcxXGnSGEQ+/fHlqKvqIL0tyVS7eV0SfFJwGA5s
OlLIAQ8U/FEhVkhuRRVFrPBsMfgv6jd5U9NznkgmqYqhl/QDpKRC3JGIoDXvu0LOhyJWtL6GVRWp
j3TZSlgXWoT/JOVFRNPPtnTx5GPiyUrjPtUKLyiJ6U4rUqFgT3e/iZy3v90yvX0QXUQ5Got97A9U
MPpfxFDw+p1rRI4mruSknopT9i0oMtVrBcCxd5cf2JbY0zl70wpeekJGglh2uyKD/NQZx61Nlcts
QDJCP90NcZakh0VVQYaQPc/CZsxVABbwvnRdQDaQ1XwpALm0vVGnvkTFWOgwTXwE6XsY0H3e5W6r
pc/fJqzDpbI4Hmqc6N2K/EBXDRLjdCwEuWD4OdzTevabxnmC948nzp3fyjrkfy8e4YiH7vZL+793
iNwY8PRR1zdi699dZ6X+fKRvfE4P/okqPxXgVJJyQ/EjnKa7jfY6DrlyqO7iLYQmPDqC+7vJa7xt
6hXf4lIrP+bH/O/u/mrA6Iqn3rGLb8r+kq1R3tvMFSrYlW+niTmjiwr494BXYTBc0JVivKAx9cGa
9JivYtchb+MwObXur2qwrKYkLpIbQU38NykCpGZrKAp0yyNc4GCK82z0G3P6lUdlPepoO0fUWSqc
XxhPxaqJj+52TFOQZ4eSDNYmFAks1lcsi58BhkkEet2mIS2xnsRjXKKJNXWtAdw14M/pDkxHkxBO
6vtH85Pm9IDBff5WuV69Jjje9asynEAr2RWI1OY5T47hSXeuZVVAlX6EEcBA2Rz8J4mwItQbOZ9o
TEspv4CGqLQ0loQATHBBc/UK75fcNWBvEZdawtmzUfx4tiEpT29Uvm0jTq17MTxhCPqwzq4J/Adx
hyY9GceQVvQ6dxj5Pgo/e4UzJWgjtS9c1Y3sjfjXILVT11CLm/etLSWqmqyOLc9gMFT9VIbSDi1I
pfWto8KvtDdpwdpr61C4UMOf4yOqJ+jztuoqDLpkm260egvj8WFZ7U5aISWRvmsWB4y+DCTCJ4eI
lCJOQfNwkatnRXxjrFXZbSqq9nr7AMII7p14O4lYdkND+uaiZEZiiFC9xnp9rFfmj+xihefKNI5r
2e5pjmGXbc32RdJr+rVs2+G9UMBkMC7a9wA9PQNeLZpoMmexsauSlmlq8o0dKLcCZE5YGhMzVbYS
b5BqavfdCtQSBgM6bnn51BhaqbN9fMtVxERyEif5vCe0PNXgydvxlmyqR/rXS6bH7HDAUHvQi1s+
48w+if2DPKWxYJm9w2Npjo5ZYln3dY01kt4Dg6mFb8W81z6P+tQbHVbiHPVDB9JOSjNhnDsSewNp
a4PAWRIlQXUv23qCL35rgtXFX0XSUKZ90dvADuLQ95nkmNzp2t0ULMRdGCSJjon3Pz0hXIrC80kP
Hl950HRgPnd6RzE6Izmk3zUOv3Jb4f3eE1y+VV+87KwxFReAr5FNAToz1rlzrT5IdsSbyFlkxCn+
MJm+p4XY1coakk76TaWosXZwNnVDG8KQYW5XhbtqVxLnNcHwsFFheVh9k1qo38Kue/wKTdq+Lh98
U+LtdoxzY2PIibuRea1PTIN6I4duu9XqcQ1lnYLWWiPVyUUyu83MeFUXYAATvTSIS1JghCWcAvbv
owt1eDSQCqwvhROpfhjUTE+MVxylr9TZXQ+7hra99JnJPJgY0XiZgaVNPfvt/Pz5ZQ2f+H+vvrUE
A2M1MZ8VkMXo3yPh6FX5KHNr4MA8kBvhmqCmSDmpjWnaKFlUBfcxTJol0G7x8CBXg3oQ3u3XkoAW
m6iZpc6ao7SsUxQv2iiCWQSZ0ymxoFM7Jqli/8X21EXsH+taoZe+1vtgW3XbvPMHd6ciNL8nc5hT
a5XA5G4COw6jjdjqfhHdAaqcpKUseDCuxWz+aUE3W640x+HzBQKBQJ69lxXA/5mr0R0q7fWhf0ku
+ZB3sCKlpHiNLMlCWhVONC3ZHbJE60R5MUC7ehZ8xGOiSGR7GDKUEbZEcjEWaU94ZPHuxH8YVRqz
8fJRTmdaVgANpVdfyjbzCZs+KRkfgBTPM4UMC5mp592vu4CMHicXjBToDp7flBeitn6lmJdBIdgj
/0i4AbT2veVNUPYz/m8xWbuAInY4d47iJJtCIu7GrTn7x9qU2tYgYUw2Ki5Wf/cu5AIBrdrIgPN9
zdATI7PPDN51sjG/U8PD3bJOtfy0491JGMZZGOGpxj9YbCM4MGDi3Ehy5tin5IgIo/q/i5PI969j
INYyCnoEMJ4npvOGywjfQWc4lqwpbR5JkT5yRNI3Jqj8moFIlOOjnnOVpUxWg00nEaEZrj9rsEn1
7Ro2I6ZRMK2nkktS0uYQooOepZGTPn3FbVfvwlS9c/8Pnz+pV3f9IO3utoduDJzGm/8fFBBMbkGO
H1SUCK+tANM77z9+NqDhqjV1CHEO+qbGXU1FiDtLgUYodUdq4MdEgQuXLdV3D4chnxcR/ts0gaO+
wivw1OZlVKftU9/W2Q0Cm0NTzygtXsE6Lrj4oGTDgbxj5JDrWeh9wjyZwCXOMi2ZmRqMbxZ8DmpD
Q8Oth12FquC3rm8CIS0kU9ldspropw4ttG88y+v246AXBn0paglqjX5ntvRBCuUsHd/D+kRCv9QT
+B/sB1H9yXWIgNnTChRjWA9dktJhprOpbWjEqB5kBcx/5ubHr/q5Tljcko58dIZCTP3OpAMZsxNE
XY7NInM7oMv7w8PK3ynl2jZh5iE3R5aaUEp4obaut+rvFd04rchxsRrh3xdt/NwhUZ9Q10K+Onte
xchIM5R4ZJ3zjwf06uP0hhf2FLUHEATbEVQKhKhq/LqT0nXb8hCMOCoGuRvyZDI/lpLaRpIGDjS/
PVhcMdY6hqLzC0fh5tZdbZbnf9R5OsWmFW0RaAj2o8VroJyYqgH7J9UYmC8h4aeDJrt0Wt9mX56u
a7yidIbw8yy1mG6xm2AuEVLTAFsPIXTjIz4cGa/5tc0SjLB4M8LEDeEpq9kdOKXKR6qXkbn0Xd3F
UDgvjJTUiUCI4en1FgCajpqHrGppTclfENhCB0HHJI6zSiq2eABlp7TXvBHLj8kCm2nJf599c5GQ
lziNINafkbOBcyv8qBO794vyUJitb0x+Z1XFfzBFX2fBxPrUuL8PlYaMlxAeYyjeDVsZYqxjSdTF
ekUrvcDCWoYcDbmwt9YD8XdmrI7/LDK16hwcHi2GOskePBCXwu5AvhOlZ2OYI6yCFJ7NFXH5zt9L
7wZQrFS5wCBl3JmcKjH3s52MHfUAP2DVB5KI+5Qki54hTvmpVuY7ADsv9k3CwGbZ6j+isU3MArNL
YkqAVMuxDDUfgroo6exh5IL3xoO/siGwz8x9x0L5Gmg/K96kDN0GuBsUlhwn5qV22RPzQnmOuJYm
KQrOkI8VzlL5z12mg3BVeN8quA+ZPJAdd1H7U70MIh5d5mKiv2wvMt+YLwUhHf2kx8F+S96IbE+q
FmZNQEZ8omVc7NWEvOWoH0ZU5kIVWIW91sd52jXo7G5GWTcMuw7I7gTZ/9omzjp3nPOwdtSU/Tu6
7/RwXqmV9G5IZHJLsAbzg4xInD7uZOd/tGVziOvzRcDTfIzRwmSHL7vGHLLEaz2Q8qMkossTcjmz
N6kTx+lfMMcn50JSSYsA7/z1d37dplKvvJ9wySO5vFN4yBAiCMiu8M3tHZcQNK0DfxULiDW8qFlU
5qF15EoWDETruPtctKTFCsaXaI6lnrQsCLs20p65GY6fnBrioiQhwRcievIRdNUGSK7xMPP8Sp9V
uoaBoFPGw4iMxSbblSATC2WQ1SJok75E4wmSIjnol717Isw0JL+WOQrjdn8s6i0vpL9Ma5vJRDD8
bRn9xAuGm4nsFEpBskv9GBU5HGzC3XS6CYsC6NSjFs9II7VWus5Jxd9dqsxW5gSrJLKUpPTw8/Rs
YdZeHGmRejjjEaBqJArHEOonosM1nPnCyr9BxiV9lHFMHTQBTBPSSrzEZPbwPw4gDEJjZsfwdkIy
kXVfUTzDaUzMAhOlkiW21oriZiU14gJG4wMvE9zO2TL1Z9viyn1GpFaUf0kPwxsYarsnc0GVmBCk
ik9ZaSCx5OIoM0PjbxKxDdKSPUYIVvvUFNcu2gtevRR7EWQn/xeXVEMB9ANFv+Hakm63kZ5V2vpC
kgNorcUbk2lOvPbVzEVFSQU18ZKOuML3Fz7s6i4ByGeKhrEHw591xqf4zlitzJCnJLmk1pOTY7d4
axbBYasuzjMNgebEkMR7yxPLSe87bSmB9cwASZYtSKaqMZZzeoF5jlA1J8p3h7urVgPLSXhYql90
Dxxj5othcmfBoc8uRGAdLIRWu+lTpZo7WwWMghvoHEgFkKUxF9ygw4HOLGkH9fFfs8/eewwWS2nw
HBXcARdcdoUD3wgvSaNruQARc1jc2vGvAo9mxCxuPt0JwumsEeAM43CvUZvqB1iWnPaqK0A9QbHH
+36V3moWD9zutrfZ8v+s/YiBxBFDlY36XompGCIY7BnnVrV0xyM6YMX1rkT/QSLlIqYNwEtEJYYC
NHKnWQek6lalVCRa9EMH/w3K7BQMga0ka4QfTUBkynMrh+cXwrz9t7RSNKE2kzJ4yjdzg14Y8chG
/cuCgWOe2a6e4oZ5Ap21UHMQxDqaLG/s2/sdzeWX2dLiTz9WYPwxuHfS9ehsiz5f8eCEXBQcBgXA
p09z/CdPJ934sv7x+Ye9j7QxAgCQVOgFtypvIMKLufvYnNWSQTURiM1+Jed+/+zGkWz05wdmfX1h
Gh72u90rb7KJVTdwF5vNgD4abEk8KqBiRmcL2LEql7qda0QDkxpucjD3/y3tu/LDkruu1TRj3/eE
NfQcTy36l1GizNqtLdvY4SuXplDa3XN2eGQBNyJAw82xs4JuQ0F4eC3WtD8py/ltew2FEg5YKELl
Br2g1GUm6kE2zIq2t7HIV/8Em7P5RyP0U5h1pkT3cGywmHprPqPW+8QWVO+oTTLNzzmEVUhFcTP5
m7tMD4VaJcALwPoZFUHNltpHEZK174kmTBUdZ1kfsxPCdTFhfriakHobEbMy6h/zjwDmKpZbx1g4
Oi6K/798L3SgWQMhgzdwlmUcB/KR/AeWLn2JRSdmMWizzLNganjCx4dTxvSyBbpCaBc8slkyG+zW
j4bqjIU7P2Whick5XG1cOQEabWpd0kPjlZk9AWjds2xU11LKe6M4YWJgW4LxmWSJrypQGt84w3Vp
ypp2m2DNorxQy8P69/ZxsM77A+6VIwzFSlGcEa2BOxIn0I8Yq3rc0GZOPekgFfUB2zrGOWbfQVmc
jPGPaEbCVzOcluWkOT3HcxVmSecxTWnDTzFlzHf8xyBNd3HNxGUIbXtlb8RTqHqpwQgGtKDT1R1y
bGketGfop7LyrvB+UJBLdsLHNS8cMMlsfSaSh4amSl9xHCcEhmuV3Nl/uruLvewXxbbQQuit8y8F
hqN0s4rn83BUNfF/YC87P1LyYg6Gfd66BUC0yRw2qyTJy/lOkrAmzTTkxaqfBN2Ba1puOryEouQI
wrB32WfblnyVr4JHsZh+jrCAwTYvsm2w4bHPGnv9flZirPXIR0ZVv8zNMj7daAYQnfrV4R6g4ZpA
4PyX4n/YJJKY2H24Bp7G7FWRP2dKTD1FiwyhP+gwUua0i3EMHyQeROPYcw/LY0IGvYr6RzfuSNtj
1UyuG0S3mt3BEZz3JvlWX7ZT5358qR3ulauHcSrd5M10/CTLIaRx0uwWqBLawR5Nrae7Va00HHZS
g/JlKs9H+fl4gr0soudqXio+dsl25KQCzNzhFH+7jBYgcDQIej9MBjr9XV9yq/KfX/7gCwSVizju
vcrtEN/2a8vkniX8VmN1h/1EgR/aN59xIBYP8BQMwG9q1EBzqhbDy/dKOb61OWwad0d8FTIdTf28
w5YzFfPq2YZPrYy9DTAeR9RnO5d8LOR6Ky2iXl/tgHcYdkkblnC5515UtMcWj9t6p7PlXPVSEGoy
qdMFxiRi/QjHDCxPQPbeNgDWkfYDb6e4RyBekvISmplo9hyfwFToGTzbV+y1Jttwf0zPueRx3hYS
2eB348uboR7RnCiwvWZY4Ph4xXP7rEgp19VANZXjIf+naAFNwqKBu6/F3uRkiAFv4YV765piMcxp
n1qAAzsdKYE4xxRb52Ot0COojC45HAhE9LjdIXxViGVa86JFKIsSsOfVjsKOwwFp/RucJvDeUsrR
wqvXU+B7C7Z+QBtEcHCnQKso06xvWKwdfnbumvMqAbr6OPYtBJVnj5EPI8ReLuWSfP1dpO9/mCst
iUdALeXStWmWsvBYlv3tzxiAXSkjZcfdGFHydtB0MEeIVvGeEzrdsfGx+AJOjsSmdJkPt5uMgksE
kcstLZVU6zOa+vZj9WNKLf9wI/TvYDJq/r1QrCryFhgGHgrX0Wl/c4tNDYeeqY3VPTMnyCwq78IY
B0WiAjRsnHiFGqRKOWzoyNQTv69uyM77GigocSFp5XpEoBVzvq/NvHCP/iCol+i/7WQFOOizY8xs
FC/wxlOkZeawn0Q9oad/56Ujz2Irf4Bntj4zI2zZCH27rlMT/YbCvsR5pbPyRFnzLK5/VBgHLgEQ
n0omQd1oqgLttLXmnPN3+22SzyeKNUcIiKtYd9mhAU1wSrwvzvc0JDzvaX/FE8E3jgsHON3/i0ho
PFTbRJrOO5uYkevn8cipqj5GeXLTsQsUl6HpqW5O61scRslqwj9Z7lSoIQhp96zTRJIx2gFihsox
iKIlznqm3A5Lt8j2T1jA4CxngDVdjj275O6vo8+ZsB3dNLaBZhD+Xl6VDAszjELTyim8RtlyNTNe
88TY3imW+PGTsBKj8IffahYy5UWigO51PbKCnq55DtZQ1gYWqQSzSoS4N7SbO+QK12n5hCRIttOF
CiOXca0AMxqZfPAWX1hDIIUfUyclMHacfLcrv1y3N4XxU6rSE/Z7MoCMM1Yk5GJYI1e3f2eUNNzK
8dDhVLO7X+63jJRlXPc/YoRdtPpT4pTC2+PJCxVjk5cEUIuL3zQ6qzUKv/CmrOW5BfNiF4HTUlTl
KJbBnbCuJfL3j0Z/Ey+Sjtq11IYJGVUK538cTB+wxlJjJnDxhGQ1+OqHy1tGko+O6hxSN7210do2
FTjpSPLJ7N6Tc277xlDCWiylXo+7rMokq8MgY2c0XYRd65LKC28UBSILK1bdzczMgIwm5gWftJTY
0AuqYl6VCCuqKNQfNIjdkLDbg2iXc475hkKgd8fTyl2RQAXSefjkaJpHXcs20pq5TO3g64lw4Ojb
Sn7hDC2hYZNof38+EG5OSdn74KSIvEFTA/6g2ZlBWW4xkSh8kJK2/D29cZVvcbABTKVNggQMAz2S
fN8Gqo/rFj25a+hkj1Ev5MQhanm4pIwaBq6O7CLi5WgoWax5YlUidlT8tTOMbojVxP9K9+bAo8Mu
bjkzB/1TnbswvBm7ZZBSeUcoJsMMvsklKTxYmrDib+oj0O+7FgwbYlBBVbjhXOdTVwY23YooLGGR
H7jnVlghcCsB1PNZmrTN6lT68VWeZBCALKqm86kNytlbN5Yeewfc0Y9KCYREaIFqdgAMJHl4w1f7
ixJZ7b1/Wzl4e98b+/P2zNWPjwUsPARuzz2ESFHSnSIP82GKiMOhufMhyNOmTzjRr87Uib55UlXT
QPHPZepedEzZo09o0SuAFlooUJRpIqllJmNIp0VUAHCsAneG/FZDmKmchYtt7ZFQdBEgtMKvBXKU
ZhiymHpQB4s7F1mjxnt5bTFkdfBaNUYxNNhBHfN/KbrvO/JTJIyIFvO0Hz88Cu4jjPis9jIXzL53
AwGQJj+f4fmG+LjYMTpve9BLDZScnfZ56ARR2UwyFl/SYNzwswkXe23kck0vmXzdFlV35N28dPvW
KJtZty62VK/FlqF2j9glITgmqH2b/MlyOyMKe3C1P8I3Kx0ek0zUZK+bhzaMjQdk/7ggJczP67kJ
ySyzKAoij8UXALfkbHP/7lLBUFtoZGKWQr4JCsxfOGO8KHigCXRzvaWWgis+kY9GgE59CyBf+Zro
LrcSVNQGwSGKFQJlEPlLXO72QwiRaklR5qn+K9w/riMZr8w9ugMcoWRX8Yw81QU2Mgehv9Ub26C/
y43bKbv6a4ET3SiH3Ef8A3YLBBUlP2J2OXEtLzUWBXXU0eZCFgx1ZuR4I90YCGdR8m7ZfSdYNfAP
dVzX6mFAXF+r8iFHhf/zaJIsgJzbOOrx7kN54QbRmOyEJMLRBX9LCgXfhAgZkBsYSj2S2SS/QeXf
lU5i1vqOUyDA54fPVKMzkfAkt5QBG2Ey1FLuHqWYHmWvnjWErgGcM2WDlAirM3w1+Avd4qzJeS1Y
BjPSD4rMEcpFEuCGlzMJ9h7CtJf2MOVOl0J8T1iM/TuDpTqvz95wl0BtU71l76/dRszSaXibH4HT
lQeI/F2qUuaHQHau8IjNYtT2rgK2XC9NJ6ndaF2II79pUDYyW2jxQZbpmvE7fctP2Dj6UQtfPi25
8N0s7z9KeLNBlxpw2+eJ9p+0CWoQw5kq4Zr+LJmJ8TvJ9sCBaSmi1jLUZoqnfAVGYWOVDrSTORab
M/3kiaUbSReUgLukLy3C4jsn6UsdOXWReI8y+3bpfLnHr/x/FkRNEyEUUvw0Xp3s7bZGAgZAOBTf
Y8jtSzISqSXqJzfTfZ6hAUobbLANI4uh4vm0xlq1fHGEm7zZ+I7X9r48ryss7RRPpo/tKn4c7ymO
Vg6a2Eqtb9Al/nI4I3OPnKvMJSjP8yPbvNicXq63kkC4oVvTf2zh3s2pGlaMjzqot4FitqDt+of1
zOGzNq92mmCCR80rdxo7H16UFSrylS8gc94E7mfteGOUMakZItbwIr+xNOamtMji/KsMyAG1h1yf
3LrrAEJZBQFa/q+YNbJQMqQhzDmV709Z2hkANHBJVbyO7cYRmnrT9S9Kc9PFE60mG8BmnuzSXvdz
1K3AmvSbZQCI2tccVeXVJxHvMcHoFu/YnWhSk7aIloxN2GZKd5/yV22mCtnT4QPfSUgWk3sjiv2T
AwRTDqh5ADEBaUsplkTGhek+Kug2b/fdbPpjzPerRi0Zk4I2uLguLJJwA3MnHRyNzkLun8MVN14j
S+dDuZU2eezMg2E6V+ux2p6lyXr1pPkMVJ9S0ixOJicm97jGuTlYNMzopUW5OTofa6CHoNdy5KMU
Uat7F0XIWnWxb9N3vxTBq/KNTxuexiiLbsjjL3Ekyb8DknM4YMhGKOT/F4Zy26dZASL2jzu2PkXI
XdlmVtXe6FDrRCGHm34f64OdEk19SLgzFQS+qo3xkiLrOmqCgSGi9yNxOMkKG/qmVQ8AC0YRy6Af
0stqGw8rMjO3DZLmg192LGbaYgKdzgjvTEIloWad+4ROeVUUEyj7b6ER2DucmpfjSXmXXM/moRh3
bltiNPhoU3Z/mZdpPhjt+4OVq5HxSlWAO3Tn+6GY+mwcY7DwtgaQ3Arebftzwvmm6lGNe62yONyO
vrlpXbzT4/XpAHLGh5yGUIYoFrn+q//cOIn2Cfi/nqTh+QCPhp++UinUnBCUlcHuIC+88N9gT1ML
333IaR50CIG3SsSpKXY9OKQ8A3QogAtPGkGkH5yxsF/BbPhLtbOhnA0rbmCUG7wjwDVeV5lHo/D4
U4zt9M9MSEqY1TqP0c4eG2Ks1eL1ffsY29n74sN3l9XtUEscqSgVgjkmD7rsaOjGl+r7+LZaRaTD
EeSE8N14RvC1q8ORXFDWxBu6HyoWBuSpbs5UK3NILwgJquNoSXSr2CkIkLxXNV+na+HlZi2TlltV
2RG9M0qiRoXVZMiZXLbKSQbcuXT9EnVaY96glBzS93Suny6FWPnpEow7PWQTohwuX10jBipPxNZd
a7VfU5F/H1KN6OASxpLA9hhyTa9v6b9H1tqP7hM0oFallI1TQU9qWGakm8H5Xfb0K6dj5wkTFQ41
bu3sQAm8b9X6uz8ZwrphzzATaIl/NUcXmd0lQ06V3MhkRv8iP0vt+4T6x8Z9FGx1oyAVPwKirb42
vbMVhR5RqYF6ifmfNld8QsWJYBuRoGAEtEw6ww3rEQC7omvyTi8D/P2J5a/w3KzJB1P2p1LxYWk+
gIHC0wztH5eUDsVPRcQedQjNpq3Bsrs70LtcxSCfJLVQt0tDEFE3j+mbQ/nwu7DTKvDhQdhSJk6F
uOXbkYEKs0CmMs55im/m6Cs+CSsedQ4tA6p5YAsiYHjG/s6WEoIb0YHMNlMzKyJTo8VX6v7InNXg
kqVRMTsF4ic5hCihIubiUThHkYlssSU7C2ru97CDHRHaTUDO8/IMf3Cv8Lvq3S+il4QAYNm3T1lc
zNtfQhq7VcgAr2JvDEmLh8Cu9Jz4kEU7lcy5+IdVrc1Tz4CGSG3b3hlVhrgtukROMDaI+eMpRexk
u0yC/wVabCRTqCq68ZSACDXr17A/rhToGC6h/h+7WGK7nok6Kiam3eGun+mePisBgFb2PcFyPXk6
ObJZkJxed8XNX3flf4KW6OU84NaDfIe1FVpHLWs06O35CvkohiP/Vk78wBuq372NVexDjHR6ro7W
BjrCTn8CMzK0aFoFm3N7KtGdzXFTwOduekiKpu8UmCyj/CrNeTop2Gsw3SrEyay2HdQlRKeReYo7
Nn4vCdkMgGU506y+O7Z70Z6S6NEqXqeQD+JDfID7iYxa+F194Tu44CsLWjf1aht0TOZwKJXlMBG6
M4f4TEPtgQdFwaqBaWK4WwdOx4lcCXQIXRiH/3hfdJqJdwb1C4nOtUQ4fIJd44xs1FThrV8ll9oj
hFW4q07jTVW9yjA+zB/35wB4Pf7l0b0xyX+//KEZNV4OSSKAF8gNb3sdsK5fYBnRNVazGGDo3tnq
Y5kpkjUGIhHWvHtqDmaJ3roS2PFGui7595fruxVjeOxUp62PykVh9e10JsI2qhiWheKscnvVHyel
i9kAQo9+1vAhREMJ8m33dtlCxqQZBShNDOi+uA1hP+tapSiolqAcE1k2e3Fhi/YBsbvUZQNulh71
+NekcMPy8dqCthYyKWqFIXkMdNm/4o+8oYiCSnmKLlngZRVRMWczd5Or3nKjTaB4oihULYPtLYP+
clRy4cJb4eKIBdttMPPc6a6UlrTH5ifGgjpGt5XchjSU81XfzLs6FNeamrKOkkHXiZbuGomCAwZ8
J+5AUi5T3+LL1JzyOOdmivt0BtLEp9jh8S+yBhozsxQmnS0aZxtcYZtcxJMgDP2P4d7LcOBeiMe4
N/AiKOdYF/0AjsuT8Sb7ExlxxRDyiZM6RxXacDblJUFVvYA40SccR7ZD4I2UXLKhiU69ZSe3+wyt
wcE/l2yZnVrGI2yxcHdMh9rnSTsTFyE94gHBLug/21DZEzOphGInsA33wrnRBg5q9b8Rbg8Modf/
1vp6mLMgWVyklPekZG9TL1qOSVlKt9AHJEZS20KzPyFXSuQfHyPl38xb4R+7+8AF+uouO+w9SEiB
IGyj8DMA9Wq34U1XkUZ+ClZZO7WAo6JybXngoV1LI3W4g7iWVrisCqePVbGqaX/kZW+RtyK358wr
U5JNMhWaHjUgSRBcusgC/auceGhanPfupVRUr2bWyPKbDivaDN/4TOY1FI1RK3JI5i+t0rDmvALV
Sq9KLYKhbg79nV6ZvciJZ0JT5+QJujXoX+EqiL0U4SMd083b+oXzgPCqDug01q1RlKxkZH+r5j5x
jacTlLwyT87zMLu0sLp51znQ9336vxzPEzaZvVOEjdSMXa2VCc8IRbXdsCeIyAas5MmXvcbs59Oe
bOAXYFhosRWVN84W9OlSQYA7saIBI4j9VNR2J4rmjg9KMWUlcATLAR/DVZxhbVVHKQ3KH3lQ+jLI
EnwqJfy033RfLpfTSCJM9t498I87Sa9CrBfofxtIGmUM0bWmFxzJrlLIiO154TEaBq/KXoVNL8xf
wGW4sH77uLwzSgbWgla9KH9+IN8uTMw2CXa4jvY5CX6ixLYhF7JGtF0fhAGbrC1ahdDd4rEgV4Lx
LFJCD99JJbLLdNwnPm4/Q895SMoc9NlLhUvbsqT+RElQY3WCVQKhiwWdMXy0PUvyWkbm/rGgxUW6
8yx8WA4nVf+91VApjue/6Rlp+PZKusqTQDb2s+2BEcBv0MqNCQjdti4cs0o/l36ITR4axJ3aMooF
pYTOtLmXpGRiWEQI53jMztpUtL0LpAEyvaKiG8DWtZo9BZgdChVkZ/ZYh91Y+wRi5tiDTP4Kxz28
TxiWByZ5G2qyVmt/zZDoEAi90uCx53tAl1Xzr7zinUY1zAgR6Pj5t/2oaIsGCOWAXmc9arvNEr3z
cCYm23g3dGAbXi1C7rhp/lXRKzqrk5lPF0Lnc36VJEWsPgKF5NfXKON0RwZiaH62Af/pMN7B1/dC
Kku1MOxl8pumdsLQf5RouY35xAnoMY4p8PxWMdxsSfNDxbW7FLKvWxj2RctyW1jqgZ8bCgQYMXgQ
u9Pmw4eCfVzYu61Ae4tpBfSH06dwQg8bauCgbs6A6advMV83rPehaE82nTIzLJBHho8mxSaVnKyN
dDu8PyVTsKZW/HrLNRdBgMUXSbfL2NnzALKZk3jx4k4UFosdjsVk70IW9PmgrRO6hL4kXY+9q4PD
yIpskb5Avc7221lx4vmE5WvOqtBvI2KPb7w+SQ2F4mWETh4NTzGKZHMVPhA52baL3+Ajgvw4/i6u
jZIINm5P4sfC4rmFZMNFL6kRScz0UDApalKiFCYwzj7l4boCPLc7gTyFNSuTBzseGHssGB+J3Fpr
qEc7ZJiemuJHlvzR2oAt91f/srR0LrkLs2q0HRDoVNNZE7iJShT8D53LY8+Tc4QqBOCLNrQAwHiN
afnB7cRaprHU2955/tIsqL9uYTyBcb7qAPxnV/gE3wNj3yVJEOc/bzdvdBfYMdwwjRzipZ4t7gdY
0tN4JViPc1n1kACqwuHf0FS0EWjwnSDlHIpKerqroVhRAIZfl1zft1rQ+zMu7nhufgfT9Pa6m8oF
OLbhce+Dq9q6f9pLWXvJC5FIH7mQbJrYYn3m6Bfa5IOUjFF+cEEjRP0eL5k3QuRcogFjxpHm17vA
FgC3zlwDGnVmOdJLc7yPC/NjFYY6ficQATIsndirMNg/GMOON6g2puQFt7KRDdGw4d52snuA+L9g
33sYlCXtR32ass1W5epzpx7nFi0F/H1Pw/YW1Vr0lUxWiqDMskZ98OgxtQMT/SxSaIM4F4VuUFt9
TPGFRMfOQ9JPJ4U4fXjnf1kMoUD81cjaRuJMLQBptiJO+XnJg/jzA+FpLOB8P10UPJGCk/Aog/SW
8E8sHtS9dbhjAHKyntwMD1oRBvr6IajlUcsyuxPCnyXBd4ej6pG39iVnguzlwggLLKibFQ0zuZoi
McDfJ4SQAg8mgJQ1LOrcLIndat9Pq6fT9fWusHhee1/HhbPoC9rr2KAkbJMnhLfF5u6uDJfl9/Dh
NUIGaYPo2a2yhVWvJh60YDruwuHaOqpfGAFL0fDA9kbK/smubLDr1lsEgni0oXQHG+ypBU3XNYGk
BgGq2JnShdKU/ICqJrR833WPSqQ8BXbTG1+LaqLu7SsytBMKV7F0juQTgcgutndGaAWEevZnS7Vw
OiGC2kZSCQaXJ5P6CfsZZpFkqapnwPeh/zCNh0QfZd5D/tVDnTXDl8I0IFevq5nA+5132xlglfaH
E9AGgRVM1GK7sUTVcM6DhTLtoJkkAkfuG/hb8k7/8KhaT8NwVo9rQrarWiUntx4MZqHOLXoEIGut
cIo3uUruiWiufJANCp2iV7KIjEmH9OWdx+vRlRpGeXNPlLiNL7YkIKoi8tVvArFUxTlTqHbjN+Ui
syI42RsXETJ1ob/6kyDPuJD/oU/GJL6OZZcRmCTZ7EhWyWYsHtW+VKJUo39gQ8OmVHMKCjaoaxXN
oNuOOG3TTc3GEU5Pf/8bSz4HCfAKQ57nQIOnXD+Pg0lZFlg6ew3PSh+Km0sJj5/OUuRX9g+cslGj
0YYuAneszzjSHhCe2nw0rpfZHivoA7Kaszuk6cdsDATaxR6HsuhsWV3K+oV0gAfarvhmH2uUIpYk
xBCXiqI0Gy1ob5HAsUsPq6zkzeqC0WoN/NMKQHp1YeY6c7P/Ttv4EZl91lnKDvcdS1voysWcw2Ea
GznrH9ceatzSaRinmsuBHj9VZ1FhpU/4Yfgf63jcyOmz/1hMFeawD5HivisgkQHY1AZKnRnGyVin
JbMSgRWIz9kobYW8WQ6wCVqup6FCXwsLgWQ8z/ryGUcPn/HtH3jQOXVjM5gsz86FrnqWxNOi97yK
dD5RYgx9+VNK9hxFe3tAAzmi5hlA67Qk72k9NBTRqpBkfvDBUZjf8qYTvJ3L1iSoquVMt3VHotJl
FgAtfStKt7QqHKEpiyYFv1ZDpQvkl/cHPFGVORQbnJA7yzEU0EJWEEj+D9JiovHIMB8i51kWRF8Q
vIIh9VzjrXf5H/5OyhuVF9eaTn0jkwtUeDTFYrPU9CZLxXIqagNFvkApHK0N+s2QLDjUd9cGQrrr
nGk9h1Z3p2ETCCnpArrqwi/+SMCRjEMPhOAHfZ/BSZXH7qDJnKMl+PJcYeU9CmEv5K+dabrUs/pA
EDZ1IP3GmNT0xjQVgKo12npsC+nz6NHcCm93qmar9Tm/Mzr8u2AjUG3nCXNfbN5NxSsM/etPxuFd
RvG3RnKEcm8VuluM3LAnSxVxDOQmz7s7cYyST/kaPdUbeoE2iCbaTANGRlhLN/gupFJb2NNkq4Bg
sgRoREHfexa6pFV2U7oF3PyEkqyszhWwa390R1OKwWlPnzAGqvr23ur5g191m1lgYa77nIrbj7P4
8ga00iZLwPymcDaUFgXb6HpZ0XvsBAxUqbHY6qmVan6wtMAphQd3InNTPCYG+h/pyypIyX+ZE4/J
rOI3+zgJURbBBKWNvRbRHXOLzVegI6pUhCXwXPKTRab/dEvbDSkvyH/dxsi2P6MBW4p2z8hnIETZ
tzFlLRmUfu0iCfKtlo3xxoC7dB8qXUtVkspRiLN6VnyyqazKDKQfckyM8Xx1emJEjog1SpG/eKzF
27BizhUJK09qESzSm87phvizQusiWHLyBPTpHDZmOyY8ksVPIpkHa08BeN7JbTPOZD6iaKMyGuZp
PijASI+1rR8LcMchmSxheXRQEddJ4dAvh72C7jQHf5wU0MXzUTgOPYpJug8NXXXtNx1gsVFUPPXO
jnfJCCmfcmYcU5MkCwLmC1sNKzpL1QbF65u/uDX+Bw5Vc9DPoyCpQjS5XPngsWAjkIrbZ9Jp7fPP
XGekjMxSqfE6dtHg9+7B5labR+b1M9vnWRaRPaTxS2H26gOCqhDoG/Wi23UgkWnIB84TxqRSgGwd
tWz+daM9utrRsZIKBH2BU+65zEQlbMVUbBoMqqCgJh8Z9gWN6Fi8EwPntcUuSMZkQWaJelgZlJYe
aT7xLcgIrunr0WZvx585fpapIULTFUnk0rgnTe9MRnHTgYmzBA3hsGX9SmbLiql4z2wz5kT0VRkB
j6edWP2krAu0sWdxdt0qPc1TMZFeVoGOCD+eRB/3RRmRjfuaP26lMIb5YTlJX+cEW0JDzw/t3P1F
fpIL3bmrqpyjAsY5OUayTvtaiQkRb8VSiwAVQTC8IdYNClrM2Y3UHjBTBXLjq2JrWw1dxi82U2fa
UqHM3Ewslaq3PvH6RoeCJCLFIzMJlNT4m8zGUfDRnsFpwrnf2q6HgKYxLROT1x7kqvI8i6EykeZ5
P2eHwHEZD5sqNejqUQwAVQCnYeIIu9lPDE2gxjvghF9xth2WO5Dm1yxyC2zASo6R6X+gtfXM1cO7
0xj5zrJCYxX6NZ6rwtBf81gIQgFbniZoX8OOIREaQHngR6lhqtWt5Ugrd9EfcvfwPCDaHOIiHqs/
mfIwKTm489T2eBxq5+MLpluQse9q218DaTzhrpSssI7BDE1jMkVtTICUtlI+Cp02fnfVdyWWdKKi
/gGXcgqZGzxl+mYDZbc+BlyPPABnm1+FYLTnokY3QbYlglv73Mq1xWAC83sAJJ0bHOKL5CPW5/xZ
VSdZ6AW3fSATB7UJ6FmEsxSAwaXNw2q2zS+Be7BlmvFy0qcehrUL4HM8EP5mYta0eHpbLmEMYfWQ
fujvcmbl7bQWpWXgEo6tR19/uXERypb2D7atF5TZFIwVY2YhO0qD2p7jVqHanAKyiE1Uiy5pHxvE
kOebpI0Om47LTPkDDXOlQw9WFuO6G+g/Nh7uYy7LTdsdzPExaiVtWKlIUaCysGyhCOC88hz2+vtH
7BWdUlrgT7pXfB2iE1gjDVq/bqHn5vAJjkC+rOdVfabrRrfppedOmd9ocWGtrsypAnhu32gxnR6b
x5kz/+mYrf2bd5xj6+pOiK6qmUoIfEAiRi9kXtc8Q5v1EaWv2nznmDlRmKEbcsCfQ0SkTs1kLBZR
hZDiYsO8vSyKIBWslc6lhgFQ7ntAt42gRmwc1AF3hrTxzQyD1+YmhJ3LvQ2JpuE+whoia1JdDaba
ZR08z4zsDS2S95WVgW10+OnliLuvmAvnAyOZh1NvZwbvGDDmuNwq2LwhQg+fQxcBuNOG9s/zeBhf
ZFnHMQbWR3yXJbfLnhMYbx+EmvJI18Eb0C5RqO03XTN/NVkVlmnwl8HqQ6t543x1HSAB32h3vfoU
hgdbJyRbTK7NTwHwdQTiEX7ej7vSYkh37ixbNqhQmW3nd6ZFF89C/RbiwmROYYpQa/nVc+43/bZg
Y97g5mWg7elnVlMSVVXuW1b9ry1U/H2qT9TwO4lDJZb0F8vbb46qYbRt6oeHKcP1NZ3vr1QnaFy/
Pd5qPspscoJI9Oz/lU9UdiwbOrIfv3y99EY6IfvHw29sTawxPIm2/2O3Fi1rAis11Qga2XcB5Mf8
8Lxf5JGBhvBgEOt7uA7hoWdKzKu7lGPude9Gz9QbOJA0DRK01jmy7WmDJwKCEmAkiin2cY9g6Deh
OheCOFKM/gy1yoUwuCo9ORjZKLtprXOErjZw02lP3dr1zGW+QLXY89Di9PoB1EQz8fRscutWMXJl
u3gIf1CyvIdseQ7n12TC7uBYD8HPAsa+jh1wE1VTVtDFQ/48OhJ6DHBQ6Kg+Z0RUE4XWYtmifUkn
2jpROijqkyzDyakNf/LT1S+d05nWRNst+R3UCJoy9wgexZMm13JLQt8dqFnbwS92a8f5UZLnEjsR
5MFXrWBkikrrJv46gkkU2UQ6elhSoviZgaS5pmEqJiq6BnBRj6zU7jR5V7MrU2NMNWjHDDmRyKE7
V0ULyuiK0giXPNQDH0+CUeeK6Yq8L9llxXSOPUkHrk57CvoEhQcDo5i6FdDGeo/W6tpfm3qP9jf0
FLaLIdUW43pi/wxl5ko13IHbg2kXnfrUG1Na1k5EkGKXA4DIFxnSX8LOfV+99bb5j81ihDOpl/Op
/CAaBPMknmzUkNi7NnSbPsqzct4j0y+M1HBPFNBlJ8/lfwIVApKF12XRD0HuJlqRJaM1bWQTA3W2
xBzHhZU30xoUjACbQxw+PZDiO4BLbfuV5Sk2iSoDRFYHmvx/GCF16OtNFXSzxvp6q3oNcNzeyK3U
a1OKA5QA9gqWZ7PlnLypaiKKIp8cl9qr9/PGBwLxXpCCJo6eXNBdiiI/XiYLqc1IkhGZZKIwPa+6
ac3aYH5I4AlrXK+eatf7ZgvDRSHsfPktdcEtTbI7CSgI5XWEOPxo1CSaDfdN1EGgh419tAJTTTsL
MuIphExbm5FMpN3gGwHMTYKa4FZRzb4EDfbOJi6/MLzUUXS4+8r6Sfpmx3AWrMSnhdtDGY0bGw+k
/uktQwLRTLvSH92vyQF5eJDfhtlqjj0q0CGTbJav5/3QqQ6Yu/8qY56/2sF+EtrPoaOv9/+KlSsk
apKMoGS2DJpukUjTM/WuZ86ZPLRI02UFXqe0Tek4NYA2WQtHmjYNko1xH+2Zmxt0qbbUvORSZJA2
AR0B0rgoR53Km3VtwBYOxfit+iGzXucDauMUC+w6wupjTBok7IZfgQCtKzvua3RQEGCRwC5i9ZSI
XCJqiNhgEKOR00mucHlMkEMULJ2H0rnmObMkkaEEiBS3monq7JbXxe98WJtyyhRTvUcV8JpaI+Hx
q/gNGGrANCVnaBAz49l7Z4Y5m1FIHuNRkdtVNVqpghL5l0FiMhxAztOk6JTD+Ry5CY3TsZ63MF6E
nnhnNDAIgmJNoChk78gVM2xpoKuwQd9H8rivlNZfo7/Ewkj6CpvFEPEJDY1KHwqgNIOvFOm9U0xI
+siRIbpBZrEzPYCsf8pYbwenLcq3vpIahaA9tFJnBoXGHfYBmTNfKOIR1luSlzdE1E+ZWBB2JAIY
m5HAYvyonrE9fftzg0dJopDcARWirzdM45my0lUeVLnHViIAhrqy2FJBoX16+TVmdrG6uPO7eW5B
lqqvhjoISGrjtrkw3Ka2dsgisFeIUsvM1YJfVVVFYPoDu5NijjbRuHBxZqWBHcb500WQ4tGy52CP
0kghvoKxWlZTqH+AP5wcOFmu/qPpjrcij3RbrUv32EOiOrPDgs3O28Xap54A4zI1nNimg6zP/797
q710rpBC7DK84Z2bLoWFDguHjaHonKSyZwp195Uex/UR6j86Zp4wVQKHaSV8kzq8YNDFWZE4eUlr
1DkMxsZiYceN30pB0eVI3O+1j5xyyJa1tPYLOVcsJVhbRckYmiSqePkS9NFJzEa7fzOUrv/I4sZ4
eD33tTrG3aixiMoUlsW6vDNdtF7KKMFCoJ/of1Eyp7/i6y00C9WZBahyR4IxuA26ihbOD+p+O9m/
OgylxLsvlFLzgKci/77HN+nOqNxEGlfLUFbpjS0Dqv4eMwdHGF0eYFb6Div9jqNGULbxSmAKqI0L
nCbtt00HJdgsAMHtLuIX/frWvkgDsIY+saphVus734O6rlHiGbem/34xajGWo+JZvlANbfNcea1k
KjgGT1ai7w1Lb/rs/D5ybBGw959J9ZS1y3PDl/EruxKmtXzXArdLTilvWA8XAAyMLxn1nc9Y3xvZ
YgBBm+0gwHBoIPwBSEMoVMAZecYKw/avXbvrM2V/fic28Eua5wlGwMbh8TJCMZSVPBw/XwzQlybT
YUmlJ6kEUF6s8sge4QYL3YxOGGcFSeEcWUFSJQseTQBhAS/J6bk80nSLHrN5WluOtKUxY/hWKiPh
vbY52LnnyQF2V1tS3zenWtSkaSCkyfvgvTsf60nqHBq+KxBxB0e8PxqZlKZ+NR9f3dOlbOosO1mS
Kbqinr3eBDcXr1/Pp0Hp3KpoZJcYPwkv54FLSAr+5epfnGOV7MDegSxTNC54loaqw9N0+Bd2zmOr
v8PdBcejxM6PIIkR5ZgwpS1nYdfckcZ5ha9JftD5HO5Mt2D3oZBtxKepmy3ncJZiSdagotd/vkdl
hNT7LHV5RSwTqIRrfbyZKy0CI7dM83lPFg5iQi/pPzecIFX0JaYBepONoaAm7CNqQH6dgbbQHtXf
ZMsnfIFb7ddEPs6ZPoCeoPEkzptsYusuWBZg8HQ/jQwomGzsvHztb4TPCrR/dVPrwDOnVn6npj85
tatZczQ2fW6BBw2Eyo1L5Uzr2Rr48WNwnk6yM7Wq3fgtKD0Cey/LC+Emz+O6B3aR31ZRIw3F8o1F
pmy1CKa9uMtf6zP2ZUgUiLQYBK2sIYa9kh3FXmib3IwRbTouGpuwhkaC+fIM6wppf3SfBb0FFk88
2g2g6UijsUAAwHo0kPIGxAf0ncApT12mSddZVLZJdbm3sCxUKMgj6ZpoZsNy1f0CE1ZmdgiMNWaW
YHS3zTitQgGqtdn/3pqxXjiT9Q9g9I42cMxvjsEqqKWMTvUhyQwnVc0HgillxWwcMJIahvlpm92L
h8zaLj4W3BDmliUmO4/M7H8RUTZs4GhBrMVpM73J82/xSXpERpusm4VupG7cn7wz/pLXe2k3cei7
Q8QLFitYDNIUL9MdtHgMRSCLwufqkTNbFgkRmumtFpH6kMZST0mK6Fs9n7XOfgpmPPr7CL1Yy9gg
Zrg8sOze9QirF11n837AZOfrjtF9NC+gmtpbMq5TVdjQaqCUB/mN88EVniuSdDxNRq7Xf0Iee9xR
v/bUeSRzFXLHh91Ia6KKkESEO4ZCsMHO7MX+K0vYFMjACXbJDHSO6w6SEs4OoFDz+mMhLLyMt7vJ
4Gk5KxSH0J1RvGu61LaMzWLoIuCEK+/gsPBFl8rC44gxxk4Ji0u51/WMJQpgT+NWAtSh5ntaNkSN
U5dT359RM0gFQ9cibYlW84kQMtYMYYQP9uhFG/skYvm5tM9d9noE7hnNodeGjTn3mvdwVeK5w0ZR
PM5k9W+dfvf8pKFZGT5T9gM+65vxzRtbEZJGbnl/C0ke/HqcSffSC5V6w3Zv30luGPw55kTj5ZRu
Eia2xGZraGvVgdEDCEf+BWN8Hwo0yHLCoCpG3Uiahugxgkop4i2MCXEMsO56xgu1+zEc7SPbLJWM
Yj6AaPrL6+Whqljq1UcBmATR8T3fsEjEpc78GVfWs3Gws9Y7k5kbW1t8ODOxLTrSH7BdqxrnIUOv
tIapiDp8rAZCZVPeagsH2bgPQJtX2WHKb/KJBI58z28t+gc8nu5xZ309S38r7zbRLWE7+U7Mdy68
7iPkkGXWk8mk4Rai2UgHMFCfDkMz4nP7uWsZSAt2t8hLWTp3Au5WQaOckV0MuSx6cMe0B8DFn0/U
qNo5LyEVZ6Zt1SqC1YwEVcnhvuZ8HwG5EAMzDDzlFbRiX8QophbUNG0yNGUtLVhOTELQ/RzuJhg8
BX82tG2+lmT5onBnnGJCefuPQzQutbVu5fb0d+ivxzwciGws/DD81415NciWRpiWEt0xxpKzr3BM
/mQp+z25cIlTIO7tJd1DZ32M0GqW1UD1iH5jGxfU6OIrKwDBNvr55IMpQsArR8Ff27Rak6ly+AqX
zpu9jJsCH8IHRXJ6jdvbkS53l4dAbhvbkJUyCbfWqX46SuRGHF1ZLKUHCJgWTm0WrWjpDUM2oRCh
3hFlZmglNR4ZlMVjVB2qB1nPh+tjLcoBZQYyEvfpQT+uRYRGu6nw5tKIutzrjm0Dr9Z1BXAbvMFY
CThAT/KJrAFhUoYscOSkTI9+R6liq3ZcXiBChIqCDly10je7LZ/1jzEqm8z2kC804ndKntgZF+Ml
d8D/YX+ke8e0cIV/wAZljusThDJbh0Ek1LVul7QcGZFWzmLRP4G/YzkeRYtJr1Oh6IDWZvAE7zMM
60VhDPtW0MOi/zHLjyZfZkuHDZv3+AaBeShNGEEsH7rkLuavcMpMMuxZHRi25UDWE0Sypl01sQv8
xZUp9x90uNr532ZDlx2r2B2nxuqX/OkuNJW0l1Bsg9DtJ+i4nVQkXM8WD0MsLRZdqKdECYYmVp3D
5O2FgXOIbnyp1XvHav8QalegTzCOZYjmV3/nOcekNg0iaU/PnTUM+MMfCBQ8zyxby8SxzLD34PAP
Z86f8vJec6vchi/0ppkBFuWY1YnatNERSD+2bodqqwtB7CVXAz9dquPkWB9arewC5Qf7LKziTIgu
EwnGdAx7dOJK8A2as1djNog4fPvhzx4OKXaxxY1E7x4Fvdfv0S5ahDsS28SOoelT89m8IrmNAivL
AEVkcKm+ybBxtVNAyGBk51pfjlIelMOWXT9ypW8DUlTE3IrvfGh9f/LcwdwCGaZNgmWFTFD7SKa4
WDIJwA+kdfct8i7PW0+N/x63dKzF/Rna51x+hKhvZ9+dhrcEssWjFvRI4Fo026+MyOvxfcFuYYl3
NTH/3GHOLLWDAwGo4f8L65zw+DQuVuBWbIV7EBm2L5Gqtoan4RjWaSIm5Gq5c+aC0XToGZaNRDY8
2xW64jzDbeoWsAIE78MEqSueeHKChzre9j6cWiE0zFLLeVXJNrNlxI7S2KGzwBkjk7OfU0xxxam+
oILH6fy/2errIgU25G1nTM6jKR9O0Q3g1JELyFNigD7C0xthI//Lq0DTWhKmMo3LrJ18r7z1XqPW
Drpt9hKWH1MbiIhjdqmXpg7dPJSWfrqCbXQNhAMG+TX7t3jhXSV/DcwR/Q20eRjMmfYyEprWpps3
WHjTUJX+kaK9J9/9JcrgKuFrXEiknC3kr7mp1Hs1b1a+wVuV4hbTyhl9fEnJtMu4Lif1oE340GSm
iXruHeURJuHxb8cSnP6PbYrCd/6mXS+ZxW61naZ6xNjdKJMvWmnx4355MqZ0xUdBy5/wvvZuy/F8
2X5huF6mlOJ2Ko06VJCUK76jfoCaWK507okYqVFZtpUhWkj8KAEk+OmV/qgBNnc16Op32biE3Nfk
OU62tE00iCVU9G9ECnc8mdOzo6rJzMvOhSdgxc42II9U4no6gzx6NN8RXrLG3B5GqzHvWnWh+9fB
j0hwoqXieiXz9L98fLYP6hlWthrzBI77iH4YRGNyurKahAaE0L2jTyntBK87Fp/CR2JxeRebAhge
pVq95R0e4+yF5vvl9u7cMwsHR7y5nVQ08NzQJ0BFM0jMcDTfquKiRQPDaxN+LqAp+k6Gg1V34cjy
OTMApStbNQ/8MXR1bw+TPY30ZLQAflt/jJKDsKME5641k0xcsPC40gMcCf8nZ0eznJdt/hzr6PAX
TkG8oG1qU2qmSLBGskGQACHtJEkJcZnXdM/6R3jCkquiT6KHCoseBz/JRqF6Z2z1PCpSk/Blzh1c
+PqMJO/03tPT989A4yaaJ0V1B7rkUmNetg2Bdz6ltDyBMod4YHG4xJ+dlcE7CrrK9dK0I4U0idw6
7+L9k+xieujn3VznbBSATe2Kh9uf4s2VRK6mrZM4TGXTjQcTJ42MFhtWVBFzg/d+lRtFC0W7OX8L
1y5yIs90V70xZk6IPz9i54m/eHr1k2MfIiJWvz3MMacVi7cvjF/lXaV4palLX2+KGI1nUSCl4DJ4
iniRfLJ1A3kTlzx593lv3qyA75fpV96w0bLug147vNtsZoQDalvHlU7N4b2JaTuvC/l6WM3kuni1
qRhAYowtNpmLmaeUPTGESnhvPi5yhcc4Ac/eau25nQe7ic1xK12djtPTAb/WRo37cMdyDFiPXhli
fTinKItnOh06uFxG0c6pLo7RXyFnCFQEl54jgoJnU+s/iWjX+icy9wHbnQ7la3+WCJs6sIvl0sv7
XaVqE19uTFYx+bNmhD2bF5cu/fnioutzqhadu8giIF5xMoKwp3qdFAnQs5DQylXYzyldHa09xF1r
eC3W9mimUhvQVD8LJzSi8eDxeS5poxXN0OcLumnxrOS4fJuxdDzFyIKTVlLUIC2lVwXRNevOc1pu
JEXaud2CkY1kYvsclwKak2T5Eik4ROGdQcrbbCEKW/d0lz2HnkWrfg22iGORNnaBHX18E6D2XX+G
wcw6xyli9XJybW5AGbjlz2yoGTI2jlYQV0MlhewzyYHwAEUNgzNlBiWaskrHb101egozcfhAZgHW
gvmhnq0ECU3QCdehB5FcnmSWOTT22g8cjPRLFMHMTmssN+uZ+/KVApOrtTA5ODw+otZ1diqbOafY
La+eaqbc9OBgRYdMdwmKnoeC/d/F3e67egAUZ162eC5t5jK2X8VidOsyQLDRnayBwVgG3BR037mB
GawhngQwiQ1aUB4KKscNvuGyZ7hGLAkDENA96hNX1zgMdHT85RkEywDfvv+w0WTYKhDb+n0IJGwy
r22PnF+2yc9yXoT35wZKLmLKIFfsq2FvRSJH/Z7eznwlpb622LzukaO4XjaOMq7ykvXmEWaPfEiW
TRrok2Nr8HPghhpStOQnksPkRqpIkxOAN/LjSSAxeUyeTKM3mgx3cVP2SgoiNRB65wv+gRSMTV/s
vfz2KHvjnlkFiG6ODsftrQ7JOe7u02xQ9OY4PhiYmP3LKqLfLfCqb0fyEypdtt2ESdLxm5gZxMc5
tlJIazolVzWi2BGgdb34ALnimwlOh7Y6lZPkC6hnVtIbLEZsY0GyMUOvJ4BWCEbBcYABqJElxJEQ
SBekj50o6jCA+38aP4D1wZQ8boQiTc5z5GqC6/ZrFWDs0g/JIp1/gbmmRX7DmXtN9wntVlagrTuQ
yrC0ZYeS23zJa0dr46QLs0CApgWzruuzlJ961B5tmNXj9W3utyqOqVkikz3pFuwI7LFICWrLbqTx
GgBjsnnW+Cm44CqXMjuxaaDVOCchjdHiGpfcklC+FhzOSBo5iY66gFWbA3C5Qcp+aHT8FRrlaRJU
cf3dZ9aQ5g9PbFo4y7G2YnLwbDpB9BT6AlvwsVXWStB2DmireB3nWhP9oi7cKu+wCNNJ5iKW8QKd
2NUachtpmGGuA5j9I6Iyi1pz7pnz7FHwPWxYGPJMDQOCV3suwM2pOLRtlmpdwr7lBmhUghY4EYzz
yK8WTmo3qzIS4mdwAXZuLui6/Xa8rITsB3ylQ8gzF2ezxrDGHJSn2IYbzpXcSBAImtbEUo0iUHMG
HNqmszPD7/lH+4Uy7mfq7Ka2UpIG7h9mg3+1/N2z2VE+uba/+miMeC45ORr5Bkoe3St/0c2cdqQo
uEPMmKMybX0uZNwKrKJZRSrucFyVllJEL0iIijEly20I/9vLfg1p5SnE8PSC5CrMZN1xby2z1Jrt
Oh5qQYn+VSY7zazU4JzETRn4zE+QQN+34m+Xglfvq+scn5lWC5J+LqZNVLvjeVOBlXlbdOyXhsEb
xbkAdNWN49bEmmTReJ089J1K0Bio3Ue59MfwwUbXaSeALpQ8uvQ7KcT0cbKltp1C1cgJTTii/kXv
s1+8vnh7zpG/cKw/pBAUWVKLjbg81U5JmIW1ppenStHgLM5GaHxtkC4M0s0M6x/baSsVLOfon1sb
CWvbNxe0PLFAUEqqrD0kGmXsoi3ZOz3lxDrR7tFyKV0DiLv0dZT1jxLJVvoasqfKkZ+C6Mwmj8f5
+h4BBrCti/T4ZyS8vyxAUwU9HKEIuRCV0DzHNo88Mg6PIqfprBAGPfR/vVmU9cGByzFcsGEklrpM
GBKjCbs02CYuhXpPXDL7+dq9pWGI4JW2F7CummBJwk2o5N5dioHaNZQwDSYPdQqDBAApBPLGi7fB
thunNKuaOuWjjXcMHRR2hQaUAD89Gg8FVpXIHUAoPvidBZzvuFB8kDdYDdzoVJ2Ba+SwIgzOGr1D
pDrqQ7L3IbZf6Cuyhg/VN6Y/1fnrKbveJ9YakZY2DssvsYFLkLxC2vLPvcsF8TcfGFFP38kOgWtH
uz5MBxlLJm5bPyybjyVE8JSCVAzwv1n9kV1wb8fghjqxJWij1+4v2vV0bxUDg/W5wgrpTmDzGGR6
BzZGfF/0BlU5WqtUsmRq8jcI8We9Km88LLZqdh7WiUyKDGmh6A/S6zBbpuE9AfSeXs21+7HgZwxa
Ij+pBJ9fHhF3Dud6bVLyY89KsDgQlRBTDbcTtVce+v3vG7tdGintPw2b94Mm5jb/MMuKo7B9f8Qq
CqspHpHStdkhyuxOmWuqvXzsmMFUrCSyuE9CiBkriWG2FYo4hTE3VLOP7R0JsUdyPyq77TffrDfk
amze6MbRJ0hrWqj/UPBX6z/7BmYp82+0V1DX1m4xJgUKRMtMhkLvpwKEugCoqZI0UUBu5AJJFP2C
mNVkAEyQqZZkpBILNyLZ1e44GUfpr/Xcn+XI+BZGYfbYs+Psul+uxvkA0BXOnSpdwcT7Pv2gkCnB
whwVm9UGptwEWA+vrETC0gDbtunJboMx/dFfM44Yasqqqn107kbWjRxVC4papDWI1le1px8HBlwo
JYYYFIPNyjEJkrVT62ho16/wkDCAh4tEDs0v3/Hqlgx6cQ+ul2vifT4rQqpx7Bx4F7sowVlqlge2
pXHnbP9ndVjbti0xOWTvReMe4vi8kJwXMN5ab0EAkPUjN8kHvTxJhKTZWFRfuOetZ71DIdXQVg/6
bxVeueGw7M0ZhBZZgEUY1dHJWFgbyn/bvTgb5IGc9G5V8x3FSbb79GM0Ca5DEDr8U92+Oomj+d4P
jONvV2yFnZThncbsmne68Qhc2ljlkWGQpuvHIbr8fBr/2JChNIaRGDon2ar/Hz9sbUqmCdSwI3V6
L0eWXeCZcbcYoAsVCd47PY9t7GHNgH36bLnRbUtreeCaMa3ZPaHsaXUe4hl2vh+Rl+KcwlKP2UAL
ud5nVgtkNhof/wTziTroYo8yzd2y233VOvWYd6X3G4z/I+rXR84gR4xCfwqPN16gu091TW+jdXNY
4DH1OFBsKyUyEGsT+e+uPpu3Ovdn+6TE/qNl0KefrfkDkXRK4oOCIkUVlbnPBjhy1DABWfdrsrFB
c6HzCrrtERrSHnseM1ztBqcsaq/kzlUsOAaQ/9oqFT8Tv9EIFBtbaKwfoRYrc7SN5ZuuzLDpRRnx
Q3NFWSG8MHTjZHWMTgYBCdVY49kD8/mGm0y6D2C92zj0zMGVzq1s/iX2iSfheDfcYlKTJPeOsMbP
u4ZF3yFAjpxYSCs7h95EK1XtVutDMaXv4rT/REePnm9LKshOVtXWpPBCdu24bJATJhltRbY2GRTs
layPd57wT4dfx81oO2mnB0W0IJgDIeYJHDZQIVMSIMRfC6UKKnsm9CF8YSAwNJt6NeNLzBiysgLw
lGj73GvbaHqDN8uhR/CmfjyP5St1gQOIp+oiGPg63SF68ktQtU6sVklrp1FBU/42R2eh0ozv5HNm
53kXn/US0oyjnHIjlFeWj7ogAmEsy5kAzjQ9QtmO9iRgfoxG6t9PUN+qdlPzpKdSeD8+j9PErjTJ
WyCK15q6mH4FxCeEXjUXzeyb29s/F1szSH4zN3gvWccyO7gR1u24kn8drYqpNR2kqw7EW3iD3h59
mk29bOnfFfK5BsI7uBh7oYCufPdbMJKmBjoeMnQqPKP1ESGr+tfc8SJZvu8HbZ1mZjT3t1lIWGmR
KiSkD2OcsvfHKoOo5h8V7o7+S0ABjJySirH71lScmoSYQewnA3PpmxYkFwpmuwQ5pK4dqpfW6H+C
DZLCKqOfsWSUj3Jg+3Xu17U7gusyEZ+RM49azoenX39vLQiThkhB+BKbLN8LEsqzX8rWcsNalGXy
rLudVKzoV4puqBWAuRgYnmBpS5I8Ol25nrPPy2iEnDep2xdbqCSh+f+ulT45jQxJhzAK/iwwYTS5
JvT+pCTcQq1oia1XrOwArJXGYhKtRQoQA0vJWljwinyipkI9pIhYFDgQuGtxHUOFqbcry8B6YXXQ
b7Z35T4vxeETs0jATYXSw1Mu8foAmd/+dCDS1P1+kGAv4VvY/i7iQy1/M8GzfwbB/zx5GOIOYcB6
jWNU5Og4c+xmSMLi2nphEY8OWnN7pEJ2SQ8ZQeVyL+akrn89SVG0CvIwJUs+FVvS4Pl7Np80a1Pt
knc042aef7rXlNAGGAzqxo2sOI9YYWQeAD08eUZyfCjy8hpu94QoDPBjSxeJK4M1ePcJxLRxWsyg
pLVjkIo8Ro2euLlPBUsZy/sIVHshdWtiPLbJvr6PiQYExw9e4PaMgMauo8z1fOxJWjpkimYHNfnC
QPSHEih8XLtvKxvS+e+hhXF1/mf8kWWV3URXOJa3ZStRMqlxtzcY2yXL/Csa5ODi4a10efiNf48j
/8RRiLpkTS1GwIcd2lcqLGeLGTW9APMHU9pRsmkK4UrG7B7kHFMoM6tH8FwfH8yjEXimLpzM1529
+Pp2fey5BZ/zllqzD+UaRHFVXrm5qlUnoTouAkReu76oEMmDvbexNj6jrh95DFjzz75t9bAd6PP3
3EH69cnad5NszySj6HWVg0ORZzVU9ABCmepd50y06gSuPs4EirapqU5jg1QwGKlBqrq6GuFFieb6
1/7rlaePco7PCYUAeJWzjiCXn35mOH/nriKmRoppq3BXLSSSeFOyT6j7A77bJYcPsFnxrTs1LqFz
qPtJHl4vSPyq3D+HngmiLBs4Xad+n27U/KzLfRJLLhLdkZOqlG1y0sHoHnoOWhEVFxLXRZU+MlG+
DC3UwVUZEIGEthlDyXHCLfDxTm1F8gaL6OoHHXV6TxrHD8qRrqqz2DWOQ+zpeuq7LwZltsesdPEw
mLTfHmZyDoR+V/bm+1GQBsTDwAsoHHHqOVYxrAp5d/xua8Ro+aJ1LE1pcxm9kD8s5HnzvQKocK8h
Z0Jn1g33vjWW90N+pnMKrBMspu1S8Jf3jWKKeL10/+4SNUj/YcnwDJtJm1CgGhf30evLlfEA7BDL
5I1djWPVeY/Q7IXvDzrCajVGlZ9nq1eMckFK6IWBCQCkGl5p/dPgneFBGS9p99ktzfHSPisAHmP8
LLotvevbYpZsAFcmu9intuWNhAGIgWcn0NAO4LjjmouGlVi1TCKmB8CrsWPlguP7DAqGfxidIoGD
QvxphA+mKXtJriJziWV+vtv/40/jk/owAPzUcwGeRzps6KEpzTPxadnTv7HeM4yfk+zbpqD79eDc
+PFvnQ+LASyoskK32KFdOXAzfnFKHQ3EgCTBDITGNDSGLayiOR5D5j/mOokR4aRyShW2jwnfJOKw
O6vB1GoYMq5YqdLZEZU8+OBoiFWIjkIsjKtL6JuA4L+bukRKfUTHEaC1u5O4uJ5Ffw/mE/Pg70mR
54O0Ziw5LIpnLS5hcsyueTrbeBl3/QX+o9AcUdDOt2pURLp67AeaxiZ/MkPPWDgQRNHW/iVPqUPy
m3xijHaT7NVi9Lz/MLqUzf+Ie2jubxcuo/46BTHpgX3ipwt/xfV2S0fUqomFmRiWqA+LaakF72Ja
Ykou+F1gf5Vfg5rJfyGMqKT14PGODpbWyEVYss+AJ9OviV098wpfTKal8r17mUMXNVsgqHsGEaOl
O9OAX5d7xq//mnj3kOF47PRdo/X1xyWhf28JpsmlrpOsq0gQrherbfRW7OGh4YcirIqsCvisWj+/
wrLGVHyRycyDjEb4jbqE0NYPacExy9xjgMiSEMPn7LLWfHFSfmAs4pA7aq6lKDBxXn9o8irFyWBn
x2qrt5eVtqQ7wg3CS8Pn/nw4Hfz3geY1Bk5ZaSv40BgXvWGrrTFkKYthyfk3+MFK7LwIck514Zoo
zV/LKYAnxOAaMqwyjZwbgmcsPpOfodmdoN3060Oh+xmiaNuQK30lsLKG/1Ea8/nPySJ46nDFNNBH
btzCx4mc+pVYbJJ05soLAHPpUHi7hMjHlsoJvHh6JtBMiFKt6urZ5m6xWCbydKDfYtxmjAlEYBtH
MZWPWmPOtPTrVUqvZSEEm7iZji2LAPu+HekZMkACHl9ZgHDabBhL+6ccBLT6m0tD/XWBlU7IPY+8
WqrihzIAF8HgICeY/ibHT7PDBdjrDUyauxZubyo7iGBwPsoDSINGA3v8gc2IcuKomkFDOOnEw+o/
AE7rg6L4hGfKlBjI1QA8ePERVJZAb+juXV+NF9l6pqcU9omh+g+0icBwp821/x0wSAnbY52vz+xs
TVkWIisRH6EF1NNNMu6WVbQHsqJBC6Wc4yTXXG0h/gAdJEqYVMZqALNJnnddsIFzPJ/aF4r17SmV
tZHEn/ap2GrDXKdeMX3hfo97DNEGEtQAkMHswmp79cSsDhYBoJyO7ljaga6RXrrS6TJyAkaLcAfE
kjUbat4MepCt1C2zyn/d+RubsobxDIHUXHziCVp4Vv1qUjcTSwWcRushlGGiIJPVNBZNAxufWwcV
8Ol0f/ETIYje74R94BiU/QXQNtfmsXv8WJKTdg5SX8d0HbNGKp+9r39IZIM5KyXbnJ1wzFFGWygc
qBeFU9im/uIxzkQJxGHmLuoIfZ2jVicjeZ2XlFREr51qEWq/0+kBXNmM7GvvOXaYqKyhi5Ie6PmB
jZW1ZPTRTq/qh6CUgTnAdflRCrk0YChtOLHJzlM8eLrU3rdIJ4eTwtQ7tj0T4b/+e5nI1k5/n2X5
vvz8XHL8Fxya640xmjlTlpgZpXvZAF5Esx+49Bo8qNrfmrzYeBPIzvSwfDI8bWI8tBSI62vlqGVG
5a3oDWGsMyjrUUiYgtzzsXP2rxTMS/ioT42KTuwOo8gzMqE+N4rlQ4ZHv7w/4hLirsyxLI+JN6fh
BCklLgeb/9cAi2ZJKApQbFtdIMfiGQdSzFpK/lIWqufwnKG/x0b7T3ZQNCHH2MsO3y5Wk7kRqrMc
QdryVXAKnRqtK8xd4P/u+JVGrX+5NKzdQ5d+cxgkdGaf7AEgE1IuGoYUFtqN56EheaJ2kAGAFrSY
/gYmL0j1DBSaNbDThD60rhuRJm6QQOlnmftFE9wML1fVXkCvKPlSa7vLHlP7Fue9FOyHlLL4OlJU
c67Czf0ntY9ys1+nVYKkNKiZkup7Tg5tXyypSpN76sgm1aioSO4GSd02dhbe5ib9uiI1xPYAIdT4
h9ubJLAf5qe0jn7b1DLqn35lLEhNpwpP6WyQO/jE+1uJEsVh+SraoPIRIzv0iOztm+rc7cLTfayw
T2z8k2EsRM1oRmvc/8WgfMwMOI8iRzy/lL9VjsdAizodpPqfASaSkGKJBgj+u/coHyhTdNgMrAeH
T919/kqwFTdxII5tiddl3NavPAeZGZXIa0Sb59IIpoz2JMmZ4b95GO2qocbe5I8ECtOI6PotrqY4
Wit8T4qgnKJgH9KCuXoCgniIixS5W7If2zGHp6cjysPblZ68VnftpubkwM4FymYgyqR2yRtUt0w5
mbwTmnQXuZ6l++5HjENlox0glHnzp+NJljBpBk0jSRpld1vPiSte+W2qzgXZj6iodthTjpk0eG1B
khzUpQ2mXSrZtfOX3dbPM/oiLLI3HmYy/dotnCof5FDKuAhkMbv6K4+IE9N98QEVvmy92ego3GRz
28rLkdh2/7z1n1rDswT15PTuGKBhxuBlZ2Dfm4Wcd6f2MISuuFejyQDcQB7Ej4FXoMLDf1YmJA5c
u4HsneqT3ErNWbbwRZesSz/9DwM/tz6VmrcT1G4SHk0k9SNtlr6krqz8Epi7PmcaVivGg7CZ04t0
bMKFyTsVGR9xOsvTahGCsvZHESF5fMF48xkJQMN6TvGgz9fOhFVHCJzm7FUxdPtjlY+XYwZb3Hx8
IztkuQonB20Fk1n4j7GSRW1s4MaS2Cy4b3dxbicAOeN3SSLODD7i0K4VZC5vkO1SxNVOyB+ZwGmx
EqUh9bjvLuAE1UgCSQM7fnd7Kwrjp28RPjVYwgWSnSbxSNhh0pC+tn/vswwuSzxqr1N7L78T1viM
Sf8RkI9uKIH/fd8BGOjBMMRU0Od1tMdLtk/+unS7+D0DMWl9oMOqPDbha2D07dmUVurNH2KkoGLc
3CtmM0O4/4KMvCkLgsSF5fF5p/fsajaag9tfBjKCbScVbpXktjC7nPleG13dtw3OyEveQvVzM+ZI
KMPH+OVOSEMF3mWzNgJyB/U47IAMgZOZzZP14Z7viRFHGA6BpVDcXdEL8mZ2ZxyH9nJQw82UHEzE
LIgIYq291ufgf1mRsVc/G76SYem7/SVHARueaQbRmHxQhcG4r/buARmF32JDLbB/RBNg8JQISDSn
OaDF4ccCr9YNB4BYfeYVW+pgaKh4hyP8+U/+tBhAIHLsb3Hxc7NHV8NeyDotMlkud7g1WZohPKPP
bsRW1Rx8u4kjSWCkK8luRmRM35iIKjhhGZnqoGTxHl9dJ/0T/0OOu0tSAqYWRjQtd8zJ3bsvcQzI
Wlv3/3O9zRVXR0WDxE1PgUFKXfvNhF+pU8AahUE3Kk6iFL3VStqAgyFESBnj+j15t2tIaMcE1GGY
cnDKAc6ogqzFlnwJod9NtXbhYtc1arMgeR7ev7FQ8nsoLEZSvH5AaLIyya9L86gvbgEyYT9goy0w
AldKb8O98W5fnzM0lDvHD9KXwIm6JdmCbjOgvQ9S/kGoHHyArrZirFYOhReqqEjEImx7Z4sRMJNi
kxovZBk+rb1U6EvTGMjr8G6M3QV55A/Z5Xe1pSxBnbw7VjHV349yzr64kfmicCfXt/sGLUgjj6ad
SED2ZUZkQExLmNzrNDAzFoWNGDX3Xjgv7X9mEVN168N3aPhoTqT6DAyyUL7O919Q67W7drEPolVg
uVFyq8tajK+k3Pm12XxgRJs4Dm84f5oXgY4lLHU7zvxvmEi2bXIVF6GoGuxC7uGQ2ho/nHc8x4Ne
0fhvIznr3k/4toKWuUq/asM4LZj012UFUGcXr7pr/6VSC6iZCzZwJHnX8Rvk6a29gmXbdYG/qyT/
XwK2Q0F39u6E6WP0fEnspjLfvZ2jGO7ziLiUcV/QO4cIeHbJgWa8lYGw28RTCVtKtFCeh+GnHZ7m
++npIZQf0KOrpEweFmhLTAkRczUfAx5B7FUG6uYLGE3+oEjFFkl+MV11Uvzno/ukMNW/E2uFSoXW
dIoZuhdjSmrdvli7v0p65R6cy0A4y8UA4skqYHmUg2LiWCLDhA24qjLHlllycSSfKhZNFLRcVwEo
nufT+Ex5S5NqHRqYSd55Bgyo5/lFLAq+aPw3thIqrtfUULY2PlcdDv7nXCz6hoLIp9LqKBfTJfnr
ibI/3b45YoKcVOHz8QY8nvv7A5/LOX07viIvNuDzxnH7+UdFR/DV78x8nTE3vzDp1g/CJ4+2ZX77
b//H9b6M0ar4i9EvFlBRQTkJ5sH8LHDMescM1A3HfwPzv01gxRruOZsqNiL+QLFkv5QsIYXqQENX
Ml2WL+aD+gCRTzt6EgPaDglg8UBLOQ3X0IqXFCGDqQZCobut8Zxjbi9RVv0negeeGz1EQB6eKxCO
5wbYdWXQag/kYuketJbBr3B9sf/9ju9ll815JSRJfOLDeb/cxGkl+pjjEIqHcp+0VCbTd/Gzm13J
c8zrSO6c0+NUv257QuRUG1wo1aQULa3CT69zEJTmAmbKXTuClMIO2xftr7olu/v8ffWW08LvO9Ss
wqrq3NPWnp8lb43eG/VC1PC3MaEiGnM5MAVvZPH6xqgx+/w7+Pv80uRxZu6CCRqll1VtkNN4MaIK
afjTxLRzmYnTiXJg3Oul2fyaRI+XC3WhOtcsQj3AHXkS+vPYg15ux1IgQ+ttJ4Mu4u6ew2nk0QFf
C+tccLyumbgzs8nmYX75XBAo29notaAupbxJTGwV4LMzQ/1Tad/Y7ArSCGghbTVMBflECCEL4CC0
AVU/kV3wkM/C0eAlIy5g7ySix8jc3PjT4bVAHtBuK31GzIfLJRrVwJ6vYOkM6fr3lR1OYm36IC12
qg8HPKRQXQUmVOUbRSlDN/7eW8GOgLXkVFj+bHidY7RBr/2ecXCil28hYG6NCuligxiFsFMcl5Td
zUdOsbDULhFz1V3/dsMZbKjlkDP6wZPpjNo6ozGjm4FH2op5txp/GDA7eJAdRkmCQsR1LROrtSvm
XCPip4fvU8Tq3w5VMYSGXf5XadQvPklNAB/RObvUX2wssLnVvJlC5FSV0YcLbJEPJyMZQoxdiJ6J
Vnwy4fumSeJom//JD/l7qAdvALs87d079ZsGXsjI+989wF7M9gHDsMfSxW+37/YZYd7In9F0wWye
mOZ7csQUxTwEtQnWik6DbZlQ4O2VmOzQJZrNqvvAEfj/dx6UQB96g/EWSYB9Yw/i8503Kd+2SNjv
Ov/l9LGNiV/2WCP+sdnnzdkqqnSqAV6mdAwVctYdw1K3MdNowM8vcJBWs6CvVMeGfVgu4KE1Hr9z
QxvzH9AaO8zKK8tYv6PRd8qXQAUnf5KnhIUno7wobaLfCa9w+1oODpvXmV5uKyO6onPsI1sSLdLS
+z3vVwlxo5Q3QXTfl1LMlVMCsiM2TXE+DzTh7GSYcVPOJ1cLiWjZvjpuT5fWDv42KuDv7hYWOpBW
K6m+ru8Iph6fBwG1wC2+rDvrEQ8N96zGDRQtjh6tmoY8v9BUPwwqcoDHVkmbxB2RCpxjJ1igOIGj
dkEOPgD3iT8TlocGzSQpMJKNQekJCXo624uqW3a6fhjfTPRtg+EdHx2T90hqa509dmZcz4T67u1B
PJbDGgjuQ3NCokEQZP0Q6ZSEIpLKhYslB8AWtp3zWCuNOAV5d8qyOcBKoKmK52OxQeG6IGvtAn5D
qvMnQsRSCRzDdjCBZq4A0yTnb+1AUFo//UeQfTJ2c9TCda6P5CFntTmSSUYbn4aYvWkbeEEZSTox
iFhXxOChjp8uXeQuqsmsh3HpkG+mnqqCW0J0zOqOdgNF9EHw/JX22DrVQbGLNV91shTzm0fbE5Fg
AVurBZq4EWqZ3aee09oKJbmqdz2KS5vDbMAwugvNsDnXR+nmgv1dDShFiUA7r7huiV919W9JnyTe
S2nA9v3OoP+SGUgU3xXjsYwfEOGwT/gdD9nbIvbrrt3J/B66CX0gdEhosP8gQHrrkcbTRO/JZ9C6
E/aAVouI5N5F9o7YJkN5xcIolPh9b+vzJ2QVOdnbwQnGVb30ju803sm9hDdun9SvhPD1FmFBANhF
guJFE/NSyV88aV/KHj/L8OZBGP9jvWPSgoyCoEvPxfh5UULy6uJCbXe0L+r6XSa/aEcchaEs3GhZ
oCQCClnE1xBUAYU5sYSPzeOFnHmgVJEiUQSE88qXLnetTEwENaWeopAKQgXsYq+7YDKX/+ULaMUF
tMHF+B666b7a/REyoLKeTdrUKMe7dPTSBw3rlnW4LJ6ozzmM0D2XK6nf9RohqrnpXhOZZF5pF/sc
0kkbPxZ8m9OqJrv0QkuDKHJxlhoBsOf1VUQRGiraIu6ypEXu/zIT2JjI2PKlAJz8/QdtRK1a4LqW
8GeND25lTXXoRAKexXfFL/vnGKQd+qGwCE9FoMRb8vi/9tFB4kIjnyR6JH+rzeTtLiSW5+7K1bHh
46PPt/L/4e/G/AgXsap5P7UIWzzgu9/PQtq7nr5WGElnpAbrkoqFTvRyb0XjYkf5m7ovSWRHZVtm
xyLezkZapbbcDZ0W4bw7DE6TF8o7/lmg2XmfYvaylc+ki+IadKJd6J/MAgXH8tH3evs0PySS86Sc
RauDQDWcb/EDpE8l9q4XX8oLhIa55USZWvB2tlYYGGBqB5/f5IA3xJO02h+D3ywOfGyBalTk7cKW
dAL05fYlKVFO9Yn5Kr8QVWEuTaJCZBXLEUWqyzFlPCacmMLtICDXRCovyTZ0Ud9KDtRkETIrSGVD
0GsRUCvLowibtdg9M2oW8rXv1yx7Zv2EhQXBLoRB94bl3TZDp1kdpuFNKOOh22HpW/SyTbXG87Qh
Tc30Zb4usWtRzukvwNlT6cpr1fIZP55BCuQEP1wQSI3yahx1aKSc89Yfu9BDcGq+FO8bgdsqk7fV
d3M1+Fy/pTc3itWBIRDTFf/E6V5hSCam7KCM5KE1fzkbSmR4XKmD7kyKXDyTV0FPSE96dq15SnKg
rgEq9zR2SoCKyQ44mI9sJHecC87Wko6bDlCExdShHdJ8jtQpycpGfkUmdzDQYRy5Vni0id5aZ7If
T3ow7p0yBLnHNdQxTW7r8enw5uJvBwhY+rcN0dvA45hoDPmowDIIkLcO9SW1bP2LFvFYeklD+hRI
wyRGuG7EDWVA9bexINiZDWtpmHFaEw/2ussd6TZxEB2t6V6xe52xVvsiyBmA5wQziO0ham12qkST
AK/v46SfAn8NwrKrWCr5LuVubnI9Ft3ncTT4IMx/YcS9jQk9DOGf57rs3qn2hEzK72T7nTCh2wTo
F87EFtlbNXLDc9I1Sd8j2F7tYaL08YYpVXNyGAS77uWxBhgQFTpedN+zaw7gCL5bZbYdZsrWG2gK
SPJcqnVQ06oOpfjDy0xf8qAhyrK0LBHWaq4X7f1RX3NxfZD2m95qny1iVYuzbY8Q8Nf04BEdBsou
pU1ZqTo4felxZJY0R7Igsf3Lbp1REZns8k9rhfbOynOsR7WZzqv5xZ4K3y66OZDm2Db2ThLLLOIK
QDnNvQbNFGk8P+lTAUNLi2RSdf7uaz85Oy2VfPrL5eM6LLvj2IeUgO5LmBVp0hcAP7imFojnSJEb
dEjgocwn7Yp8+5AjOgJxK/ZGp8105Cb3aSaMfDf91z1S5z4VAiENr3vprtAGLxgb6nvb+kjdW6UK
Fg0VTKhXaj/wrYKh2QMaojbxBaVOrPWzWQN2qoyXm6lzBr2bsydAPnS0XBVse6b5NhnbQtHVGE+F
TwWKaFwS7aH1KcU0c29EwjW/yGOM1hJ1oXLqyR9jGuP9zTggllbTAWlwAbS5CikJJNI/UKRzBG26
oAo3guP8xXXu8GRpWQgHAzJf99+BBmWUMjoMmTNw+FRtrGdo/LF7upNXEFJlZIBsbYIy6b0/iU1w
cqWI/MrqUH4rKFikVTbgXU71bOuEt5Yfw2Y9MCm15m6UAVCnqWdEcZ+tK9DmPL0lpvXPXAeZZgu3
8KwBRo4BVwmJybQzJOXh0jbnpJgB6+N7UupWaRbf6aeR9F8vp8ztnBzlIAxym2IqYvNm/anTTrWZ
VDOSDR3mUltHjh7p4qCzazAXOaXkd7yzFHU2McVn29Lq2/k+DoPixWPRO2z6uDDfCwjsyYzYo4Wh
pGbwF+VI0vIkae7GsSndXUb08Pjz9923JKXUfUkTE2NYpsS1tq1HCo1xUPcqsElL/C+ni8LTcH8r
bGv86jKXKwswZmtZe2yj+SQOb8wdjZdh6pzS3weZk9awHMIGF2H/uU4aJOOOIvLNDPGma+m/yEsM
Th6ZeovWnLNKX3TiLx1eUNb6sse2dO67N0UubpvLRCfh/gh9yFmjfNwuuB7395/PwyZuZ4twKRl7
z8goN61Al7SIoS+poEGkx4XSq98BWMvDCukSihqfbCfAA5DKuSoaw8GpARGtcKU+MRbZa8SbhNbg
VVNeT88+BbHGGsJBRBI/absqZXbRP0O4a9HsBsunCHCO8eWKkmPj5ZDuDQhUtfEx7kZjP10egoDr
4ER2VvKs018CSH+XY03UmyTbXhj6QXKHzxSWcxXWsU36XX/Jq9pH/yqWXnFDyTezvFu383ecfoUh
VLeqweYRNUtpkWMmvr7arC3AlQ0DccVTOmrHUQJ264IkcpAFkCFWHjtcCbYZL2zgmXC2a4DYxd2U
wkV8BZULTaafYE2S1OURia30VUUnw8BuJFKIpsPPjxTpxD6k0mMtraniv5h2ZkLS9x9qj79GEb58
j/h1yKqrO7CKNKhPaFrzZe6B1vBeuNQ+INTS/qkNHw2pJtRGG1zB6q5anLAn2DyHikVbVYmPk8Ey
jB5lJXSO+jRFlx+ZFcunRkKy/iejZevD03Z8d1grqmEl2z043ytPhhVs0T4UJpqalaSkyIgmvFG9
1HDo7hZSfVl6cD3Tqd3vCHVck4NSebEDycts6mb7/PerHdNkGKN/Jd4gam0y5PXWMPaxOU+oUL+t
2x23KEDQi0DNLcSOPhRyWe1G8oSB2JNevF4KXUYPDz6NpDJmYQ7YRVii4c684dnKuR1HKulBBsIu
gBBqPHiZXs7bOn2EQkITVt+LY5556n8o8G8BXmesLYch0fzi3sh9E4p+JIC+DvLNZu60IPUNxExa
taJZJ5StTF8+x8U8KinssXTBb+Ua4kxu79x8IsbpOMD7IKsqU84tsHhfJ3HmtcamvLzFdwDfJZAr
786WiG7h/KwvCPKvqaW8gx/NVhr3b8eNoEnAga6rY6mFzVSXmTEtAQmkkeP47vHt0BaOWqzQyUHJ
vg4P9yedXFRWKAy7amk1iW5U3OCkJ78gK9AtJkADP2sAh4Mw7Ms7nWpFsQ+gxsPDf7iAQ0A8EYm9
Um0qaxgxR3v3iWNaSyym6+PGzY3AJwdJDr7+GasqG6cg59te69kvHAfzzXjd23AdW8PjqFAisdUf
jl6zmDiSQje8aWQox9fCv+eEmjrqelkuyPD3fgujorJj35cL9Z2ltLGednv/F8iuzDh4AZIsf3Iw
USEFCufatmK42cWNdNr6/01EfwQP2MTxWPBJvwKEW2n0/MNOIMljOLXDuZjSxFHo3xdpp65jdAS/
vCpPL8vD/tmXY1wXuMjzN76O61XqA4iQoKdmWrJMfI2FGAoG9eDegg6fJ32lIw9k7uGZmmCEv/5S
rLxBBVoQSFgTQfcJlqsCZsfhUtIFOjOhD4rL/1uCXAVViaOCmb0/B3jgf1Tv1pBIWJ4bVjqcbKQS
LxHF5pAgRx9QPBnyb/gzzMp27XRi8OBqbtxb3LzPcNHdlf/SzxX9eJ/Qpn5i4raAFEOA8zck4dCd
pRwYk1AsqmXezv1+xOKYgw1xJNfkn7fcB0v5OihzVJ4wetltZFlksWD732BoIx57znjxukEmmqyj
ekyQiHJwsOxuUX7aOfCQTM7GOxHiHIz/TUxRu60PKywSXBGSxDMa1WaXxjhf8ahg8CwTUDMg74No
Tu64cQvxMOOryP8fWp2LNrCWONpDfbQlJ6oL5SbNyHWaN6q81qlURFaeh/FvuBJXUGXzz9uqWRG6
mLfaoQq+waemwLHeN7II53QFWmOQBtvuE9ePszFLWvn7RJ3VubiZUII/x00CspWtOiaavOUqkeFy
Vyvkw8U18bqjLGfYK2Sg41DC25K1r1Gy8vvtwWWcLWE6drnfhemsBLWIiIgYKEHpbCT/zhElpwJu
NYaWBN0J5ipCdPkf/1jXzLUwbD7imvuGSyDVfMk4ue23giAvndKBHelZneDQhgNQIxB6lhucMUJO
34GfhZ0N10q3agfh4zmXAyQFyeZJlFpdHWp/qcpLVYibKIyzlyV4w3byfrpSY90EPFFW4jMLyDnj
n6t5YhFVV4pyFxtWP8QmOZ76AG3EqAazGBE8LcdzqwcMh+cSIYYinL/zrWRFF3f7w53/D3RKa/MZ
1v9ExNGhWGEh8lv4vQ577dE9RpStWyR9n/0z8OQL4bhuKd7NpojjN5a5Dh0cnNOhJYPctoKEsO8v
op/C3NX2V6R5GQEh+zAOQ/1QZA7xIVMVe0a23Io7PScdR1uoxIr4ksxfdF4ShvpFLo6ZkuQ3jda7
p5UWZBK/IKD1zq4jW6jFGBy9yshkzBTdzJttLDgVkATeXOD3KcoeW46Iwki8sg4q6HIeiSZNepDU
fH1XU4mL6yU17+xmJE5crjT7ohcZeEahIxPGfPo1EEe6RIFuq4cfWcAB7o6z22euI1kxeTxIKsTp
tL9ReOdqe5LPdkcDoz9gx6gQ2nf5KXsu1hC1bqkxCn6QzmjWjrA218yQNaveFgrJROgZHIjF18fi
Z7Ku5S/PN7IvZdZUcAoVOH9lPq6JZdiK4PWbkP5QMNVwAXg2szHXkKyuqZxiV5RWdYm7xDXMNbV2
8kfEBVLZRKjikZgPImIIbXq6StXlcHEfWHdF5okrTL5kjh472Sd4MxEjms4UNa3lYbCGHwSrI3cF
gRm9hcPV4fqCns7ih1i883AHXU8hZhVjmQU3EdPsV3bgYqV+prb3hSNWJAMuMU0ubnMOdg8fxLFQ
u4oYpDpnW0CNp3qhitPzPw9cayTYa/jq16fIfm5qowKzhlikr1nO51XRZUAVOIGSt2sQwz0gXJIM
DGOKoLiUTgT587vMRrVaa/DMQ6MQcYY16f0rstIV8R+oycVZUUJcoT5IMJnjnDcwKj2bpL+I6N8y
bEyZz9VOPJZU5vUmOmXKy25lh3hdGcFmoPyhs3vAgpL+mJ1KUVPLe1gxBQF8XfcbHN1WKGCzeYC3
GgRgUbEpj5aBvHoMqIWY7Nsm1mXAhd5ZXMhknUYl3Ev2lEvHmLvldkW3iqIzs+XgufKfn1ZtoE7f
nU+7VnHrW3JtPMtOHKPHMpvofRLo4dXh99bi46Sxxdl82eiStzOBp46Wl6yuFgzLcYXOb1luzRA0
Wjw7vO/YGmDeoTNy4e+9ADrrSoSZMaf4M+apkaQ96yyp+NvgPoiyBL5ocW4SCLcqoGP++lbupTto
OMTMcVsYJPFmdwfm0CdA7fGyz56ENHMaCC58tRwWzs/95p51wV0bjb6O+1v8udIX6JvLiNOXOVq8
aci/JdgAcXaMrPGI1tLzApabXZ23uI8qOHeNSQXahJ7/7Qs4fKXa63fgp320AUiDOpKpdRweprPL
jhZBZWy5+55fGzShf7PGpZ1ZN1mOLAaUBMsWYmde2TjZ2Q3tpacdqZ2VkxIxPDN0RCfJE3+z6ZLu
91Yjixa7DOh8OgTp7IrGbS00GWxMGJt4DmqrpZa789JwC4qjRBdcwsi9gzgNPpgktzyEgXrLSBjh
mGwYipkgoiNpRKRGA2hMmUE73qFSFAP2CFbOAPwtM6e9MI6zoZMUyfXAMBioI1R9xCbx0khf/1eb
YeOOU6IVHE1PDIzjgmhQ58ZYUZvhj4+LP6JPzHB4jDKYKW7HbIsrc9K6HwT9HhDU3/3Zr9TALpwm
dzJzElYUB244R6QjFz14VhthmL3hI7HIFUSxF58c5AQNzlcp4tqJQuR7D7csO3p36ALQIWDK8N8a
C0KsPOxtTmwwyJziOHBtvqZSQBhPbnSHZREWfgmA6EvwH9fC58XBOuVxs0GFXgomkWBhhe/IEssi
RfGZJqsbGgJGv1k+vHNVRKH7lWYuyeFPHIS5ouAIcJ3WZPJmn7xBIokX9NN8AwZEsqor5TsaGyjZ
e4EM73AmiWYJKOORqfXb2o8rzmPF1DzF0R2g5bcBasD9MwvGdwnjfTUIX9Hf/9YGg1gn0golYMwX
YZ34XZ6STLliMX0Fj40HA6E5IwO5gX+CAxBjwweEZ9aihofWlCgLiP9i9aImP/XiOJx+Ij7Uwwb8
6V7kprh1nx4gazuGF6RpaSEsDbPpnnjKd0igsSMLSK3q8Ofyz83vFV9Svkxx2UNQHL+QhCDhDql6
qcUG58MS9S6xT9YIYBI+Rk9w8KrRrAY0E4OSmOOqQLedyGfRuGyPkMqQyFTc7RYpX/vrHjcxLp6i
UvLoktwcVyBMOPqw//sE4pjur4pMz7y/uC44nzqHgs+wDKdtOQdgdnvS2f8ILcXtIapdaVhqAHai
oWK7wUdOO7g8Ldb96fxUm63LKdLEHwm/aPrExYJLb9GdkxKlwZGZgAGRERxF8Wd3oOJ3iBX4p8/n
6NtR2S1Pq6CmPgilcXpPSMxPYjDDc2R0tUz+Pkoz289/h7vhnL/5faHIIpT0HKDtS3vHj4KscVJJ
cAPEusbfEqiSQFqlY3QyvGLfeccs8+zJyR3Pa1WBF6IqWptwCVcy+we/uqUri/zmPjn52kY6V+v9
YqfV8UTM3fcRrgFjDCfLay/aVFPg4pBAS0l+R9BglneHtC3CqSuP+vxJ5sViYfrvGPCC6B8GsG9P
5R92gKEBHtqDnT4pTm/vzYhgOJEfMOtYWo4j3qPZz9pFlMPSRNw8zd7N8UpZwWNfiEasBamojf5J
TT8X6GSuruYTov7VXiEnmbuom/poW5o+lpxEuENEGMzCZVnIxEpICZMbXK2hl99HHDwplHQrySiq
5L5Jgb20HgKAEmkqYxzgGxrDQ+3OIpV7FTmsTQUZ8l+CIAy/mCpoEtayfvQwcwmY+18BmB3jdj1W
hHPr8PadARdR8sBz4Z3Hb2/Vt+OQMX3gEquF57aAE2fcv/iV2Eq1Vx56SIA2YcvAOxgUGSVfpCVv
g4VA4/3dl9soRO+9ajzbuiE2aFVFW00FuYFfBfzmnSCd+Kl3BR3/Wes4NvCbBZ0M3lwupKT2rX45
k9o1VSFvCwVZcQ7T/TZmgURhpbVost+lAjfWNxC6aPFZsD1kEwDQvUP5IxbNI3KYPhqcaWR+1U7z
evB2dLjrMuxRACiSAHIhSW9fDK2yRnAHVhbkuF4i9e4rpCOVkPMUYA0FJOl8lm08AuyjElizPYwX
OTmA0j6Hn5FtatNKKSikeunuyMc3ioObX2bdoQMCs6MiAvQlEYmI8aBaZigIJpnbXADLIBe05eB0
iH1eX5JLU6HoSycJbK90kWFtDgMhBLoSmkbMTmdswRnHMmMwsN7RE3zdGSsbaCGSAFliY8VWePh6
ijQh3pCPTC4o0kjGGz8OR5qWSSrM4E8QZ31K+s2OQmVeSfkIoDJJTFg6M23j3cOn2Vdz1uu6/VgP
NeMCv1NBOEZPNWJatJN9hc3AJcHeQdoKBOksvuoR4DKuNaIn/VxwKEJUAhCqhmwNwu3El+kCEtBF
wv5zKRKdhRfo6mFyNPwzl/XhaqI9SaloGfkJv99alKDCcq11xgm6+MD/wGhiiiL/C8qrvS6m/HsW
+vYPvKr/85SRR2uhsJR5m1uQOf6Y53FzpWgKPthN5JdbGZnRpy0qIS2O7/YcKXxw/8C0cL/hnwxi
QMusr2lSc7pth9IUrDq2dDeKaD2SeGqk0eNu9cGC6MEnKKiB7+s/F84eqJy9dpnC0FnT/CK8s3mK
fdVwNHFQ7/9hUPrN+XfltOes4XJEU3AHS5ayYqwtbfP8QRr/IbRfV4CNgEa8CL1lkZx40Rvh//xA
V6+TDUirGyUuxc2qyFprWrU/vrmQYl3sIgnrWS70z00YWutfO72j8SESa8OP+1x5dSX7OvgmGemN
aH0P7nBbK20tP2PvQtDzDlLAhzqaLjTbOK+x0z42XDx4lxeDBDOwSpY1/Vl8QyVfXWevsE9YshFV
XtdrbUg4aJhJEgcFpcSF9UhjL8bnyqzmOB39Cn62SjXUie1/2689hqBkJIT23dcNRP0GxE4tfiis
dZ2rV2WXFqpr4RYviTdiB0iOU0TmZ6UPaLmie84x0KHukcIiMwYXDE7/hx1cVyWKsbxOeAH18aac
p1oGXURn8xp1fUgVbA+Yy2Iw8xZrspvEZYwlSSVT0gfFbuq3hI2AmoO5FZl/rQaEmx6v6iSkwk/P
ZUkK1BoNgtufQXUcvQ+E8qCgDL0eXeseI1fuNLlK2oRYTV3tZ/J+9IjAs0E/bnD34KhfUjGhCsr5
NdiebZdtxBIMrM8cwaCmplT0OuRbr/p2vuWrImJ8Ds3Zh9E2sRnskNEOtjuInIdmayo1TgsUTHGA
mvzEJs5EhHi28VTg0i60c7rQu9H8H7AhGEFnE/GuMWwqlK8RDJjTkfRA+NndZbeTzHD/jeSfu5Ee
ALvHHFU1Fxi+kWgtFYtw9spgxJAU9g6fXUEviW7X6453G7Sg1MZ38aLcwmY9xu07/wArQBLHbnTw
LWZbtwkaqlYU4aAWpjKwZC6ZzBV4buDI7w6zGSj6M5lxXZ2s4L13Rxicdq9p/WRyQ2VYZheR2KDJ
pVWoZJfdjGCzQL5LFPMPW0/WEKMiDx/B+Nlwbzb54Osdfci2PWZizf/oFHkxnMCQeFQC2KOID3qk
fp17kWjZVtLGPNAjJaQX1l9VC+kP8bdnLFVfe40jY+GTUVrTL99i9iE+PD7GQ9mi8Fq9AYUichjp
Ibgkd+KAXqlDHhqY7Cdh3PgPMhXKb8NSO6ge+k1XEW840goq1/sm1N7glYhSCubN4cDYsCkFIE0H
vUxISzhwWwqLGx9mlp5jlC7FQYH5gFnNYd0H+irTGvbQUkLoZG02yDXBTBq3IXQettq12/STZuwy
larbnrnnX1qEKQU0rNzyzaMba387fRsUkWsGrQcF3gf6K8Eg0F6Fd7PPErBHl8n8syLKS8P1wDYO
FBzMVrETuMn/+cVt/fgGuLKW+36SOZjsF9zSK0OLZXoC9G5KQfPATk4RvDgD4fhehmytjvdls22H
bbsnwPZCoLvky81NpffWjxiODiaklXhmVPN3PSh9LsUIwjvI6iVAUH2kfOiU2DgwpEUknNEeim37
0VMcRbwKcXmh2+y5nxsy/Zgj3cHP/0zh9zzuOS9TbiH3efd73bWn2CQ5hGo2DSwFhwo8HugMGKwf
bIfHTfCFLRvXx1sUyJFNTWiYSV8kbaenRPDN2+78EMr9KjZ/95X/cUCb4pECSYDCPi2cZwgdX34n
Gz+/jRcukv5Fo864lSa6o3LbNCDOYKBYqI2I5cpZgSlTgTZRQ+czmh65G9ROhx16ycIarLWQJp+f
FTseP6u3iCxuVJw1hKx3iiZPfm/BpuYcsaFUvhieVqxa8KargIt2Vx2ufzgapBn4oxOYeOrMrdv1
9iU609xw9o0DwuTH6uOnxynx6F/udDhmRPv2C538wX3UTkYIABMazJ+SRnaNwXLUNGk0PR8e+Kev
WYE9LD064Ri6O8mFialkUcc00AFJAF429Jrg8OSQ8hWXbFy+QXaA3//0b8L6DW5+Pfvs5fHS9if7
9t0ynL1rckaxq/cKRw1b2wX66sMycOjkaPljMXfS6/WaKrOMZZDn95fgtBR7tK4na4MVw4Csc7O4
cTkZQdlEPIhxa+dBeQK1pX3VmOuvMyY3cpVHrJjsfzeec9zZyLlwY0DhovcK7u9uqceL1WYZNh4r
PCjpdqwiDI4owATjC6j0xxHjrbeUxHaF8GZVRDCSbpBvPOc90nHR9l629GRlPBNSxyWjMr6Irrzq
OKR12zSr6pN91v3HcDN5iocLtrZ/pcVmbtR9M6wU6iHidimPTSbIhznG8fEBucwBETVrJS/u7Iky
CBoxf5NEFlYMWdtyzMFSa+X2Vz3YCIpIQC1FRddMuRbt2IxvTGzqNBcmth/3C2onQGVfcAjDHPjD
zc3b6kz/imkwXe924kYdSVbrrZtFH+eZEyzxNHt7DjgmurHiRHMWtm0N06BHa3LvQrcqyOnU69an
iu9cINzbrdjAS+MSh4Dsd2dwkFeXnYzRr4I8G+o34TO2Rivi2quVuQIqIxVW4vP9u2zY7UTZ+lgs
TWIk+5WwKDr1Ga6jbbjaiLn5Io1YMoGQwPRE0KGLjIqENkbyowftUJCi2CsQJjl1L3mfP3qarEzQ
Q/JYkLs7RPX8Chc9o9WR0jfGuNMS8OORHHFd25+rU5Q28LYUA4TBSsPFcgkAiARjWry25vg4JiXt
vK8K6hNArru0UwpHtq+zmUFdZ+04gsUrdZVqeI7se1cQ2syuTVRpvCrDKONLiddkFqJs1YyDDbU1
cC55rI1b+OPLTzzZP46TfXCNeTVt9ufW+qWcPYqtgv/Q+z5FMsj1PZEvC3NbQuWhUcicZz6pX2By
PkUBuKVE/8VAYphJWEA+Fh84vUCkCDTY9UJ9aA4WFotl9CpBkLM52WmX6relxAdjlUyUr9E06mXU
JswMyL1qP7Z4w8TxvZ19W1e9NQHNYZRJAIjnp9VZ/T6/J14C71s3Xmx12Y7exL8fQdVFIfxOfbQc
NSRXerGyIBT7DcPmRrvMETGbOPgjbuQnJG0Glaw2uXuqRnDBuLYW7R7IpEDj8oeMxvsDk/YkwDJ+
MaVmhuWBYUKYroNuU2FAFuH+7BVe3BA8bytPl8MdF47DfMyPf6o/23PoY3RSKLQ/YmtHGIxY59Ew
I5F3KhyUH6tNbLqi1r0Vw69/XfPIrVMv/JxZuNlUVc/JuMqlFazoOYoSEPNq8pOPErna87neBvdC
LUIMvYWM1/Y5ydE0wI/cP7iO5x2HxtDtziCPMlfEB5N51o2eSJ2Vy3aViTUHg6Ai2A7384NcSlbA
sy6st5Mnisx0tDpst3SlXToSGn3DHpyOtNN5q7ZGDUCHba+mlz9VnwQONwrMDuOhmXuW++O+Ieuo
HFIzJcTtwsz2igNBv95eqhEHLlFsIk1vL80RLf+wjJZMj+vK3TtPY8JCUNwKjTklmzesGNqCbcHM
NuLwCxAxdCTXL6M6qkjKMRC0Y82NHNQ4FF1qBl0xVSJU/MK3YoYm+Wvb4IeNxitQrN1kmT87x+qC
qywsFf53/PhNOGIQ75zhhKu/LOMIvqMApIja28nQVo9qhEJwKm747OWLGlFQG0cGzamlTaA9HXKf
3mQqGKqebae96QB5ispLJ54TN1xk3lScXWk+oXoc/bzEBPKzOKmVQRC5xAcUTks3T3EhrAFb3tY4
7J8jFr2REnwxel5J4Bw98csQgKe/z0IpD+dXAbg7URAzEoJ9QdbmB/VZDH+yDDFGDqxMQZJmg/a8
IFSvPI9gGDzdJFbjDxsOP0xXLd3+XlDbpL3JgytnCUWL9ar6NRnkrlWvYQnngJFJUGPclG1OoN4s
IvAzSk01Cq/6AFTVU+nNg0MNPm09MniWdB4sEv7Tnao7eUH4b4G0LelnE9+/6uPLM8/aVAt3FEDw
jL4eZ0u284frfm5CGqD1UJLK3wwssYu7qRg8uaDmAk6+d90DlVXfJI2Sh5YNeCOyx4YefAIF/5AE
LQxqfbtCZqyS31skv+fRxbQr2xEL0uBmJoOod180ekbWM184SeTahZP37elq3T64EIt9cm8Ei1lk
E2ZRuQ9dbquCBNvJ3BqaQK4QmQlyXWZ8ZlAfMv+LE8CZO98v1pNx0dgOovmJQQigEIrcp7Z3hWq0
crQIrmxFUwwx/2VfE1J8XCuX2dkIBBBImg8RYmTXQBaluW/cFjevFI5Eds4R6VjizMkSyH8e/rQ1
H34qMmmLpnZNApEaa7o0KjfoVXxokFXyrmg+Y8IZo8JGuwTPZjULwzvcvYmPt9O7IIQT0mRrsGXL
t3aJFNf88cXUdjBJe9w2IG9qCW168SRon/JFwNfjImPUrReJyrivQ/pIkbFSdDWkoGV1rM4tlkEw
5aboA3hYHZM6/qvjJ4mCAfPLgnhGFOrrWyBUQ0oIiHJ9m6ohXpaH3GMhO/S9utGDkWABRUuJJSWR
lzPgO7lWZ1zTypjowRVLd9IaGKjswzLL1jtXvlEfAQ97g6X7rRHYTo9WvcEtILjpyhgd7W9vc5uS
DmPiZ4K9f1NBH2DVpPMcUWQG0zu3a3rdHsbRhCafMHzp8rakcPBaFVuoFIYKmDCCVrAxtLyx6K7d
c5FAZNrQABeDIYa4LsE5QaweOD0HkH95A2cTtDTjeZcZqJmUQP61pNc4XdKafFrwdMQaO3GpczD9
kGbg2U0FaY4nd6YTBm/2Fmg6TEDKDR1N5sXtLYwsQCxZs3F1Z44kycjxedBGmaIrPNmTq697Dmzs
Ny1db7NhwKJ60VpXxUhFBV78QQsxuuZQPua9TyMJg9ihNt5HGTX+zX4MozcJuGe+Om/CXbtsuUpP
V/cDbvlv2AODXFS4sjeiIZkPKwpF2T4j7hyZXWcURoRRH6VcLdE/hM8BMAHJVNaF8F2ibTen3lOC
ZbyXVecpBiekZ4jfuEK4XSujYf3RXGlg64J/v4YHlqcKe2Ghu6hMKTKpYGLg/FqRhDOqcwZ0tOBR
6frRmG7zwx6d1vSv0sT50NGcnumgPE4aVUJlpH3gsUBWDSdtalw1mfJI2K/xbfDQZSOsUBNAjhZz
Q67ZWCRKb8CJMuIpmqvM0VdSSQT3W+1AnGmwQEgibalBeFMAVBgX/RETWy0Rk/POWoaCwD4iScEw
yvZsnbAWF/+IxNwIMEL0i4iD+ijEAg6pjbCjVzgcY/iPKrxMOlAa93dyHZGtsP5qhhAOZDuklA8b
eBihGj0/zC0VWQ/Ay+MikLYUA5zYFGuoYXrGumz9hyHgtteXzF6ESDYtUQo5H2kzWWjqiOiHnj6S
wZJXTmsdyd+IgVaWx+H8brtHLWqFZdN/MYZq+uhrgYpUIrqKFsNiSPrdmK3i3rBILutlZuwseoen
unJgA8o8kFsIdGVH8q/uVBZFkF3amELSvdx4AlwcMa2cqkUWFjTfQZ/qGOKMGcgdIyzC7uxsAtp4
BSoX1cdIto0/Tq5eQLc4uN0yyucsm/+npiD8YvijfY7Ps5Drr0zNk87tLp6qcotIHuARkJCzZmjS
PIUMtysTe0SfPnmLPmzDgjrgixNPRUi6qPRZ9v/2962ETR0JfQrLmgA4Ads4hy4eN2vUc6wRxIFe
G6WMxQTd6LkAEZreJrabw9KAEqwHTFInuVc4bNRPAeU0BET0D6GCsyjcgyJakpqkkVHxQwX4LJ9O
a/6qFPzvbXok7rCOIVPBp1lCvSgvP5/wNm2KyW6NnYgkBB6t5VceuOS6bcqYWpDOh63zGCVku9Vj
rDjnYHAzcTRSSwW2Lr/Sx1c6VjGn/wa9Ri8K4NkzGvNPzbnv7VNpO0l9goFkud/G+ftG1VyL2yt4
KoQRXOKSi70EREULmnx3dhlKOZnlYYNscdedxRhQR7h/MCawY2YdAzMtpQK4NiqBfczb8BNmVCjm
w0XczV1E8t8/JgJryaXKP3AJImADQwNVvfKBr1wPXGBvxAXMsNRuEbfa03eLnHpRD5uHslka1qLh
dDrk4kmzkRbe/YFABo/hdJfnktJ96MnNlTe+oksErpOKkCzWF1a+1E+8D3NF9pWTkcCD6scuUvjR
D6Rs+jGsl/TPYrMs07dnUB7CYXknTmcUFRIUihVGvhYS9UqSbecCEJlRz68GS2KLpGiaEQl4joym
sQHuIPuzT06MrtahzaCX5Jjln8Ve0Q3x9oOo+gVUfmO8I6tWB81MaOtQ6cFKo1TW2djf4jOSoAul
Tj2jP3kFH4hL0Mu4/M7ciq26hhHDztcJMzYCWKSFTiNg2vOcdVJaw4tj4JT86ZF5I/rly+o1zQlS
PQKLuMMRotJ3461EgPNNegtfnJv19p99DSRGdACfWLEumZ4BMrWouJd+zK2deO+jLfNpPxQiDeyv
GJkALEWDJXka0jAJpgC5KjdQ0b2YCE3hbvIUi7pqJM70uLoEvFBU6pcrhtZlAtX7KnZ3h0pyLVGR
Bd3n8U7OYAmN0X5hqE4U/OERjOWevqrmGbqqAw6A2rxhJ358IhcD9LduvuGLPvkqG3Jjq8LW6+Uv
jllMVl9BbYKVoOtBaMIm95JoJIgnQTUWdrGfcncaL2nscV/qgdRgYKcE4gdgnaR8MSzEV8fHN6YG
tzFXwDF2QV+i38z45Pg+nmhsmfh2yXoB8S73wmarMeRp0C09NOXuZ3qCiWBx7i/7tII9S6qS9jeE
xTWmZwis8FnITp8UgoOXo9cv1Ii1NvJjBmw+RCoruXzqGWP+Ho3A4zyc96yINaHM/8yw6GJp4UJp
QJQWC8BQb8mlgfeuYLba1hvVkNw7mDF+iUm/BKF5LqC6JEUSqvYYcwEZUN2U2t4CbJfJlf3eLfiu
6RLs7jvyY8ke+RSjieQPq0cDOAJs8KU3fK8Xx/ynEb8zf7c/oXh/JbXbUdkzRoQfJlFkA9d0jlkx
WDPP77oraUU5QkdwnqTdmE+JICZuCMXJqSYqBSp2beCSYXTcVZ+jwyzs4wLYDxbCBDuvjZlfD5TF
I2sSfF6E8y0Vw0ISdgNcJlC818/wx09jAJesLDU6AB4v8+CnlHL8ovJfNJLtjQeLuM8M77docuWx
JJXCRlshVCZWjRW9J9HCCUzA+5k6w22JIfB77B1WCisvCUhm5LlefUJLfbExU/AFkUTNYNhDzuM7
V/4he3QFnttpGwMsx5Jo1a2SSOs55ucuKjB9cL/py53certGNebfc8o5BJd+Nh2byC7wPDJSrNya
Zc+xEDdB3nPomFHMzfWopet4rnm+D/eFfer9RCLsqIqS1iPjkM8rMymwopgWP6Jwo9AMREo9Oa7Y
9v5HWNDCe28Ettfn3kJLuevteRYsdRwHJHNQrxd4lJyStdUCFbkEtw85LsIq6qeoQmjcoHXIZLjM
h7jAVssSjs5fPzO2b/gxJgKuQ9fhlH/gy3XmcYh0jaxdwPFZ0hyD3mpkUxwC4uCzQiai7TDh8/Zt
EYKPahjQpo/Su1Mc2oab43XiDfWy5vMc+Gcc/xRKR4vkzu2iswdkxVa0ga8w4AXuuXUAegvbDuFq
zq8BViYjpgDeXZsP0uU+grdGxWue6I3LoboGX5rxhoHOKYSfNxGtkbsP7CxFMLcoSqeVQ7934jln
fyNt+cs/eSNOdRu5ptINFkQ2oZXX0qRyZTsrO2tW9OgLjyFKNig8fV+gW2daLmfkqF5aHJY7jM5H
gQ2z0MqdCYfkp/7lFR+xIy4nVYdZ0G7krSlDfPjy0fE79Cc67xaL8CudrTPORy1Gs9BBlTynfIr0
tfcd8Cr6W3Frt/ESTfpuvFaV0imFXc3Z2JZTewZJkpQTsYnChbUtpZuQnkh9CE5hugPzmRV+SQD+
n4K6QQRg+VkaQ7kQ0bvrAqHTMynX2+XYQBE3FfkcGmfQYn92IJgFP8wiJ1ts/ZWau1vljX6whDKZ
xcSjbZo/pB9EoxPRbeHzLUC7ebqauynuQm3HWFJm9pVLFh6oOqLChHgLe0Qirewqo17ElSzXoSCF
x5lcx3wXRvYOHBDIEip/m/ZvAl1AOj/6pYG9/I+bYJlpYS2U53B1a6FJ1WNjbRpWbT5yGkOW3MSZ
NOcPpTeDXaw0Nw7F6NSjuv5SgHmUwhxapyU5fhA/7npGswo6et06TfTIHsqi0Vy0p3Talg2z4ggf
vw0n+1TU9T5LobcpBgHr2/G1QukhoZ+wCzW1R5u6O8npO4uPA/KyXWP1KdmItIMQgtYoiYAMC+xt
6FOwB5HK8Bb2ZoPej52k+1cQJflIpWo4LcXURLvX0lMDFhqXL8iteAp3H28Booqo6FpHblmgiEXy
3oMuoF2W/NIv7twASQcd4GdWjrwpoyDol/Ei9Pj8yMtAmQyeAQ7J/7Gznj0+SaFWsiJdINJgInM7
GRrbYwmjyc1g7A/+op6MEhCDJ5//dij+hy1RZXTKL4NLf4fz3VcZCprFts+lEO8JuvRY9kGHq9D/
F12+eXebFi+g2pfS+Bnmno/lwz6aD37EFGSQd2263pU5lH/jl+war8HU8gBcVUjpvKY3oXxYgd5Q
cx1dYfZaDELYEjtM983MZGMCLcEjGlLCXZXhrQMEmo4XHA4S8OhJV5HS6O5M4h6nJjam4YSpGXW3
XUEWVLlzWX+WNPqNwtnCxdt3YZ0cPhQdzomhPYBeRlDeiJpZ/VcXcBNZrXQbyz2THmE5H1CzT1SJ
qDKTi+Edli+HkipUW/N+md47JXyerpEBENhgDwtqWcS7ZK095iIL+P7sdk5v/itDTGHyzyn9JStx
oAiJPXMpDvvzGovvWIHgSQPYRNrLwOd0XCuGbXq3Ouf0xkrIEtX2ZHcAclB55uld7t0t2AeZg0m0
kk8awjdH0sZnUUwR9Q71y91ze8mxxt5s9kYzTgRBls06dzQhFxWQ1E9OWOVQ3BFcAdQ8KljL41k8
uSN9kmUZa7uQrm/ZgE516cOO16rZn5RCOaRHB+8/Pzsvk+FRe9BLqx5KHLyAGq2XN4V9vMgAKahB
ldCwCBwMpL8XQlg5FhOlEgvjJ378jWS4JsmE+chQz6wRqTIci1yBJEl7XfTAKNkW7YkvM7OWW6dr
IsT3lLBmedGNgkrbe4Y5RwAyVbKJ8Eq7xfkm810ROOK7/FUFabVPGLExCGzSZE5VFtS7RTgdIX/7
GLzeKVTXojnCPtPxloEX5CbCJhEBv2A1rwUHzCSO+8gCtyHEsIwdRGH/33N91DQ3ITB91UK0syU/
fbortEtDCfHqrs5X4JCh7rPHayIJ7r0UfhGS59sfIpQWGOyGMou9n4sr/IHccO2s3IZnmNeKas2S
rooiz7tMfh9L3UTEb6LUyEwBsVQ8FMg2rWLkPLJWh3EyjeBwyNHZCrkvx5nTYpFAQSGdeoCQnGQ5
IzmfbRo42kJ4ThalwKByD23E4i4x4CtMXLxYE96N6QuRqXq5b4voiZYQo8w+uqFK2ZElI2O2n6rc
G4RcdGwF+DY6s4gt4uV3zVFP++R7Lv5Kw5++OzhkQeS66v5/bczlKxGd8BoCg83r0KCWlm1XJ96F
LdY2rlRuD+k+OFDU/x0aB8aw0ruHoIZNoYLIWUxvryAuvwm2wSq6abVDtq5usL8IxH5UqqDQpCGF
+TJ6FVCn8HWQpfHz+nALoek+E5Xx6YYRL9WhhuTrKb7InskogaMqbwaH3PUdECo8zlcn2tk51EvN
Xzr94EEhF7FlUr0XI6BpRFcj6Cw9Gxqvq8K1oyarAr2xcS4gxHUca4X6NnqORniMwxB97Z6mk4/I
vkmuqOeG094OWJdXJ2PLmrJZ3j8/5DDD+twVJJ6u1W2Pw/wSKf4Pu7ge0GqPW4cDbTw6EV3ILgZp
3xL7ge78dDLCuKeilo0+N8Sek0RDp0clguvFSTDxpuNzBECk+9dk9td3sImM91oRTiQ5/lOwLbCk
E4Lj6EaXh6KDdcGHN5Is7Jfqvo2NTHancQcNNHtn8VhltTLXfXc6GJjY3MQzi5I/tqcGz1jIj3zr
wR4fTNmkH5sI9j/FvRcTGXPogIVYLjTcrKkMV+zlnwNs8Mx3kt0M75VyJVJiZm+rYaUc5FXRE3DF
S4k//z2O4dhZs8qvDPDlnURbA33ZiNkKc7wbql/rBljgfuq5FflbAfz0kzcvsXmEmFQWD6mvX0xg
ZcJBvuGPVLabfu17W4ZTfcSSPA/2bxrqPmeMg1h4sYzvqFi554raTdVLsilHBgoMdIoLiDIIiyOf
+PTM0IKmULphe49ULyfNfpIOvymW3LPMJ6psBq0wT1+mkglAASiu66/udffqBANrLVOvjv6s90Sh
fRZ6hOgwUyLNRgaKBuxwhQE9pPzkslD95UvRjg++5eJGo9vjs1qpXFb/+XDuZ2kaIeN3lU7l8woR
MpRgZ08jg/STAwnbWZ2Kkbkks/SYYMs5ycPLzyudvreegjxduF4sFX7fwgNALiLz0ZxzXdld7iPq
5Co6FBJ1mcIjtaQHA3+xCfRT3enYhEDB4pp51iNKkyEq+5N/lsvxoPPww6iGoplJHqK5UNZi/ewl
h1FwKlvfxIbfvpc3vm26q3D/89h52Ju6scWJNF2TpQk7qUuVx0iYBs0q8oQJ5wwI/2cPAdJM8K37
Yshmka24Gmdqtcz8507PW0kqvg5RP+FYgMUytAWQVJc6RwziGO2nF7tVZGyGLdPHV4jNR6/Ws4ex
JnDzjZEczlAW3ole3l04wBBxRKxGAXl4cjvEP6Py7wKjskK8k3BkJYnUoktM5RFgf8o+i2rr8ny9
2yQc8+6r9eh/UNjpmo12F6LO/Am4pGIl31FosfGs0+dtJ6tTO5Wf7Ks4Sn6Gf07IwzOozmKAACW3
nqjBQzZGSMYypSXvaKbNJtvtAn7iLxgHn4CmDNDDSn+/iY1b1gE6blhoKNXgPKMdhbsXtbGc/X5L
B0MOzCI01kGY3i9JIu2XOEFadAWymmokGUyuRQAbtHJqEsryDg/oGsicVcgkcJiI2mxIzEsRgREm
XLiNn14/mg4DMh48QFhxGcJxMASPELDGulR0z7EhFxydtx/VvvUEue4Fv3KkZFd2R0pIxOzuRQo4
UauZMZtft+Ob2tn8X5Wjlu5tpwbeTGxPZ05oEHq+/gxSQmgYw9tO//pijA+QTbIM10rxuZQVeKzw
wpOA1TcISPe5T2NgHzte9+Di68sGjZm152hN7JKuRHLWNY7rG9nAX7zDr0BIioQoqF4awaynuaV5
Fwbz4hLuM+RVaKlk00LFHxtlLQSxlAfCsjotNvsN2gMWoxwo9P2nxd38N6KXNwqf9t3Y0aBZU94u
bFYuFlPjMTDgBYpdpz2RCRLsSDkgp1ooM74AIgbUAbg++dqw+DVKUxQuyQ5hcWWzsWiRScE9xJfN
xIDplwdtQBuYiMoMxkB9mlW9rPShDbhCnhQsVE2froXtsRIilLFOALwivc/FuP50TLIJ7Jpm69F8
sA+my9+Fnf0mtQ6+OL7mmB6pLwfpweMr3e1v1o0sIxSpb/JT30evQVenh9ToLyW3Mw8Bn5nKdJ6Y
8YPvX69t4qNsorvzt7Qs2yMmrkJhATbbSEZmonozjJxR8S/OJM71aF3TfVrwrrS3bQ0210awjZiH
z2gfnu7l9q6gd2V0O+4vbQHIdEreEmp1X4ct0zrhZ9S6E2yiAvk9ooyI3yAjloih9lx9n5gZEa6H
DS0zPtxe0MJC3hP+JTgk2BLvUfnahDpYxqSGNmYH/YB6516WN2Gqt6fmRr4ESZD1/2h/aLTLP10y
Lm8spwLbHmFgq0SQIT8btGm8nxFXhU5r2UmAVkWMF+ObA0aRl8vqiKQM02fq04+jZAVBrmY98Drb
zVF7UqaC4yguYo/jbkW2P+Fh1F2hq0W7bs1N0Igk71o4OqhwGcvZh0y3eBAkFEXvMwV5GkUfWuTB
ewhhPjAB1ZFl0DhFtXJ/xXIpa5R2Xr/yse3Fu9wCt4+R6E8sCBVyistQcBypTnHAaoQJrbyD2w1V
tjuYuI5nw9gqqLcCWXwqhBPQOH1gxPAUFwze/6X1CfoABqiWQAA5ebQI0xPoYRS6uXxFrfTyiM01
z+LwGkqm0X5iPgS+Yfh8AuBpFqnEj6tj5QC9PR5xzaPvwn3Om15qUQwefFziuAuGg7lnOgf0bUKS
cIRrLxGpxZje/yuY4aM/GHGVxGMUNwYmloJ3M9aAExphqSHCsED+poNkbkwWDbkNZU1J4+xwxKlE
6xpW6Let4q4OUVbrmFbRudzVibmdSGYTOtbcmbS5Kg2wB4X7I7mImzrLdAS1S/veBILNPrQGkxMb
tOz1sqNzRg16R44PwPeO17SKJctWa42tQNDydee6+fSyWmtFjG2ph3zcJ5fM2IGbJDmiOIu1tI2B
lh6YIUmR4F3idf0cFr6LZz+PjrfTo09hFL2n604jvMWzsj4GP/syn5RPeYjQeolN8f+WYFMAxH+W
YIus5yT1oIhLg/ZCPUybnAb8fpDk/MgXeVnVrZokMirJBoOVm8pzAu/8gN1levXd8tZVbKKcwEKf
jb80/XLvE3VQbpUigG8o+zkdoEm64/BoB6nk4Hc6Yb42lsr3l5aNW7jCf/4goAbx3gtwv4Nm2Svn
6InKzB6ME5ck+4NzrupAk6axQ37AzzlGRv0N5MZmZGcS0rahrAAwUFwD7OSh2vF1MtEDWwHcqrnx
29mUKU4ZQ7s4jwDwq/p/V+mUCNPFgF1hnmQAEnq5TUbWG34zlAftwA93oWKCrl60tzGJl0JlD/tI
org2G9r9fwFSyzXan5zdk6q3Dkq4yEWKGtAR/OFqFXcLYpH03NUfF8SzITROpuCzhyUYl6rZ9TSp
N0C09oLKwuv7+fK4Yo93R7Ss4onq0jdldBSvrDm7VkRmtADrwzSvjzM2Gfg/NzFLbr2QtWc+muis
bMOJhzFOoTCCgMcGFucwJczQFzWB72eh+U+fy5uO/2bthvsxEQ91tFpjE9HVqv5AA9u+Hkh2glyv
kir3nqAyaKaFXOs1tBkhhvWL2VpWj3IUTEuZ70YG24bnqYB3aaWgyVHZ8HDzZhi4aPCQCYBInODn
lqBp0gpynZVYuTnnmi4oFLraec4h7nue3xJpPZXEpFjuEnVFWInSE2w0dp4y31gpbtbLWXX3ntm/
G5Goc0JbAl+pUz97DoT+FkQK4fIM4FboL9URCltVpkqFUzJ/0w3s7aJHEtX4ModJAFgs+6ZpI6JT
7hoBsdEABcRlHfLDBkmv84OwmbXei0PzxvpmT5D3DGoiSvrp3qt2NUUPUwGhFethZT5W7whB0Y8V
SSE5VBI7cn/ZqcGDxBx4kVRC4AzRs5s7NAEnXvRifyEnVXmQJ4yZr6eziPTLlw5dhbXsLacIsNYP
bgZSDnn6lLkOlI5RvEYyNsxaSY2B8HNdEpElgmHYBSsJSceH9yvtRdCy9Qbw72UuX9+kPn5EgA4b
DjKfiigzOxWdKpn0HcDVNwoU1hWic6KpNs2zZnYozvcXgQ3OvGqrB0VDPghU7w3bMPhFPBbc1mYw
zTKAc64tsZzjYvj7cAfygcWePv6VL0H/IWsrOSUbSZ18MA4GuK8ZaPcuhD1hOPoMlzGE4gGyvDmx
/MNEN65MOcbuZql6x7aWVr+aBhm2vwbmtY2HnKxzDz926zLw0CHH2oM+wYdexR3jE+X9x5fYaJtz
/1EXNlVdF20DiQhg7ZmeQ+5g47P4A5o+tmDMjg6OYXdz2T3l0xGvwinla0e1DGe6Ge5gK41OmIMl
gd6XMCRxqGbZ3EQxpO4ZJfXu0T+/keFaV0E0yPFbMBD/5dGKVVSV2dTjEqyXyLcqmw+B1JLD8b5f
CfRsf+3Mh9Q1YNX76dADcabRw879RHr8N2v8NOq8ZhmbvOqp3cBLwFGWnKgAWIq7Iel1AcYTkTaD
q1d6Ky0TSeOHku6cOq6p5BEQkgPBeg786RBmXspMqyGjIchdUwhgBAouOKyBVeDx7ege3KlxH7t1
WpZnUL21zbqDTK5HIGiGAbHVjvU6EmRIDQme/x4fCl/o4ZgdU90Yz/LyoobCDnEAP1/Ft9V5A2wG
7y2zm4DeNQiwvaw7ZFLmbX6gvaiAO1d7jqZmNGoUTZmYGZomaTNO8sFiLN3YGCcnYeWnW+475rwn
QYyE1HYJ4Z0mKmab4Q3EvI8iarATzf6RIjh9Amh6JiLRCKXOwIfzBADBwmryibKepoQJNRLVBCtC
iAsqRijaKLF+PR9hDiIGarH2nIxQ0oUsslQ9NApm+SIGiUsFHPfjfNTkdVGckSKMyngWvyCggQGy
yJE96wG0ERrl23uNe8qhp5tsitwjT9kJhfWoqGF78AG3bAfW6FrQqbL1nHisxoSFOE6e3j3joLSE
+M5SzPlLsOp3xKoDwPnQcl1DWCRThoJCy34Y9/v9GfC9O7e6IOnE4Y7iKB2utcX4o5VUdsuUGcKm
zY6p9G0DC/y5iHAX66MSv5r8a05wTh1t9ASzhA82lYwjpLShqwkDoMKzW6qOmgs+C4Cbj0nnreMy
wqeQzcpWVUj0sh6fdmWWJFbvCMZ95INAmjOnj63eFDPzquaF/DWMlkwdBTnrTSr9zAftWi13WFbw
FeiPOSixYN02fD0EuCUGgtj1mIiqUF++IW4ElUq989rB/Imhd+iPsQl7tWZ4PyL3s/0B1UNkpBf0
I8djmkLk2GnUgvkNKS/vs5KEGbwbqUO3fHq4/6cWtfbNpO8Y5OWF/9Ov055vi4WsxDNldsw8i8QJ
xIHU9i6dryVnAx9o7ZYFC2DlG5KlXY3yzVLdGToOk7mHErFAEBNT7+3aU7Tu+i3E4N4r3xLpSGmp
EL+z1JkZILjnTXcf5cVMf5AJSKMPCpmrjNWCxVKy0eoiw1IpHOptgZLzTcDJ3b0re9rV/MX1GUNd
5/3cfx+lESNLynqJp+K6/cNYdWpTJBQKXgNh3o0UC/0kkF4P/Dc1RlkaMwq1rzLQWr2ELEgE3H3e
kMb6EJ822vLbEQUOF0lRetcYByZWXMcxtqHgSNFMI/fKnqpw2z0c8mhH1wt2Ii3r5hq1KSG3enJm
NKcjZ1CH8PKuXhftXROkKt7LoHcDP6RqgbBw9aKT8IrtrD9JuLe8BHpribSCMp6PZEkniFLzjXeh
Moc53z+Fyn9YeNDzKh7gKX8XAbeiIRjXtU7Inl4YyJTts0dTnyGk48uPRm5vC6TWJ/XlH8iaYl2K
hIbGm+PsPa8BZY1Z5XlFtZA1J1jHf1cqWEZZnFBDXM67Nqqb8kOu4o451k/bmzzG31ZtUJdmqCGE
ldVij1BXS2+hr6/LOl18vYr03VboS71pxpDVpjG/lK1QycphvXs+ep5g9fRuDOvvQH1FXPxBjwRr
xuqrQXHY4hS57ZWPspT1adeONgQhT3siGAQ8oZlIS+hdz040940lxvLOH40mksDsIym0cAL4A/dx
0qqWGHavUOVXMVUfsLGF875NDkBTOeG6PLTVhugO9F2eYXxhmd1AW8Ufe0axQq8o8znDWz/oY8Cr
l99wcF9P6GepaHPWABZW13LXrTfC8NJ+a6Mi5hxiDWgMjyHSWl6p427j1O/Ojb3dHdxtyergeT74
XvsivcDnjzY+k4rJDdYe4rNdii2bnfwWyWd/5PMWRcTQ4skK84SuwL5+8q9jubPdMviLkX9EjzaZ
P9EPOQh21/oZEpuJ99dR49SWx4qco0TKrcHIfBwpyXJdxcRBE2vgyEvz1u9OtNLrPUY8ZlBvJaVz
xMxhhfKKx1cE7+RMWBsVQxP/egHjqBunH+AZJNjwkKBxJV87tN853kD5Oj90JNZUb6g2FThqRJx8
/TecnglOO2F9zm63JJreZ76XWl/Gi+24P5jFht6QcQRimWlb8uIeBK8EUG5adiwcMU04013OTgYO
twTCbBMUYWNmU10xz61aZUVF2TJad5o9a19UDVIOU98U8LidK9qy3Aw4ynsRl5X8dt+U6zMM5wBN
+m79sq/5b5S+fok7PnBlK24DSBorcT846ftO3fYwuq3LdTRQTmDzRQZAcl61osgkkbNcIN5AQUkm
5SkDt8jOo4tg/1sNA5JtpMgzu6hg42/BEyhPmksx2+cLvFCWV7O6QOQNfxXxjevwPU0yNHegPjC0
zNssEfXxmsXITgDENpz2RMarhYT8O1AmqTuAwy+quTZ8GTH8iGcyeoPqKPagPbzInD8LB9EP3dAl
asqUMw08sCQ8E1r/upDlnmBjeVbNJsQCQ1K8DOFiQhLbIyejUGbuOh3B/sGZ7gZi8yxoayg35klN
QDtgEVkGhisd9hG3dAPFBWhpo7bNeyREJK5Z0h7grYGAHRBS03GiRPXRp3LmsnQqr5egqTuy8dap
Nq3dUcazTVz3pJfMqEkzFemVXfKxBuCtZimJe8s85beSc3HE5cLT6rKjsHRK6JguRpS8K1TOpnGd
cgXVZ4zJWKG15SaHe64NZTtICdaiH5f+sc/axmuz1cYRlH8Znpvv9w8vvQtgnd+CtqAoDkCXtWiO
L4VHVZyCJoK4D0CB9Aat9ki9EtfKmw68DyU7Q6B5Tv498m/WMT2Q4n+1MWO74L//NoygGbTXk07U
9/IyfiFMf4EZEGQs31B7cUksu5NCagxsguwtSHoFhw0JO6XkZAxLZutgxhbHcHHp/JsXVfJjdXYb
ZkDhG5yxFWH9oB2IjGA0qGg2bMj6+KY2V73INK+M87rA3xi4jp6DdpmtBiDSM/gVxfpqk6W/2mxL
dolC4tV8uJnBAqffdXjyiEgDu7PBG4J81ZNB3uaGBIpjN48fAhieHWRqUofhzs7JMBXoI1Oshwl5
I0xy9DQ0KsA7OYWssKxyI0qmNaxFh1+qSupMslP251XLC+9FbvqKqZNIgQmGZQBhC7qwzmPL404J
CmREwKcTIgmJOe7nmeke7Xdr2fGrGf4M3tRouKgcv5+6t3y7GT2PPxjhVrpQXtdyvxHlt2kGjBvz
XmLu3za7VeMM9r6c5myse19Q53O4cZMukb4tmpJ4FMyIpU3r26MkN9J0pRbn3xlmCIXoBXbEIVjV
epC6tQe2JbnyP3TymWOk7Wgf/Yw5TyLF+vOZRGuw3gbaVRl4BfdgKSk4m5RuTkqa8WLr3bicFtL2
ZiGfnNeY0Y55w4s0+6J+nAhHmYjhzE9W4UFU8kz+vu/L6yqixyck1la0ylsKH86Gr/ePe5EpEX1/
L7MYzJKpRtq5l02MT+4v2BXas3tC2DDMnHSek81ferkV5gF+oZlGdGGjYL5j3Ia0xl6a5vwftILY
gYkhfeGNxwZUEaYQparzkYzTe1nbSf8C0CGnlrg/c1AAyAiPhTdG4HTls04J4Np5kAzU8t1MrfoL
+4bUoi0eQ4CXRW03+9Gw8onGmyCBzXMA9VL7Lem4y284ao7GzUVqgmtNqvkmEEKKWy4grPY2pMyH
g2BDNkCrCVlvIQ4cYEu4AXoxTLcTVf/3cFS15VIzhxekdb4sLamZNnQWK7F+8jTotyrnAcT7p1Yp
ogpZqrq9BWMmZQVg2iSlcw9TEBLMZU2nqsf7IKRy+0Vysel5X+N0N8Btw1qSAPXvDqByomiZMVRc
Q0hQubdXeVWWA8bFH6B3laNbeMTz2P1GKA0Us+pCd7tjICxvYIifyV0S5eURM6ngTlDD4KpbjW2D
6I+8fGrDVn4QsEyHKazUJSIz3OcDFlnU95ghrU/Ajs/FNmPaKRzSBQ6AyJ0Iimo6Orm1VO0DOhnz
4tYRsJmCndkVeabNQ1ir4j0EIi/FkAFza0M+aex1D/pCf54DpH/zgumixuwaiuZ1P628r/VYf03B
gBzNmopdBi9nopDJzsnm+mk5pcdwWb5CKYusSP1hF0V8Deyd3qwiEHWVbm/lRRuVNWGIurhPbHaW
zv3ng7ZKaVzoWNb9UB3iStiBSB2Q3osFgkJC2D/Phaa9jYd+SSnne3+hJx+zVFSS3iOB8eQSKO2v
KXhjQ/4Ea/tlaa0Ix73RiZnc4g1nTu7F7vrv2TJBMU0r0IyCpxhxitCA6i6PBFrtCe4XC4K/4TIX
zJn7fjfwEMd5w7DhfOb2ojKMcWgEXVDNhuvfEu5sqoj29d1W2PvYzYnzSXPx1r+hGah6jkkI3BTC
7aejyGGIy/NZAj4SX3MYempoGzQ9MdENVh0PKyDVriXLYctt/dod2sDwkR9SMR4AW5gBWu4z07E4
XebCXBj2FdNFTELtiul8gGArr8coKcRiqBWJHVeDhqOYhqojvmfai6I9G/nJJr1jvS1B0wzRFMuM
Pl/cgZ2t/3rPUg+lz1bovu1Ff31WsAx8LFkzWRJ0MdoO0zTJHEsr2IiIJjz/bNBhSQd32kSop+GR
OFpfYoam/8NA5CDQo6WXkMkUXsrRMnBcLZpKQQ8Ph4SuvLYsxBjB6fteot/6IIv5yTbIONeWN0rm
6zbgOHGMCcqEITfct4+LzPRoWAsQCj4jwaecfeKsLKKv5Ssrsz04wxKMaddXqO2Aeq3OUXJlIeL3
e+4M7tYzYZKAUAFoV3BXzCIvab8b9R2bwajlLpN8l5l2F91pQZcynA7KPfmAhL4p4fjsjETB7ppO
yfTOaiKRwv5SmYsb+HIALoantp7S8CUNsXST2vnXfZihNQU7L65Vto8lrmjYIUnqTimh0eG2ldGG
nm2tEDT6wOxmfC5B9+UJ7NoWIFxv0nrgUdOkK2mWTxo4Pp+K0BQiOzQ9Kvu5U5nvu03VYKohMuQ7
n8xgVGeTCcn2nZij0Zpj8ErUgRDPmdEvQ6CsEEIFomfhceA7Xn5PQYxKnHmwZo7xIhlkZvTeWkmm
x+vnmwVD+kucUv/bw0EtCofwHu80Ywr5f1/KBkaFNAgokAhdkQLYAxLgo7cS9cxl08ITXDzedvVh
UqP28dyeFEGn56JmTIpzqYSkFkFUwSFm+7d1k9jXkjTgYKlkq2rUNEjN36T/gsXii0g3bXcYs+ur
P2+9VDke7/EwGflEzqahXAtRjAxJa1+1z6qHG2qFTpVlGM1eiwETzr74FZDyfACcOa1buugixl++
7l4EvBuPzRpvRds+Lg1bE7a/ej4AmHZZApI8ScqA4LI1PyNXd72TILc40gNAPDO6x8QaHF/VZrZP
IPmH7UDEWOpAEGdq6d0p9uc7pE9k9l5oIqzKJfjV07kRIwkxP1b7RIm01+9NNmiIpSkiTq3s4VI5
poailBUt8yeEFeVPJFxn92mRbk2E+uk8Uo0cgCyHDVrpft/JAg/JkO/FwMxX1gMu7aeESfnRr+7r
DZO6JAwKqj64qnsuTJDsJAlsk+rmdxqRDWJVTV5q2gOQw5zBujsqLXcyio60uZuG8Oj8EruNacoT
1zhCdYR6GuCzQrrNKL+dB3jjQrXS1KwIHBdf3fOtkC0CoeOlE+WNWnbgKeMXsq9huyHX6v6R/0GF
fILlFJr/St/4XGAjuMbLbBdIbrSAQEZbJA5Do2vX5KiYsuZKQgNtam4Ja+JmtJtV2sbbl1XPS3P0
36QLItM3BuRWC1XSQW4/ILooVdsY0V3dOtNhjjjnH/YwOfPbXTfmDdxEcsEu14xgUWim7ayVjDDh
DD8FG+KbgJxDrpeVRsbLt3EguwD4WHwedCJpQ14qYktJ+xAjnYuhTH+59dIzvDTeA+mSUUnJMCiQ
WQG5qSgGdRl20KfVABPY9Jf00qWgP+wScg07M0Z8PGvRnc82J1ZatEvkVBwzgFPZ2edzmOdxysU/
bKpHCEWw1+s6u7VDo6g718Gz32Jp0yf3TXB6L+ndszB98etmfGu/RiaaHqRvzpcC72ZSam4uaW0J
o/r/pcEE1mmHMbuCRcXzbseA6FHnmAnVn1V6pigOYN40tSSrV3fxHPFw7w4DFuuGgWGtxMD2BTkS
Bxs9gvORR0i4K4ePBtK0GDaRcEsynl2Dz8JlMHFgVbjr4wV5BhkPupqYB8b4QngM/XGwsFtr5Nm6
rn+r4INreiJvUSB31hPStWDPYnMf0/sE7qR07ZWWUpTqLHGvP8jTtZ0iY5KKXzQMK/D1a2zyttBn
CHF3TettEgapegt+RyzXWkH7HZAqaQgjpWfcbiGgUp2z4mzTIsshzKFPU0VSo56FRelz44bPAioz
/yO1UraQRL4OLXbYS9ux405Ab7ITALd32jB6X8jTPRDi6Ny1JAlpHEeevUFB+NaFYoA/hmczYW1H
hgtKsmhYizhzAZIj/cg376+CND1yP7ZTT4mfOzl2zHFjjLtnhIiXXYRzy3eey1OdTjGGgpjjOftc
HLQIfDmN6aROo5L9zRdez6JxNUwY+CojvOAeMKAoVqOutLXUI1lS2xwP2+FEqRCJYnCTJ8mqDJOp
Zj3ZIVWEWgbvZkKENGizcHT5Sx7HsPZntgLAtwSXwlPocvH2foHddt94ltY9czkJEqNlls2DzPdX
1iLsOFoik0P6ARpwxtGSn6SEEll3o07+fseWlMD6tg6HcHBCLhzBRvd6xNPx4p46rwKs/QO5bHQ7
xEC2JEZdgPiaf56ZwkV0cDeAUkO2zFkXTQAcMLGyJw97WoCPwe88orQiuNo2vF7oerdCBpKTPxJy
vf8ayXKYy2VcQHzenXk81UQAr51yj5edlAcHL9LI8fcK2cP9zfhJ+/MdTGd9wQmeX1Plqg2GXihk
95tQdnnb957GPsogm55XDvP27UsbaISD4f2WkmQ+dxiLNl6H1vI8AhOowzvdDSyIX2SLUisjPhvu
Kmf/Ic9OJ8giyHfCcELAAJ2SWvyyMLNDF+ey+ITQiVjhIklGWtFS5ojf7iWXNHwLWpX6AixzaLFh
ZDDLCTXgE2H5v3PUeLGDQi40YCx6cJFsOXSH2/tEMlpkqVXA6J+ltdsJI+yOzqnV3Q50kRTs2uS4
B47QdZmvI+0U/ZL7rfSQR351iosfzgBihQb/TClcIh6ird6GPUKQXb9CvVIu2JXWJUynqL92U9dG
lAU+2ohUCrj8DjbrGwhvUeYf86O9Tdb+zu+ztuttiULe78JGXAOBI2gXbcGW5+7iD3NsA0J3NrJI
7Ou9p6FJUbcZ6FIc4GB/qbyUQaRkqYMqTOC7BdwonBOZ32ZvHvPsSi+6YaquV900vFyLpsjj0tYg
V5biCnDJ71FTQnFWj+xhL54Hb6KThI6Z4JeF0QdhKRwu83LmFgSUs07Cz5dusDokPTYXvY2s0N3X
7vtFXzS/z8yArr7D21UHAgP67ZfvC0Iw/fUs5eqy/91Mh2Dmf2sywRLZeISiKwIXCFkl5Xzv8cHs
0FEyWKygzRteKLRMVp33uUaTWuPQeyq5FbonSMqaNGjMH2rMIhnGmxdrlij3/s4VNKYvIu2SC+V8
v6pxxWBWyAbvFs1mbzQ5R/ePDs+xDgl4n3iwqehW0sQU3L9YmHWBlnz0EWhS6Cgh3wA56XRm5yeJ
bhzEvFEGa01g7mFUZwVYJsRra7zXBGvpZOpCFXHw8NP+IzKlH+jgI0icWpLBurXLNoDO/7tC4cXM
yHAs0LWNUTMEkslCsI6HBOu0ZffQxelC15M0KXW/kNA0V8f2zr5dz5iUPNXkZuvziLUy/seDIPrT
q9rOt+ONjnQTy3y9gOZEcC+ZtEiOq+Q2EkGx4WZZdAz8dWWHBUVjeeJ+SwTEThY85YVGlURz1cig
Y1yuc4wMxXdHQoC5mXyg3/WkF8ND+GyoeNHatyr/qOjsZiBayOuFsnUHFlctrrJtdO99BxcG4DWI
LNQv2WG5J9LEKjzBT1hOVe4pc9FQHRrMBtcuze7ZssZi0kwp8XoZNuLeFeFDXhtw1niwfmcgAsVi
mq0E0qZxoPudr8dO98/0nBsdRmtm3NwN6Y6RxDFlG3ZihyiQiyYph6jdA+/bPhb07fnjVlsc3/eJ
HvwgOGruSd8fo4asme5jE7rfyRm21WnGNr+WxqvuZoNy4cXp8u8p/obLqJdpBoAFwJd1sti0CQZ2
+x2dY91o1topnR2ipLNlGL8njELR/h1LxhH7D8oplunqP2T8TqN5pxZCO752vpRCFJ44+fuJf9kE
BTYylkVMkyNrdiE3MJ4X6c3Ntm9Zn96F4p0tzK5BTk4rh63Sl5KqmEK3kB2UF7EHDiH6hpwId1xK
X9GKupUj9ZNetj1rFvidLbQ92qMx58oYjDYoJGZHkWWKL+jSzqrwe5X4C3dBXyfVGP234b7raIT0
6GV+/A4tPPOcRwU1HxbKwE53E4O9LVKe6gcSJRDjJGf+SxRoL3U993A8jHIp904fgfJ9P41UA1OT
7/DsPl3ad5jYdFm5MY1Jh0cmeSOh0VYNGxPnbSvxytd8Ny0/8HOWrKgdoipVBftVXGgQFND/w3Ly
3C4CE8KG2PRY2FnUnwRmUQrqPww5B4V4NRbNklR7Jf3v/WXWK9uuy9MULA/GwefnsnsaVssoAZgM
9vwpGOmPxGEhjVUeq3PGcZLDuqCUe9lE8kAX6YVGywfdLMTsQBSzWvjzQhaquzmcMS/xHLZKnRUb
l4aLpcthRHfi60wfygf3jbFi8I5QYkudfZPd16pq0n/Cdt+noYgfbmd+Sn8/Y/sso59ec8hVFZ+o
CbYHLtslFvwRZaeSYKAVQv19fOQem9KZJb3bX8UFZAhVKKTfwAnPowC2Q7zbyQaiMAf0nCbhjtI2
0LSFfC1sxicyCEEo4XZO+3N9iMp+SOM+4/7WLwcqJZYHcXPmUNfGiDMlfxyS83gBRqwHsojl5brh
YJGepIBmRC3Ju6NMj4wPA3RriNlfz9OPEa/EUzJkfwFEkO7Bcxw0lnjEqNvt69gJ5IyTKyHLsonJ
xXLgurEMADV5dcLnONsuFrJF8kdYj2RNK+Z0B/K2OI/d320F2gnbjSOEnbLOO+DW0zPonGN56dDl
CEIGHU7ujsv92rE2y6iSKLlJFNEBZRKSkyBzI44u5AOeHxQXj4GyRVdBNLzPeKAtqnGNSPa+xlgE
O1n2ZcN+4bzEUtmJdNFs2/evYv0ocM9+eqGcdyu3DBWA5QPH3ojI3XhiTv/HLtyHqEEllhtPzRUb
vIxYA7Od5iSSokQmPaNTDP/nUFJMEfB+KhXG5I2EfYW6QnYhA/DO/ErOGSHsuhsDynzerxAefKpU
XKXXAODjTcU03s/5Qu13hSrd3CxDdbWkeDqSm0Ifz7d3esm6Ga+5nLKwbX/kX0aDbtlFmZkEcTN3
FoG7jvGLmPOlLFBIVRYKMOGf1Pn5V+7zHPYh+BAbuw2xzQ3gsIgjG5u0N4+6U3Qcb2l9TFWwtXWh
t3zHbl9v3pmfewJa3KMCgTNJ28LSwgGwMk1q4+EJH+4fw6gxVQhMQGAPGadlOLTp6kVZMQromMER
Czg2UZfJnDPjs2IHx9nX82V0lXqO73BY0VyPjOi9q81UkjCt/AiC+zvtC23wZZ+Q/VH0QozFdv9n
mGB4bxE9J32uPfK72AS3eAuAtQc31fT1NT0Iny4AR5uZ88yIpdlO7mPLqG+Ab0l/X4Hh/mqzfuey
hCZSylTsq4xToDS8QR0593S8ZqxVE0CLXE0N+eCdUvHFIfT97Wq4mHnL5nFICJaAUwGHKSGBk7u/
m5CBjQzJKc+C4i9uLhG1pPOWMrqhZ8kdMWR3+e0h0iyx2pwiU+0BOlMWNL55CkvOEIakebzUMe4E
EAWx/HvLU9cTqtvWPEmXaKmPPHgxIAZNp/PH7jQ2Q1cRfiPX5OK/hynMIpVuDFXF4N30NFVY5NQV
gZVyDvYkTpaSmxYSK4XCo+GEBz0oFqyu0v+pwmmN8/dcPQo6r8OShAdub5RTTkF7StyPEuo/Bbq+
4XVmHtKmLz5YTKbk/NFMAYFWqhapbMEbTv7wIYoZ3Bm0HdwUDoi7Qy0pDPQI4JvktbJIOhjgtc3C
f3IHSpBpOPROcOa0v7Lz3BQrXNZLHNPvSAj+TbK3F4jZQhjioUfH86hgKftSdotvGorz2HY40y1k
QFJmXXPvIkg4yT0g4cnkVn1ckmk14O7MNyEV/shFXQHPBVvxbf+5O0bFh1yqfxvxDrcA2AWh3hMt
OIry6kg1xpb7RODd7u+NqbYdfvPnb4XtBZqGRx83de9ZW2wDic2Xe5zs2B1FWjhyHEKLpLLM93nf
LzklRULuTy2fExh+Hs0Wi28nxyvxXDBfib0+r8LBAmIzptRucGLRJMlfT0WXykPppdChTsE1tgy5
ssbg1hHOnIXR0CJmwUistBjIaHDFOX5AANJrKgr6BJ3QjpdyQ49hyBPU0TBNM2TxxO/SPFG1A6mM
xN2JGJPis080FilTa0grTjkVa9h5mKOCyo+QviVUg4pvX6CMDj2nq9vw41iLZ0y1wqET+HlxT/5M
krt0JCwsIYoJG3mVMpzitXBSd53So425bLoveGPYAXcySfkCiRAqZ7Tr/tHafdAaphY+BomHLmq+
DXWkoUbYVeN7+xphAr19HPwAdP8FGqZsjsDXs8SX6HRflfNgovJHZqSxMKoh65TWtS3nn4mnTKLu
vv0waTxByCcCUk+fISw/PPHvJQGaT/l5AG8EMgejrVxPi9EzF16lz/dvGbNnYCumeFv//CGKGozR
ycG+peo9LHplT7E3xuJf0u80nLyagULt6YWQHNk9WveCk+5irB3pmsuZ7WoTOSQ042BEjFFfOSGL
D/WeSvoImmg9jbt4ck7Kh1lDbg0vuVCC7ElEK5ZXq2NUu3rbVTDXZQFC8kXqpaLdSea7aoMwlJpY
miaUOqvbEj8mIQ/LVhiPEddk87MHsnBepSwDHduLIjN1vk5lem2LA2ijeZJQMFwF2eDcGUtCRcej
muAXypg8+Y6Q0cxxcnpRo8c8p+M86xFoCmNw5emVaMVia6jh/PBjsqwycWJfgyEljqvfezVqkp1l
s48Z8K9SSFTUfRBnvArtIuhhFGNRcIrLt79D5CPGD8Syc8kbfDOdJ3Rnvv2hAtqOPHbNojTfYdCK
kCTCz6AVlu/D9tgMhX40pY46/ISJcZImBd+jD8sT55qSzq+AizJ+PKaIKqEqtP0KNG6NAyUDQ7uC
nKqjQSfDoCFcxs7pqQR8LBi1ozJcza/CvWYhQ1FbH0mTHR0SRZJWWEe6hQe/6Lzqa3nXv3StTkNz
axpYK6Ck1fKLTfnK2zEU9KXjiUFy64eIuYOJ5Hr9PWOdQqyo32R8W+5lRhhs1KjGj2ScQsNuLG8i
RzTS4Md/DHLcTODMFMtl4AOGZDBRn09RSxohE9/Nae4ZNdYj86QqJmal+Txw1NKm2e+dGz45I9y+
zn9lX2R0vRCcs0ZIHx2jNm4m2WUXG7AXOMxCDO3GQ7jVuwVFJmHqCdn+FJoI+OHd9emymQWPb7MD
Bva4k0UWVc6rsLHStta0Q+V0vpFm2OpmV2qkAfNh82iVrhjCbiMZnzN6j7m/QOPNecmgUCVfHfX2
ogFVXW01dpbn9nXDpr6ibwnit9k15T2LkdoX7sxxj8X5NQvh2OFWt54yDwy/q+Jr4wHEHlukxt7i
RmX/APMne+FnF+kVJCEgQ521ZzdzFu7NHbL3qNdlmPh+9R88eFUaQjkttCSHW2PE1OLs0wcwKq/D
pGjsxzamV5zePoXUhbppv+k7cRVS+EWUW9ZZic57ep02D3LM/GAq1V2ZlpVA4wpvkCqWqXdkJ8V6
G3kJomzeskCkDvQ1PvzQxBiK34ZHClcGMy2ybLCdgUzXYxd9bbwkuNHe+UpOHBdEa4tpUK9UidZP
QbbyOkOXcR9L4ii3FDJETcWuSnM38Me8YMEbQ34j3pl2/Yw5Hsdc3axEfd9s/jq5DZCyIEoyZ65S
x1zDaT/Ni/hB2+54agphcOohvDRkdABk1uGIKzwxPc1IYOy3kTPA8iUVxK8zmN6ETxkXXxzovYrs
B0sFluz92wRymsXh2OfucYNSd5u0HhSdbmyr1CTdiYxk3YPlhlbd9LFsY2J3ix+IzlsSVDJiFu2d
eYau2k95l8xw0FNaGON7HPFpGO/6u2hxS84hulu99RCxyxcAYUCAofNfzHIZejNZgxVunliRJTtk
umdn6UxN3ALlFmaa81/IcJoz5AK2V7z++u93oxKO/ecKwFuZEztw+DNrsPcTvaUkdCtrDzbHiyV0
+7DPflfNiTVp+wSCvKhUbTJJgV8C533HXPFc5NolOKohRyCoTWaQBl40PqbMolanwJqKbMuUTz+R
+l9xLa0q3qSI1Tlt2xYOZe7aYivJWjJeh9UFv5fbFIzUC/hGZhdf8LnFddLbqT9VCW9NLYxMLi/e
Qge0ZaCdLIZxga+Ha3ImlRwAAFB0VNN6Fz8aATgAapmPfhzNwmHZ7nqEnuUAaFROjRhBkjesEm/+
1r29xsm1QdEjDdYEEu0AgW0VSq7H6rxWArwcVqKQ88YqK8k95BOtI59U5nwEkLn05dqUyyAnULKF
uGEqRHsAt1TRlE9CCNwnraMCI8r3iZ5V+mXY2QgeobnEAWefo9wJjhCo1PA4yhlLz2UxKMg5i6oh
0LlixM+ttxUiKPwXKrXx1yjQbROdTX1gowyN7fNkbIxo25rj6foUl2Qz5mie9fjYuA13sdmSdS5x
2w564Z200ONK7IF01LsKfwvYxvy6+LSGU90/dwspTEB2/8LHAcbhjzNjmY56H4yANgrKZTp21Hhr
7499ODoszpS5iclf9gsCyzR07mNKU+rX9qAcOhFFX8uJ+3C4ytYBwjhnK2LZqrtpd6snxint2Arr
sXIoYc0OBdoklXYIeKEBYmErOTL2Vv+k9z+xEPgPvOPy07oHuzIfllqhRtRiH8AWzHPn8PIe04l5
j0Cz8AJHHFfOjXA9RcSjJMfUWmCDpE0Okwgr1Py2Wh3I/5lEvecuhSiNeBndJW7OSorI8oai0I0x
PhYL1ZMYR6Asfegk/l8ibiXPlgFevjO3tJ3lHn0JmfKU97N3NV4vNxUwvoLaY2D0AE2Q5oQZve0z
11zJIC2xHV9qxV+zxNwi5RqhDD5GDUl9+UUCF48Z8juCF4G05+u+v9cqHA9b7BmE1D8b9QVroszK
S1B3+BZfYqyLOt88ESAc+3ql1c5ndttKjOYodmGFavRgRMNAm2Uj50t548C53UkFp6Sfk3I64AAl
xsppYNmSz2Kh/HFzteemE4HGl95IXeEa5+HmN9KwfVa7nnfB8iW33VxLE0G9jUIMmIYFT18acoue
cH3SqbEtrMOpl69+q/HsSde+zyfUz0lUC6TrZVIG+7PYThgQZ7bRK4c7BNVziZSWaoin8I2TbFgQ
av2JtmsYM2kXT5xvfe6s1yu2LOIlgl/XxL0uQIJP3QGLSlfYOKQ5X7Fl8tXDLyro62Lh1DTI42WA
JK6u4+eCwB1Whon6PmoaRBRDPR/lNLnlrfTduj6OE9QWCTYjZsmbi4aDvxwtt3lv5oKw6exuPTd3
PfBWuUPoGnpTWgZ2UoTy8oZV/7dOhguu2HELpf9RCKdILvi3OIfOSZZDTpEVcT8dL6C6SFiIhU94
vUCnC/QEmdXXke6nCYEL3ddBHMCAqFVtALpqF0zBNyx5wXjSJIeDBsnkPmq1g7Ltb6N77kK1+ZQk
wyKj2cp9a/0o0bAk8cvlhc7mbYmpM9g4PoKCRa37TbGJ8v8WCNb4GUitq/Fj73qHkZ3CWlILlYDv
ED8WYFPJofhf2DiuXA5NSbsMcqIDFv32x8H71zl22q3zB6y2j0PSTKS04vEO9XhSJBrK4nC8WjMf
7aoTWuQAjwezkCMP/1CpVqfbIe3F/sY340Ccg6RDhCG7IJk33MauY1dRDWIVIM69cnt1Pb3b7JkS
s5V7zT0Vh/tLzD2XT06gjGJjapvniocDCf0vDaghEf3IyYdlPkMdx3R6O/rVGoe0LDGnSh1RtjQ0
ZgAH+a0DCbqmb0UVSY65a1k2mud6gbepIlol5EOxg1U7WlYnLrhk52u5VYrkX3uIVGgj8wCQG+ow
XnSTnLXpjArpKLJELe/K9zKDyOsYzno93kzs832dq5x2PIfEuWZUlpgG4Kzm3xW81xlpbq6DTfFt
H2BnUYjXXElJ50G1x6GFg37Su6ge/Hi+aJPlg+MBU2qkpFPx5OLO2WKYvOfmL3a4l/TGg6/E4BYR
brMrRFV8bt9aODWM2BynQb3oRKBZ8NZQCYSTk8zaBQK1d9aX0qa4c9ve266LssI+Biwg2FX+OjFD
w3DQUTdkUbJbvVUeSt9kWK+/L/KTM+zp4KiKVSsUVrVyrF4no0pDpQ6WPNkcm6LiJ4onmurnTVP1
yrkJjdOKx1BxHHxgMLS7sO6dt9DN6M1qJe6wcw2yMquWLHTVv5VLFul0Xxw/HrbhizprtlipDzKk
pZLNwnRmXu6vlKet3/QEk7dABuuxJnoZVerPBqMq0CC6ZMGNJslP6QNLGL6pE8dXexOt/N/thMB2
eJbZO97bxIYgBUshCJC7MfBF9IErR0iupaTQzilGtjjMC+M2Pp1Zm/lVqEHafxZT4qJMObiQ8IT9
0xT/1zYmPWUzvWOr1SaqbiUNBv8ylOe8I40YYm4Qc2oSG4SwiQbgMPF/fOSEIQzKtf8EU847AT8C
8AQoQ+CnxPtZtyTfrvB77afE1f24fpAd4b4njMsXv33IvECy0Ti3ZcmZN3HziGAd7ZTXwkO1mXu2
XxBgxsl3TqS/+OuNbmtl0pqiRl7CXVmQnnKzSsCnMhUmUiCFbb8gfdPygdVpxCabg4HGIzxtJc1N
u5VZMg29i2IIX+89d9Yk7cB5GQ4S42sUv/0LgcJVB2p8rNr1guPsf/0QWmP01lDpU4P95bFueq2J
nYKQi0bFu3DKRFg8Um33M5PwvgCWi0YjM0egWp7nsB5iLF5kXRMTukaG9cWeX4ctm9nUGYpE7UDk
wjpJYPPURMOoq2O41C7MEIlLtKDH1oM1H3Ol4PsrhSBOVIjqbeP4T5pdBPKTCQJIZ/Nw3ujs4M/+
9QZRZVaD0DR7my0x6oXDwKOHEhJhqTqvg8Zt0+KmpGE1stilmrNBkbDkzjRlSB+nwi/h+SViHEcT
OFEx0gz48vxQCP/J8uq9HNTaFq0Fm/wReChz/Nk2bRuDSj0U3E+QjaJLIgLVcblNFb/1PF/sNlQs
hOR9opE69J452+psApVdYPRU3WVXMTKcQh1M1hL82sb/QVI7expFEOqr1YpcGaQ0YA6l95EwilpA
5DFCORldjVWZ769FctFFaYLigbE/3ZHRFbSIKpgh2XFR2qyLk82eqbrZ9XkJqe0dwxQaBscQfgu1
nSVfxgIHH6qTccOa0Dd6+oJyQ4qhvIBNavkU0M0SVR774D9hWQ/oCoo8o3xgrQAYt9Xmy5SBS8hq
aCzpCpAclUmVEAvKuwHakpFtCPGSO1B9pbHUt5aOC9sjI+MqkrJZ6CrO6IS9bCThkCC0PZC1w6Zz
h5VQBO/7VtkB9EvqI/xBCSrt8X99u2ZcWNFsmYu1XVUnZQ1N3NoUD7NnJVNczFdqjkX/yR4PPEH0
J3Yg59zCVpr8Gxcq7rMD/TR/YyHRFUWYnp8c1vQqwUDpMESUI413QQH6msyJR8vGFZ/y0rqqFNcW
+KrZgjsTuxk2IK3527UsMZGZ7qp0w5Q/3h7lFZL4Mct+/J22LBENN1/m7VdQauw77oscVFons2zC
4OdHUWVii0yoUWiZzx1xVXfbtFbLF/g+TcthgrQRqNrQbc0h3w9KeN+q29bIZLsfHrOHzxSYwoFb
75LpUt+mn9iVWj40LU67PcspLRrowMEaAwQUF1v5zQLL5Kt88gVOUe5j6LvAfPXfaOSMk0MsByYH
HTkPPNjkHP7kzZ0FwJUPSKym//LELmOYmPwTk6SQCn0Q+2OLTapQujMyN1ec9lDHBoF87TOStWTH
jq/mfQiVoATNoyZR4M3Uv3LyxwFctwtfy2OmFsVvsLovo+oEBBh3Bphygy08EDRRWglvBLqwbCgI
MeTZZ8OQunkoLVbu03hnucPPrEA3a/bF8s86y9tQ6tePytaD2qN1gqxURRr4QgVvWG4KZE5HWArV
A7D3EuZQrmkgtjvot8a3uB+VwJfNfWEZGSjRgq7Q0bVQBRR7kG79ohPhLzrUSidCuJSmbC4OqiSC
qPThTsQNmNjlSFBLDDz0Yccr5AKwIyKhiwiE38eCEg0Uts3rZV6UXCQpV1ANaYmzFl7ZcqANwY3J
KT78PBE2EEcieDkwfXT7ZKzaH1041xxSQ3572IXb0Gaw71JL4zZC3yC48wc2tGteNOjXh1aNaSY+
09MbsbouMwBNU/u8GhifugPVwzvyP8kh5zqlmie1yD4K34TGeeeqKdER2jAyiu1kCzvZ7Xo1S4fx
6JgLu3MY3LovuZBIu9LRTlETl9EshKbi4PcDtS3d8ogU/uFGb9rdHjwk0pnFKIvdTZSRRbS3+HNu
x5FFmEZUjA84/QBIW1/WDcotf8CQe0gFzMJvrZfPtFyW7VvAJndG4udC5YFZCZoTTGJrPbC9Kns4
VzthwNJlt7eAAn12Iz+bqo4esd6cqRYAUsawtfewO8PwpnOIJlpsEMqZvE5j5N3xszjlpKmzj8SV
gd4hINFdBEHApTrnEmHaRC/Asb0bbm4/mbKXYsfYu7em1s4xD1pDZuQYi/JBR7gQ6Q9LOsklwV42
9b+BNpmumbrUeu6oY6Vjt37JrMOxZCIsymjR/n2l7Lep6SS2oDWsSXkvJRPOIgLVTsULk0ZKS1el
JtY93C6/Gclbq3TZjkorjbJA9q1JNpj3XUudzNm9wM+iSn/APX+VJAf+pIHGV5rBOnFY2cZdO+CD
pnJQYtblDuu08KbigvnGYQM0LFRpPJKCe5pyqkjNJDgKPUjyx0V6hp6UVBtyqroKf03l/PJZberg
OYAvaiTy6J3vxhaPJ2e93UNWDXh5RJUXD2zIuMH1GmMpjT7H/Xr8/TTCgeF4j7g6QMz5ZAMkLjpy
DqjPirzP9D7BkFa7Z9xFVP2w9ta2Z9lYtN2ZM3EmqOHcAmYu34foQbIoDodR56No0ulRMfSdfcmG
YUb1oKpwVa/Op+OLTZHh5SH5wKueLLS/Fu2sh32tbWfnDAtVP0Di960q0BqGnNeOhvZjkScorwIk
ipBVPMUTlq2FnQ2Tk+/300i7nrtYDyF6YAq6SG5SQttBuFT6+3/bNwcd4eyNn5BK2KKf4SPe/z7d
beOfFGzELbGZ3bI2HeUQdO+RDg50VjJKnvZISW747bNNN4z2lWU5sh222gIfGc+TM3EN9JxB7Npb
axamNYxahzzcO/7vd+wUkHWiXjVTY6DuekI60f1vnHXwsCVZpM1a7tTTbB6Kku1TckHBNQ0TdLoj
wt3KbJ6kNU9yN+2ZQXKrqTM7z+RSGB4eSTRKh08vh39vmn62JxZQJZYX3xqUfWrNVIh9A8TjG9gW
IhxYWFm+9B5JylEbZgmWTeApvVHJB6aG//utJFhhcxESc3pnjTbH1j0r6K1/Ka0Eb5kpeUIP7FG8
4LO1qPK6idPruSjddQaUaoN/xhZGT8PVokkcDKfPq+1vMic2oTTQXkOmMpOQMg8eNoHriMsPmd4H
n65IqiAM9YDzA+KKcn6Irfu4AZCOkLdpeLCxGc+si5hi9XnjtLK/ezi+4AGvG4RHfNgLP8z2od7+
DuPrsbWKryCb3TXlMfmxGfA+rf+DxUHqow8O+WjlJEQGQCEC+9ktgeVH8foUBHv2sN/iem4w66Kj
Zm3gm7NuOTaS32gzsCFA7E61T0502Pu8fDMlkpRnxdytaGIrUfxURkc9eJ28XYPgu9ra3pECXzZJ
vQcS9G8PipceUNm9AwDkzvDLuSaSJ6OBAjf192zB+7o6uwpMjyX0Uh4nRvethMApWLONAjE0u/G2
t/kno7Kh4MwmFYE3dV9PTvfT1wMmS8iryOcYnWmTK1ggNAN10zfIDdXhMLFtpStaqGtSrtsrvJk3
pYG49+rL7cQV3+RthuIWaaFV2hoNfBNsJhRfIwoeY9zaBtxXWDWvD3Pr8zE2NbSQKcwCCWXL4Zsr
QgfYlUrr4UHkIqaydbbg6lKC53n73LrF7HwCmSaD6MVdQqwkb2Bn31FcIRNB22T1ifP5l3znWlzK
6zpXJJELbdnFLMXrQrFXsgCd18FyylKJ7ZVXwTSfvbddfB4Azd/DdvQU3uDek25UHAP/m6Fqd2dY
DJlHaqzUpWvRmU/Q3PVXLvCjj1+VoLDl/nIUModYhP44AwVSGS2awR04noWhfwOGZeElPREIk2MV
k4fr9I8UdJFd2Rf0MK+TJK+Uix74xyVxnoLrscROqerdEVHLJ5EfrZoWjAN5clw1cchCIObiKUKr
KrSmfmXxiq6sM+OnVuxlqPs/XAZBgcVJn7HH3Vzkwn2q5Uj6096hzqmdn9A4ONfIv58oZNy7qJK1
CLR0HRFo/31YMUjDtfjdBsOmkZoZVY+HOugM2snIO5cYG7wOk5rrvQu/FoetUTafr19mrYL8iBz7
Taaso1zex3fuHnekK50Y9wvKA5GwvFBn41sCZPBDuFfxdhjisP1quCuREm+mTvDqdS7kjHDQ1wGZ
MZ8ht3x7tWrl4sZrBywA0Xh3Ab+YRh3af3MsGf8efOi0S3Iy+7BIFL6ub+T8dQEI0SdUQNnbIL66
aFmtJZoilUvJg2ONFKOhUV0qf51SLHe/uO+Fa+bj/tLxKq61UJ4GgWVoNAa50Q6i0GAnegeyz7nm
PCqTGngj/nGUrJLhFMOqMo06wLWwhIXymalnnl/lsslyJchrwpNq+bMMoE4pPoQnn8qEBDJpYbrO
X3p5Ne28GYkIn3Se/0572J3o+clLYdxCgaR4beeCPQkiQxnqvUlc7JCnsRgVJJN85SoVrq3LbzML
0he6gIm6Hqa+Q0BiMl18nhAqhjm268epINcTBI5yDC6fps1DWlgfkqx33dmOy2s2u5hx24LjR0aA
hdNh3XP6xlTlLHoSMSUKcphDIEHUEN02m61jkVSraU3W3rU/3CXE48FzMH2UupthC92QELkSymMP
WqhdMk/J5Cs4ScUeqazvq4dQ6raPYmLe+CsXROfWiuInzYHILs6zQFUzZH4v7xi40h0+B7O19f5X
cb+CPa66d6Lha9QjjU3DeOqYKDHgt4/nmz+8xEsSAJIPMSWQRQmrmV3SkpDHSp2lQwI6q0rLOLxg
aTrW3TA8PcrvtYsQKLI/QWNWMZ7mUZjvskbkYJBUF5kxhFjZcZAlNkjqRuBLRQo+Maz6kaWPU5h8
t/X0ZDfemlzlhrwjlj1DEhuV3YQicBLdFSK7hPiSF2BydrxsOpjDuFFHybWcpUIgQGZm8jeSXDlE
5609SaqXmmSxPkrw2axjdQBMq3LBzbolD5useuoTCigmEe+wHq1FqJC7uJSc10nXgcYXXxdJtmML
dz571h7S4zSde5YLcL2U3yeGgaACnt7yoc1QHjd5ZsJNfVzAPstmJzDYNJ/fyscVD20PmVaaqDRX
sCw4dDuw/HviY/fkygwFxHbynuPChMuPkrD5vePibPWTf/vSBgfeKfqeibwZMfSXcHRyMd8nYyCl
ZjDCqD6MMr1qh2LYARXx+zusx0FBXskELR4m9HU0WyQNjdiJh0TGJPO7Fkw4vya7d0Uk7YOB7XDc
K0Lma5l2T7eNxTEW5a4JL28o+8GlXRXy7vclHv14YaTpxNNkwk5d4qQob3mOQr/FkFWMsuxLLsJq
qq4CVSSVS7WZXfqFp9a64GS2BmMp6ANcE/QKBoaIVpeN0Bx2JuttPh/CGego9FrOobik8/G/G5qm
3MV7azhQZePOJYm4CaZdutFhYi2mg/Vr8AAodKTJLEgyzszbNI7wMI2CrTYoQcenubmSi2DtBZ6B
vqSWbtkNXvwnnwDZM8jARSiL4PsLf4GJ+qY3VZQ5VbxvVNhw+ddSFL7zCwRTsqtOBSA36HgtHZph
3hf2Yg8WqgikF9JzrBN+d/iFlwTOTZDxZziDLAFCCBdw+YVEzP7iLDPABU1vcdWoHV02cnCQvHzw
qEskP2ltaM/MkQmj0ERmJz+ui5SYoe9OPgu0cRMe5lOhePtdJ3pI5e75p3to+ciVaOBEGkIJWATN
vFHXllwc9EOUNrDW43Be5GZ7b1dkXuQmsOyn2xPupc8gD048E6VSNmTlXhiNI0HEBpj4G2j1TWMh
Yx/YSTJKmUOzcOXN+MY7zxwlItnOzwUec0yF8rcNsb16Gfd0nCdBzf1RH0euMFBrFa319QdQWOhQ
NWP9ow6Q7eluNiD+a6ZCRcacnrabmXCawAtU4d1qU59MI0IHz+6YOgSH+vEVve5fhtRyTusenvf3
5TWS1hJg+KJxPmIXg6Nv2QA7fxvjjFwPRRrO4qtpkOD7DDoVIDDQ6TiQ4rjGO7o3ot9gz45QetKQ
jUnh3iYOu/zU8zNBlqCOtan2owm5BtJOfm+ar9rxRifqFo7JcEdip1RkMV/ku63zSBVttRY4B3T+
jQD4vtzKYhEJwLR8c6sUbP3cvyRmpZOSGmjISkM4CUpGPztjzk2XglWQPxpYt1Q9th0CHXtOfRoO
oxl7aVjt8sGLi/S5j/r+4AS1JoKkO9uXJ8C89GGssJS/XkVKqTXc1EXlow/3BxwE4dgMZ5oFEKdQ
w4VP4B94MshJSKZkBN0+rF14voVIgSxYeV3P7HVVXK99hpBYJ8YAPY3oz8hnvuh3GoYmrI3v5zTS
XabIEvHl7FES0ouu1vHJK1EmbraqgwwC0OdrQ+vMUT7uoZpvHIeYQ7I4Ux/Fq5oXIK3kdUtP74u4
vBC5AKkm8qVTtoh4nIyhQFN+1Nb+8Ha1XJlGaORH3aFiY/jQnSGvQYUKiNi57EWM7UnzxphpZoP2
519X55FjlzvykBd03nNqjpL93R45eeG1gKpkl8qp60VMDwO6FMsqWy2L1POxUSwY2nAcwiPSBSm3
mwG14DcnuDJVbmz0KM9o7UH2hEXecOSz5Jj7dWsXioYyTpd1L7wyREz3ZfnTDEbFwUrqPyKVNfmr
rd9nghTNLIkWT6f1vAr7UNIhVEmx+OzswOxMQtydINQFezoA25D/cxruR3hAtUC7mel+ZkB/Uid6
SZmAIhewDrWjKj/dU0fXHjRsQfO3Y++EkHUPpWR5MPtJDuoloIt8A3fKc9E0oSgFOl5qnJzu0ru2
p9+Jj+fYqHXPeh8DBEoMwJbguxyzMrcqbt2xrXTRuOR5H+IXjW0lBj1vIYXJrWaVc3ma75KfmhRW
Jo5OHvryd4IVWw+pgtcv/8l6DBaljlrcLQqAp+qnPAhvs4bEcAq0Tzr3pfOJYf+YbHdjm+8ZAkia
tREY8yAuMpCI6iraOhABIucQDeylCat34uoPQM6IGQJUVIAcZD8jnZ/zUzq4caNH8qpfp+RThdBh
EQA3WGO5SynK4YZEJPFc3p/Dwy8aJEDCdd5TiRxcQSVaMWx+2LjGKkAMms7y7Tp+Mm2ZCZ0TiqWl
r++MnCaisbkDDgP+9XmqoFWRtpqUsHz5ad8BWow0ZWBrB2e3FH8JQI0EXCo8XJJ9tCp5aGOP/o20
QtNqzQKWcgsa7GCxvE4zl0pk3/YL+tdsnzsAvRlYjJF3SVys2P9LWpAofPsE1cmXlszzavsv+Zcy
WRQudbG63r3c/uv34KXErJwpTXZjeGyv5oqTpxoDDhKroMG5krTPQZiJnyCP68kALkEQjTCgJPd4
Wco6sfet1se0EvtpUQYEIHmyqMv54sN5T0tTeVPUlr68fCxdvVZ+TYr2I73245wsKBwitcbEiDSt
9qbZ5HX7nAA56TNiGHnIVpyQXolcjByPfTxYoqo85xJALWOc8DZObmILbkGCkdMxzUNzeDuMUY7B
ugM4qMGTQ99hfny2L+N+Hfn59bWPKm6ZKpnEayqrSzIlYkcinFUJYL9MDwUmJ2Eb+YJIqpoRRrEd
DM9zQgfq3i2EuTSPY71deMRnuFpH35WKu5shBCt7LbH+J9c92v9W/+7d7uDDHwcCcVN6auAb3jP7
qvAgg42G4h+0Vv36vafPRmJhK6zEHTA4PEtRrtiFY+evCmuSzWhJFdoE+vF+AQQI803a5tdR9dCI
u5yU7bOclJPtAVDVpHr8ZJuithmeez/If8RvlzaS+axq9S7HCL7beGVLRt41H+D8zRfsaezJYVGQ
WYxNAaxfPRZU2xnISor3jsCvrRDxFeuy53qTjWhYKtskVzoYVD8mGD/+pqOyUJvYhk67c1ISU+KT
mLHDZ8hAB5YjReoKc9BnY+aSpfyhB92rM8LD18wKMzz1wVz738YvVoAmx2i3rEGnJfi3u1Casgxw
VaciLVRZdbxg3vL3GX49F3xywNtLSVy+255lP1qqGuENnI8Cg29eqW3owtChMXAd3qg9CFMMRI/1
fKPye4G8ZEQy7qP8S231xMWhIOgUWyn5tsOq8hX+eeeKinL3K6HwrnCS7ZK1hswaO6TqxRJEyqqM
tUBvgbvGp8jIacgZ/VcJCixqaYJm6sFVUjyHnANmtK0Q8Zn1emGg1wW0b8huE61EpJF1Nm3NTdKU
D/yMkD37iC5bZw6S29B/yvw4eUDbawSOEyyAv179r75uMf7lxi4H6b7O2Dp+7qL/WUqf06kpRgaO
dwwJz9cZwx52+WnX775faPcmu+sCZpRaUIizqoAjQzip7py7jyGsjXWvs5aGY/MWfbHLAcNL06mp
RzGjC4puimYHOPHbVzpmwj52S+P26FuA74rq4cZsa8koYdrVMp05XFFSUeuJsdSJ6fwvJRUwPpA3
HBgvYz+IsjSOv+3azgpQyx7ymJ8aw3AyodGA6EqKNmaIHVqk6cK5a4d2c1Dqa9Hy09tcyLDThJzr
JEe3ccfM0ExP1jPsl9WuME+wFvgC3ifjeHMwLI0rrsaD7AyTjSPPiGf+8w9UZf37jTcKWehrsA9U
K1wSjJXZ7L6oa+EQO0NIFYM56Guv8uI8xRUznJtJCUwiwRhA+z/2M37wEOCOserzruHnCG/2wcqf
T3+g+QcLLWjTcGxPVNi8G8PqiA4xRzLMND82vivxA6Ch6fHQqGwMu1oqcEnsB0VJSbUjh6ZO4xPw
g5CGZ3OujE11OqNhnX9pDa6xoBbI4c1qknoqGAp88TBMU85Wnf3eSaDSsuwtC+uoZOkjYuBPpkMk
YC4U/bsx7ShWTA82nUSFnN3roPU+rpx6eHWNHMmKRO3yhoedflg4HkM92JnXF0yDnCoMQw3k+xmz
UuP/0rshBmyEbJlO5+nqaVKoMnSXmShmCYB94h2cOc2Wri3Ba3yAYLoaWrUP1CokXe3s10OJEHdo
luOcZBj3pypVbgnm4Q34+HQBt4QicUrrDob7xjew+Jv3iDQSbp441IxFwnJ6M0KkY9IFp8crKBWG
vySLYv73rqnrLLqW8hTO0RU+LH1XIiHkO0PdGOAMB2gZ+KjbEtxAGgy0Z+ZimLkGcEHDGcD0MHhe
HKG4VD6ZIPwVyz2uHxqmL6I284+51IFU8VVIqABq5KvkDtTcsd2KLyDQJkofD5yOChKfzRBBUwd2
KHRdRyNa0uydzzaHhPV1IOwxaPWT9u7neyGEo4HXMluiFTe10VGrQm0XwIc+gFWeEO1seRKQ5GVy
zTN1h3nVgrnvGOpENfBJfoBbzlGN79ClUTVqcb8JTTUty2xjcUu53AVCKAB/3IOoKb993TEH3leF
dJ7WI/QslCYIem7qe8HlkvKk/SMqCFSO3grWC2AqVv39lz+fD3353B3WZUHdV52XEIVbacDAxDaJ
0rHzLnTpdM6UCxdwXzjsSd78fiJIhDHnKN8qk2WsS1OC9JS1Q4UC6wOKGEw7uz8TpegppET0wtTC
3NXCGdPFtrx8lXKnCYonkvkEe9PYYUIbYKzUKA5TCqcaKElwD3pYF0R7mLX/HFp0qDZpv27swoAH
7ZsT6UZlLzdzeqkvoFV3mnIeg12MNk4MffnqF7lVjKncVfhsIzTrSMkvj79hUOjrlYmy4d9d2ZZe
r5o5wEf5sOBuSAT/kxrY3LZf+5fiiJz+sWaL+j+47kdUrzSe+VnOfuRAr6vgxOYuqH50ZbzaQt4d
cAIcC8p6yy4Vgbi/Alo/t0WncQlUwbjj/OR5q9CDfL8lNyBzXg+bfFH4U9ZKYqNHiAEDT0iOuYUk
Nfqy8KIrCwtKA9Ptxfy6lGOYoAL5Y5rQQM4AlMItnK639LBsL3nH8rFINXJRFAKMOzRj08SEThlU
KO05gJk7XGEA2JqH6jlBCl6lpJjK+mWsF1ne5kxoboWef+9tW+n/jN1N0kQYBmUKgIEKlfQ/t9Z3
xwA5rvNG/NZoL+Jq2P/2KtNlF59QDeC1unMJnfn74wnA8dMOLRrQLUWVbYdlvT/DNy6b6adeHbNe
ApFz3jV09q4XtogNv+MYXiPUJ3U5skPE9bZCWtx1Apd5PMATTA8eicvglJJLF4oDSjTwW/d/ZpXR
5Geqp6vu/FlKWc9DYUiIFxz8wTR01a1OAmoGznQoj7Yf41iW9DJzxv2ntA8JvOHnQ1jlYeLQ0m20
P8FgKxdNlkm2CVPa6wcA4gpxHj/VBTp5SN2M+2HK8Xmthxm/RsUwgvUpt3Ngns9fsv9o2zHg972z
HmpX/5QDKI5+yc6eF3ZybT+YTZW7p14XCj52H830+GeDoUVZ/TOWo+8UAmdD47c2mk9XeUZRCccm
r53YB30d4OKK/3vmqqiMoW/TJrHKDuHf7IvI8Osy6cNu5P6RxsKcLKzapVDVqPEgY+QMWnYfXraH
AhPuEFFSJT6y4l4OQCEBFOMdq6LftwkjwFrZzaYsn+zOZl0HyPIo/noQ3pQ3/FdIfiUn5e66ftX+
IUs2HrimbPBK4XZN9iVdncCCL2q6/uXnMlO/LTl4i6TCv1ue4VXAgPBFCAGVSqMM80UHYLxJGKX+
bSszMrE3aF035dX7YUE7+LGu989zsCr81Y5fMoiOKY7/CN7GqTA6YEAB8cZrieaM37aWjKZu6aHs
IwHI282F5RNx2ZcMMt9+MOrDGw88hzQ8kR9cUVJ2m9mIGEOTXqWGDmFxSqeWHQIkn+Z4C/QU8q3g
xrQ9q331joV8xT7CvBSxiPJik/wIVY4b/eaSa7IUn+pYfHZX5wc5FIKd99TCWgBN8zGec9VViUoI
hteIoBDbNNM2ANRAUvHH/Q2TqXedZsBPbysGL2E55HyLDDoKj8524ifCOB+UW+flXEq5nFHgsHDA
5zmmkLf+TbTOXHilfx48W6dA9jhfyDRPyCD8dSIE1mauKuxHp8Mf4jNdRT24lsMQepDKAEPyM6oI
Cd8qXSAxf0l1sjwCYwQyGnJuxx++GjPbMWZDHZQhu/xhK3FVNqClLdr9XlkFu+XyTzgoWGWhMTkO
0g8V6ukV9H6dCa3SeFr2uRzgGXshStDvs14CcrmmDdo+GML92G4k+HCBqzQn409gvoifhEEQOeOk
fFEhO/tSDrzJEUDUB3nlSJIg5tARNmn5xQH95wSxtPBU97meeUZ+gdsemjTMI17uc6rbcOyvKHdO
iRoBNUz3/GWEfv9/Zv/59BjpP57XS8mMBGZZTwCfyJg1PD6tmMMfCGw7hjo/1tC7LdOhgXdRV9ZU
Z1IW4Zc1RGdfRq4ZUoqyAevdJKaK3WEsLaMcwSkrPj3JVaxxwd7ggtDuhbIklD6xWm0ALvH+jecd
NYm95AGIOxQ5IAUaP5pf0bb5cLHIYmBDyYugz1t9NwaUASnNAnwstVwUlx7nNyQo00moP+YJ7M80
w0eiBHojaJWs+fczpZbH2hQ23ZKJv/CzbfuhM93SoUV3dRzHoygyBQwvosCRkNdwcGU9hdClfBl1
+sSOiNk9xR/dGU39wC1eIxW96WH296CLJFmJqd/DGs4f07/wSf9VxMLoJrCGNhZlxdA+QCP/W/TH
X2PkuuUih4AI5A5VDX3L/lUrw+fXqmgxrDaV2R90FuD3gUKX6isV6a+PJpM0iek7pHZ28rnto87m
nQcEML2/cfvD5UthFrBlYk1EsAj9V6aBSfHNAA0zgyu+GBGqsXmkc0pX1ofnv1XHd1d/lk9iEQmP
AD2V0mdw2e91Zq3c8dvFpGk9uqWgX0+c1RxGULp65W2QorZKEHsE+EureDW8DE2DMNVEl7/cOp+y
dtndzx9u/uxZxcVAVJQXF/w6ZNCL0WzeCqm5TOrpnuDVbwOiVDhidaZRk+d0kQw1JY4AwBgUuaPl
vPM+lWrt1Sw3nZcSjxtJG/oA95kOLBKcHoDfiPmQ4s11mSN3tQL7YiG2lEBdfrhp/PFo9FC20ow7
0ZXSztzBwOrjP/TqMAAsi42UTz6nxeGyv0kjGCJ3D+3eTBONC34+1Jh9ku0rT9/afimDmv0g5aRX
yNiURlo/NF1PIFRlvwqY/dLUSQzU7atodi9EqEXSK/UKBbCHrTUU+EH5mJbQz+NMHx/+n85bA5ob
F/6yTWZwUhPWKgvJC7aDePczAPJTUCmHVjjoa9aLPdIoRPcxTwoj57yD7OoM9q3SqIMY+srL+04T
m114J/xFs5fk5e3QVuvSysjolQpX71ewdE6Vx2OiEEBHYUkUrYQ2d+QcIJtU1ReoDL2jFAKeb8It
OLYCIVyXo4WscHVYFNVGzBOp2sze6th414F5c74Y9zde+GAixcDoGBt35hADyvA0fu/sYBO4+TEi
cfvfxYBpUg69QRjw0dCEIjdagh9dgxiak2qzMBBcM8P94wxrKLCCT4hpBBrhKfMo1Vx+ePj3oGiN
zU8+2x5mYYqOzxPSSbFC950N4mzLi8ukfCyMSnVwZIQ8nD126+gOHRBYE+ol4ALXqvLB7fi/s6Fh
v08rz3PFBMBR8jvah94NF0wb5sYdrMp4PrXjyDyRHEXEZame785CGt467EVmW0nZ+w5bKwVeuGq0
Jljamg1KZR87fUiYn02+CgOxDoB77zGrRXX1plhi13XU47JC2dXrj/XjVG5xOFERlt2QcHJm1WZb
jdeEEZjz50/43/TexAxFWV/ngdowPIRvCm5+VNaSJlp/5TjaDZykxeZABpbIWUXbajdiMndM9ntU
NWvKzohJGGlzptcyO+L1y/GbCatsKPw789pGtEqOJAjAxboo6haLktslYiz8fMoJik8Y+TqsGvt1
ZEvdp/PvheaO+DfcOES1a4L7SGZXx17gR2C270FCr6t3HIzaXdE8Uw3SfuWDx8nKuEntQgxRU5r6
u/yBRKbLlSWfEVnxd3DyoMyZgK2QFcsH5QcTHP1Xha1uHiiigBU5PbkeNGKYvm26Y7u67H9AN4+f
MP27jGuR9mHitXAphFhjv6Hep+zbxgVrP7bmNrHDBV/Qm6JTz45yqWrKgGmlswzks2DrZ1LG6pBl
VNa/kRC4K1vWZ2nMp1iVVkbsYotOqoz+VuMFrSzBk7CNEVvaVzkyWz1rCC3tpr4eydlH9qDIAQiq
HzKQI7k6FExR7GuLa0nB5u1bD6wupZJ1Rspk+WNBd8/NINWVJoC5b3vJBb8Phpl39+ny7BUrGV7G
ak/C7oYRtCU16RPihFHlfV76defhESsu86GbvrHOCQLYJl5aYlpygc2GilDz7QWaKkUbNzJvWiSh
uaz3nLuCfQbWikbFYXGfC+iOAD7BOksoMIiSfASnav7qiW0SMxYzJqznG9VmiJGhPb4h2G1AtwwZ
4k8Sumjs0NZP4nAXUS44oRWm3X/vg0ygmwpaAx21xbA01UDSiSQT26oStgyUGSngFb1NoyZb5GH6
rbE6aKnqy/AjhFMR1bNixFnc7QND1YcQ555iVqyXrlH05kZeuz7LDkGLXINlzbYTX9L5Msfl2cV3
aMmPXIgocrE4YythvhZTUQWIgswS4JFkpzoP38Tq6atTqzvVDx5m6ghTuJY4KDyDCQF9oxTmAH9l
tA0bHnAnOw8rFSXq8BSLGrZQwqe7oX2AMeqV0TsPjXbdahxkjMHYnRLDuQA9US8Xp81p60i3BVRa
DFKMzmbRuJ/oCYvfCUqXqUeT3jm0Bp8gkXlBUo3uDo0q8XHiyNe6/a0hmrrj5IdXwCmsQhhjFvS7
Yr5UVqhZdk/tpT5EvCqnOvbsEltZuptgXDpihdI8uuCOjoNBX8O7RKZja0BWN/Rk/OFUwmZvRZ2H
jIAarosXSv+MlN6UiT6QeMLE2qjbtstdUGdRMc5kH1LmioAP2wM1/+fC+/cXJ9b5P2onbzJCKkWZ
BP+PMj6w+xh2rST1tZlBLZYKIHj8b5U0OzG7WZ4plFg8GJuSfBJaQhs0n3YD5nstwMX0009dksjd
ESeimLLpTZLcKhYFhYcEq0ehxlHxJXj6FrLjlprkPmIu0jGs1Et1GYlj5UzGs8uDZzghxvLP1hKD
IOq3FSpMhjO7Wg+MSNc22WOk8rQY+sm4OGJ3XH3wWa6FNlaoMGjIJVWYOpiOdSLMcn7CsBPfod/2
+Tm81cKKdLp1Pzl/3eGESuVsWNODZg1HyLCsgtICo65wl75fpNm6l0K3Kq3q5oWglKG3/r1hfMLe
vt7epYpEBebjyESIRLm+4ddQFNs7+xbhIUxdUKKRNHV7IT7tLjM/3pF6V2KVrmNlNv+uRn3HXonL
zyeOExVMJZOzYA23Q0L7uWKZ1by4hFdJl6LMrhT59DVjM72mMVOlLA2Ack2OWVR5t4bz5E5Wzjee
NKnf0i4DTK7kR+6L+465Fgte5EYyfSzHcb2qOhInt2N8Y34PkfiuOeLtFTCmwDiISlDkFCBHDRAq
aR/8kkxzmVbv+ecLFm46ADri3NwDLSO4jfwBSycgCwQndBvwEbr5YMjQDr4O1sh5mc0bwniPan6D
34iGR1zGwKlIYP389VC2ZfwFhYz2K1hufrsL3xxePOOq6X5hJU1XrSDFFtRf7YUFyQYa574Y/nf3
uYMHQ+p2fHZFLzhR5hHIjWceTJNK0EcsMg4aP4ZBH+vhoFC3vFvFNkMIl1LjlrhB5V14zvrqylyC
MbI5hd3p1iGDcJQEmRuOZO4Zi4qh5+I7LJonX0J5hlRo4Uze5pxwMmOGUvqzIC8y05oGK5s6A+Io
E/GtscttynRJbG/CIZJwX1SsnNM/42hFjVkMwnFv5FdQVtuDs86viHn1IygvxXrTy/LWbFO2B4Nj
SChoeZnVmoO76H3J2iAL3yEWX9953WZYzsDJdTIvcf4QP+v06kPxLk5Mse8Ac7fq2bjGy742zZ1U
uYP6Mg5EpkBgnlbOUpwGUZbWxDyZiGbRofkSfcMV4zENwpFKQbw17gDD1mTCOmuX/FmX2pzGeaUy
Z0co+XW2VHXtQL2ZunODqQBjZPsdvoA3z7J1iSzHrxkmnkJ1SSBC9sYlsPanKdZOZEQgmWnXfsKt
MLdySCXKcZ1l12QWyUHgzBEKJ1OAAZZMONFsucwB3cfZG3BGPOB6ybHdaToI8O9zkCbL+pfGZc4y
eigtWGKflYT2mBuSv7m07xI4oFy39tPIqCVVsJQe3Tv14vuDP6hSiRzkpfO0Doz5kK7T1lsTmh3L
4N9tX4qN45F7JMUWzoljs6Hp1JQJ+aaOh2Oeex8SYNGfLjOE7UN6qQ14FyQ7ahOT5Za+osUIlZrQ
wCwUC6VTKfDe3TNqvxk9EiLVWLaxlWm+iPEdydytxKdvO68puUyU+UYimdma96yAqMCPEKw361yQ
PY+OHBjwlosAb07w7FgJs4TTKiG/KlQlbr1B2F9n34EODMq0cJ1HdEUhxzZ8Mmk49Y7Jvp2galnN
Eo/piTwkoM/AZbKzo8ATs6HtJj9IBLfs49iaURAyd5W95rxGCu/Kfh7p0XbDEm8FNnacvSwf3iGn
MHET9tGpITDWkFUdtfANpUY437Fd9pSa08N/jsXomvwJdbMeF3kzdNK3sQDzCgA2xhkWtpD4/5cQ
VFyymFHjQeCMut9asoroaqY8TTehs+q9jRl11Fi2Ugq/V+KYrpSNKbLNIhhbAjU10FG1pI95tctq
OawJyIfrHF/n3wcelLFTVQt7VmXVnKHZ1Ew75A73Co+YVMlOh6NQ1T/B9y9dLk3CKBvLCMzcGBNV
oIFD3d9vbBnGr4Yfi3HfIQW65V7yCoPsdHa39fciRsibEY+s9OOedxtPAehTMOLgIXoE9lbqLG5J
FXZ+RegQ0CWbhGIVripz5n/uF4Rvp84pjvEZls6GjKuqYOQjeEu4WodwNjdQc4hwnGJ40NEmOxkD
CL2P74TkFwjU/3t1Sw7U0h7DuORCfoV842UaZjv6Nro5pkf/UdmZhLMX20l8oYe9MqQRcVFkwB1G
rKRqaWTBPyEji5q8T7vCXnTM92Z5ZZLGt2SiAfV4VpQgemWYd4QS6l67S/BifkBGCII7EezSuhqW
GJz0Eg06yddHquYupRo05OZ5A+ghMvsFI8eMy9OtDSyl+1oil+6VJTTglwBKFfVM/0UZEDzccCUg
HoP2cVTQ+8Q757DW4AWAWJjiJtK3xT5HZEaIdebhW7fNiUKVugC821s8ETxLzjJYymciMIpQTcL4
BXZJdpBymUGwsR4km4sdtw/0Oa0cQpQji3AvSG1jOGIqBhj9sekDHQSV2Ax75jWKhzq6XrCTLLuD
PXtwl7gNh/6Qd7SXYoK2JqMCrzCCkK/R6a6kOUX3s1Wd5wV6mmiLRXUpxnNhXTLSP61FObh2Tsw/
dmJv+PzhL3xrd+EJjHty5XYnLh4TkSX0RzCq3Rrj4sQ/CPJEH3RFB2NiE2RtrIQcW9XzHZSu8daE
4wcDe3i16rhB4tKPwxtotpQ0aVwllTauRigco1AqOvtShvUgk2Bx+f/kJ9eT3glcgXLSUE9PvOTD
5ztov+9haO/qlVXEPEhgCas2ODpraMVpnsw+6iK5H9PBdW+n6yaQ1kU+mw4gxZPtAnTuDIn/cj+J
AFEh6nIqOsBlKnOTWsjev74KVAMr9DdO6eFGjLKIlqBh2vwJUX7B4I613aIFaR7/Kahzf44bV93G
3646hq6ZLUnigfyc+/nx2H7L/zM6vkDyXafZM0fRITgHsFsOxSE0KSDeW/fnuaGeK5HUfe490Tdv
kXwy7fzFftdWEWpofAzXEuL8X6zVPel/pM2UtEQgnfwK2IFhf9u7vTjkQNuu58LjkWkysdJhSetL
wMWQhHe0TClPxFb5hSTGkU/So8gYPX6oVPlBRs2IKlK2bIjMNkm6+lqcgdqJtLwhrYBonYe1HgYP
gz32sckYFdFEgp/U5cKntL2gcjHnXu4NvgFIdbnhigDmgm8S0SrtrfQEWrAUvjCdXeV6iBpMVYXv
hEIRCZ83y97tcqLxl9fHnV1LKrNZtzSrQStogDZ/ReZ8AxYcDcqzmt4ljgLyb8nBB54v/Rs6lYR6
27cEyTwR10o0InJovkl0LWCE0cWiPGa5/T4s279YPvxbmWAnN5i4exgok4NC09Dk6hpxvJa8QgUE
5boGx3oyJoLp23Lq5U/jYq+zz5weighARx/cgxDvf1Yxm3sm/qad7AmWfcvrFFnQh5RIz4XoS5h3
bjj5kzFRmpamx1/nJpzMP26Bzv3PfVbQfIUmefYq/Jca5X1i/YKPV+4sWJzS3Lps8cyzDIpmSUHM
/TW1M/bErpKxoT1iSMR8tm5OwUUdXfF9IdlWoVzhmRX7GLKSq+qnL0+4A3xo4ubQwK8hqDxh72PN
3aqUCXv0Px4T/kEMX+0W+kchM5Ejhk7c+JihKg8TqC8FF1d8LK+RrWueR98WYqPcja2Z4PWpGt1Y
glrGv2ohmPe5vpdzluTqcwRFDhQav2E02dSeanFFAqwoUeCIyt7mp1iiIFE/B0p3RSHQDLgx2J6p
WZl+0LS/YkKvJN19iNq+7J5WbSYl3cXI5ZKlyb4wjhAqZql5j15mBKkpdy1lAJxFThvvS0pWEUYY
jpoCNgRIRMrdz78XkyldnPMEErg0quzojH4+kc++117rR6aWuROW4JLjqbVTf7+j3qU6ajqk5aq4
RP94qam8TIl5ECVnXDs6YcF2uiDsfePt1ZxilUnxlcfZuFPqBdY+fWLsNndjRAV/G6MyXX9CSTD+
a0iI0TIROKeF69XRi5WGX/K6SUPFFVa9PMxrfku23m7lUgc5kBD2QseCY+kke8lwck80FouCK5IK
eAjfS4zZLalxx2hfSR2mcTYussuL+XmYQXfdV5NvE+tyiXz0fEjA2gD53I88xZmDP5jRv5hnaJhR
Xy8G+nGZNyIaqPGTMmmWN/xmpUn6nnhujBhxHK1sgzqC4iNdUxa5hXMneJhpDWKDt8fJbdeWeAv3
1gCNM38yrETvsGz0UKPNoNksMThz1kWKKCPm2oRTwufqODGgx2nsRYQa2vAYF6p4r4V7ziNxv7iI
C4YzuCKvv7gNQsn+ms4294fts8Nogyq9UbmIZc+Ow+XchJtvQUm/8MGWQYASfdeMNsaoJghoU+Eg
9qs54tBRZS3RjjBpChAKEs65lBgzJ+XRJA5O+I2ySljav66WAn9uLENdcH3r/u3UoY/GXK8K7xKy
EgH6B0UNQU1NkiPZ3TfQrqnWqkteCR4UOSKKpvOeT0n4H1/+911indB29n8tYcDonZOf1xuAFGXr
g/DonZ045QJCVLTNHmfn/qWUwDRfqLdRfQ7plHcsgHXWD7RjDh8lr2419OwD/57exYn3ICgodLNZ
U6oR4vPz7gICg2AGNbXHCivQj+3tyWAOknzVcXXgfYEKGcPpdUUUqAnBulXMASmCK86iV+xZ8cId
9A9+rF6kZmdsYWBjTrnXJcrA6h9IXuPmoatNh8451YL/6m9p6jK4zL7MjuIATvrKSDFuAX4mNwff
cFvNst660i5UhOj+3hCtZMEHaTU/NBO4ixGtrCOvWRVairpRfLJUxszL0yQIO6hAPm3t5TiS8yVd
RPqTMFA6aQ0R+qMeUbt6JsDQb28CoJ130NhyqtooTYNPq+AXnas1uSpWmONXTtfMJtUF5o1PW6R/
fTrXiCrnZCZFvJPX4gLAjpkeorh1pNHlhGlMx8zTPiOOJxtL3K7YEOb+HDYQzggFZxferT5KYKMQ
0PUvTNSYNSviL4LLSVm92Ya/STj9PflrsAa7iUrtvgeXYiA6tZbDFOTKo+unngdZ1I5ktCeGlgpC
uF2i2aXtBKrh/2+n8BoXgiKDwKc/Snvlja43TN3OMk5DTzrTpzqqW1j4/R4bJWHCzr3V2S8vhqZR
Av4IlQvFikL4hBLqlaOlvi/yvzBJqF6Y4T5HH2jMplTUPkJ216CECKjwpW9+f8uLAvFh5Z7t4zYC
tRyF3SDnva3rKowjReNgTkWp28A1W8K61SjWLhNRT/v3i2j0NnYnpjhoXJ45P89nhozjo9INgutl
t9GkwpTUcOlkgfqRNxkCYFfKfO2fx4Pc6w+C0DoW47OgtT36IOVsoH5ogP237koDnIO7Ws7Aq1e9
HICUh5kXWporN5tmkgS6aakngNE0jUiAKcR39NHipAB0rTQ4eNmp4xy2j2A6BXFjBB33+pCn07+u
v0tqPsPL+rkKWpt/JJExVXqNcw2NPVOUXuh3Jc1Sh//aAjhXV7GfWfWKx3fLVP/55B027881KEqx
2y0s0qChz3/caQXYAcrWBQm2cR2nrFLSt1AGZaOEdztorxZ31hKRDFjtTfvlpHp3oPi8zc4JRYan
PSY7PlZp3KMJl+QlMnCPmkzkFW6oNr+FJLpCgqJo6qiuLnGzwsrCf3Y/qxcaWRygCTxYyXOjnAoB
qlYqheztSH2UiEFJ1iiB7NxY7jUI9178J4gKiNxyhUWGA8WbgUQmasEywgpRnVsnxDJNXxFfvp0C
Evy8y2TR0CDIHWLZRX9y5DLNWIzTG1zzy4T6K0oK/5WL0IP5WPm4+aljT5/DD+icKh/gFuYop1fy
frkQng0P2MFE+XD/7ct3Q+qWOOmPavHdE5NCpHVtkct2sBCl93uPOqfzfLTqVYNvNVreVoKiDA2l
hr7kOyjg3JAIvR+uIdFO5YbNUm+jLjakNqnDkQTm1yvRciGlWgNupTuA5bUo9X5Nf93A8IfHIRiq
bdtsZZJXqpW3gXxlXFX67gsAPV9Z+17ES11EODLIbSywWT1MoMfvkO+36p5lKb/MBpIYr27iZ1OZ
HNHLJKYT/OCJsrT3ECjctV843bryaK8+dp7lh2klEWtEUp99tqD7lOIxEpgz/1++uzzBPoYWW7vq
FYXfaNSOkjEKJIXElkmsRgNVc0flRHlX8yYOEyC56rWQX6K4IzKjYlVpeEI5Am9xvtJ3y/cy8kUD
PS0ozBRQXsfVihu3OB386rzv0+eqYqIw5KijGC0Xx2R2RVxGUH5/LTHysrlbTG8P3jZXedEAx3mN
j1oSNGsRt2l1xGzL5rRzSXadbCvoc14TPfgq6Jy0L5ZkktDxP6DhwAqWrFWlFX9/RAhVK2cmJTlk
bB7YkqO1VOWu8qCMC73RYd2kY1BfVQNWhOcStlku3Spb/WL6HL19JlAQruuy0F9TcepDBFBsXa3m
udqjS1BsjWtPd9onjT5HFO95O+lnz5rXRIc1uNImZ+vQDU4aQYf9D0K2lUEcsM9fHcmWZrbByKa9
YlfmP2wUH2Dl6sbU+Wg8vN/joM6pU++1OLU1ygSVmUCbkqnTYyux5qjdNk/HDcJBU8aknboqkNUE
Y8zF29bfxrmSFo3pTCkAUjQcbAFBa5jt4V0UVaT6h/gJqdyZu4e8niD9Do5Pt3L8pgUJn5YZTMnD
M9mRA484MXG9jlMJkmavDiX5SxL29RogZ+vtWujqW08g6MUBDJvAfUChQfDlNLgmPidoVkEnjFwd
roSfUHI79BebgBzmg7JHO+SFLpI2IW1Ag8WPw25f5V3o+ptHJt+KyXa4NeQx38iHWJ0tnx1bjcWj
7AU7l/0BnhSg5BiCAK45kQ9JqvJ1/luWXEoMomaQq16JGW/Bq4bosdd5kelIiOv1rlRQW7ZDDk3k
bfSn3nnqA/efh8GTysSyShT7JzxwDSZ2pwTvYhW8pHPkyMWC/imNSfCuIMT9h6EXVTQoafVWdmEb
+rjeH3YMn0Ka4Pfdx0xYnctPlLn32fRTNXoFxp8DD7OGXtO80eI90n4iN8y5ZcNzsFGhcal6TlV9
ddKeBRyWTKHrfSqkdQcRMVfxVkAFWHKqKooBH/EOOMqfjIN2RXCe6uoopMrky/WJF12A/Feq4liw
JqFGJkmXMYjfPc/jhsL/Yf3xnRjSSv+DCzmPWKeik5QRdKfjjQNNQM6dcdOUDn4apJUM1223JyhP
yo4J50gp2QxSOqelSMNDp1YfHTCFZNmzBzy4Au4gaAz+MJ0nVoyXBhQMh2o+k+GuuGesDVUv0TIP
rFkCW8tAY4Jd4QW8Gkt37h9Hp3ydWGxnfkSEl0y/IcSzooRQzNcbUcuVynHqGrJi8t30s0vsTgIR
JftqGe5JTIeFtjcbRZx3WlbLHocOHP5/JhzpyK6BiF5urt0y4LLzMBaRdJE59F1oSpIUlHReRT2F
LNd5zT2ejSpFPNYLtlXosaIx4Mzcn12AGUzZxtmN09cswhIdr3dJj67X5Q9lKYL8tQUg5FuGl4WM
yHKtedzBH9r0bT9VZQc44ibkfPm526/4R5SEkVKG969kIzi35rNazwhRV1Ry0Fbu1Q7orW7cvrHW
tU4lLSrj4bb9SBwlUPzTiSDcXrqfwdQYYZpz7EPj0C17KebYWVaFQk+M2HE9CAu8wzkOmDusD0T8
hRYLJrWK+f3T+rAzpECi4MK7QrfNsY4JlFLjdg2zksSxdUYsJqkRw0yNN0HYO2T5ItVoah1XyPJ8
Xxw2PdaX6kr78cxusSHEW0ObcLUGhW8iP165ykZNqlOJN3tB9rDxz8CPI6UrLBnyDj7g9v74vrxO
Yd3P/Jk3x9vZ8RFKDMmnUsPbHcbqrW+gapnOTHa+cttHukQmBGrz1HDigYZISPM3xTHPphdkCD+5
CXGcBjx8ieVBLsPU9Ihstm9/d4D8v/902iCUKLeNEJ1bY6Acc0PsITKspjfAomB/VxBZnPh1k3Ag
kj9xMFqy1M49SBjqtyLF4CQ3luqg8otXdkGKzcA5oMpul8WTHN0wM0OsB7ECU3Z/R4Xbax5THk6O
LlGNyIzHB5oGApqQdpXGN8VL8c+T55qk5tU2bJgM3RttyMHF3YQZWX8eEf8frAn91YzZrHTo/aod
MRZBhy1W41fAWR0lpynM/AhGhfN9rKR93O9U2MO7BRmoUJcS14mog5KrM3R2BDV62vLht5lzNimm
n+er5eVgh0MdOAAr/2laobSw7D8YP81h3AkW5Eg53kNEcLph0XkQESnLSGnBzc7yo9zDOwWbYVkH
Zimsxn66DZImBdHrz/78aYt8AkGd6vKH2SvF39H8r820ZlnI1LnES0il4lJcpRFEWLqG+JGXZ7Ra
7fJkergazXNsTlig1AzHNDFmA1NT0bN2u+Q0x9gT7Aqq5bMEbMISN43pjhowRLVZw+Lx6AvlwyAG
8CY7DZYi747Jx083FczWP/zI8Nk6c7/nDPMFDb21P9Mt03iNF5zUwHVY3lY7uhPY4yxf8edrHMJA
R1q3qzoo7P9jbeLvN6ZPU+wgwtrle9JUxKAefJcTP+UTLIHopDlZCfiyNgPqew7ILjSeqztWHScN
8lVS4ogFIR+gL/A+DCCjftiEyvvyVbj3yMYQFM3mnYj4ppgWc2jqoFQgCabjv/HHfCqSUkPyi2qI
A9wCO0ZsbCl9oSus8nrTPL59MiCeKSZSiksWQRhJy17CmmMbvymmwDR6s4xUNLMFa5bmZw5ne5Va
PIWexy87BE4kD7rZhcTDvE2QUqfcT9VufIAaEst3WiJmzu5l0yJFhrciZrwMmcTeTIwtaOaDqeec
gUE0bGpsm9d4Z/YiqEN2hwehaLZ7sWtDO2HQe0me2DpXOR36LbmaukIDX7x1jgAdLQE7xfmMv6u/
OXZlIc69/MwNYG50y7c4HWw6E6PRJ0P4A9KpkU3mGF+IsgJYBMlVVhXnajwHmsqgEsl3X1oOhYtp
alxyeVg0shUaLTB7zjSYPhQNB4GEEgcDBk+X6omgA9GvKW3QPwCkz6IrK/Ha/FPIPE5xLwTmt5VM
QpmXMSaN5o5oGtN8F2fqlJ1xbOtUpCRbhJDmTFhDnx0h7w7F04QcBmRqasTBVPxIy0/wBZV6JXcV
A17s2OTCv03JpjonhAkirBqaGUthhCeUj0vs0Gyy7iDQ+KTWYxz2vCQvlkBq7zbUxW2h0AkOP1J0
kklmwrXIM6+kWOxlw/5CoCcA7LvsUyTNNz2Z0zb+yEePnorKwtxCnWtRuWoYyxBw/G5A+NMeXSpv
G4pAqxNi9l1h4mQANtt5Aho4YfW1g+MXOT3DG5ovtMtQEEKg5vnHI2Gh2orBIGQGQNl5F6VMhX2+
w5BN7UDR8nbLzJ82I/78FeErxdtB5rH7ypU20UzBlV4gLAp6v7KKdaQrFfydofTZV6PGDp1wCvJR
N6XQdPEMNu7xjQ5pKOYuKSNBpol6Du8NvCvKY4KtCe3dq+rmBzZotAKWdFzkd5CUawvnJHHIm9JQ
IK/THjvX7yZOMv0u6N5msXfH1XZ3AwXEM/Z+nZcptSvq0cdfRVbK1sUL2KtcI8nntSi55rI/Yl3I
vzvRvE5WEA4QAjmPVAQdPMt287EHcHkt3e5/0oFwd/xkoHpjszw1aEOm+QOkAP9TLia4b//oN+oq
6URDOjLUpYHr1y1TVtSJz8FI0encZ+cSkhJt0gyoqPh9KmhwwQhjGunewz1Y0PofGx+4ZoYtPiCJ
vaKI2Rla6WtZcIeI1waxQCYW3mBzlXbr0O9n0YQj9F97B42uBri3aqc8tzo6Y3GIkeBp/mZhpEnu
RxGRKII/te4ZykyGOBRZliIF+E6N197KfZxP7n/MSGUtzHQPrXmhtlEF+j01ZZJRAUF31yIea1ko
pg202+nYVaHjiRPGY5MVcmDi5q4wTifhF+8BmuwWda6uhB2vbet99lZ5iWlP36noTylbuDmj6JbC
sRVQaA20Y1YjD6reX9CbvNYFJJCxvqVFWN0dkMKXsvy8iPZklem02fYnJrzybXR3qgjDvTuHWBw9
OE8/zrP/7so3ROX6LfWnkIr3Cz/hOLTOFx09hN0T8l6Uze1fLS0MpDFiZH3Wc7CRjsg68bJVgs4G
liWd8RxxuEHJJOmg0VS4A8hzBBz4gqLoNHe69ukhqmisl8gFCFa2lSvJIslFBYcVxm9kCJCbIdkh
Q/cvWM8xyD5DAr7unxaGD1hu1GqBHBN5fqefaajrDxnnEr93lBZOHcoBgoo3iwcNASpsX9dsbUVk
j/ZtDNsh8dcMK9Q28QvI94AdiVhSRdIw206mImCaqrzgAXdb/iuXGxkbKco1lPiQL9QzgtlwC1XQ
iJoUtzuGDIGteIaJKKR0HmQ1DyfYYn0NNJ0xQ3byXpwLf8hRZy4+vOyLfIpbTgrBXJkybFp+0d9P
rtTiO80mdZZdQGbm7t0sjfktH7MBJZOKX479yBNq2k7HtjMkjD5Av0Xi0NZnkHlJXk08Y+Ksyt5t
QifpskgDwA2JzK++BLV4zKCaCydxqodjOYqZP9BRU9PdP3VuvYi/EdmEJUNhON7iROCKFTqWMlMv
7+O519ypa/OrIPK0CYYZ6Bu/m9LWSiSvjXzmRxcjir+YZLkb5/4tpaetqPCDQ9uUF9Sl2lFy28ix
9Y2UjWNzxTyEo4O5D8GiH7aB5J+dqLi63gDg5JnXlWgM2yUu25mUdiJC/j3b2TCAWghKf7vr/KzB
XSP4YCJo+Z6O2R5Qpdoy6Vgyuw7GJpugDEtLvPUc7IyPRRC4G5ZHS6/M4ZcdNxGDPrA+FaH609hB
UcIk3m8iPVrIqZJjn4ibUOLH5NBVFau3j/gYGm/ik1jst+HmV1J3WFTyiip652nxCsq6yd6Hk/bB
xUuHiB09yEQ6Hw5dJjJs3/3ll36AcqZI2Mhm/5hs+fFHpEj6M14RHx1i/0fH8T5Xe2nSXfKz85yJ
4IHh9HQ/AFoikY2iEQ0oDSNV9v9K5rdCm0JN1RFgpcpkmCoc4nPyRVAjBtd+Ahcnwm43yl89reHJ
XebTPJSoPC/xPK23Fp6p/s1GlETtjlhLMEhfkZAS2CmPY7BPm/PCKOLlpxweJ2YrhYcpvin5qgB0
gqyckgskGP+LRW+ydPE3n1INGCFtlz7rYOJfnBPjIkdioeKjw9JHAdCv+zv10/W5MPSHn26RYOo0
mDHYUO+YbHyBLZWgYnHsn9GRT84Rs1aRctjCv9bQ45P9Ya3y22CUfAlpAGkS1d3yg62jQKccLvd3
v0l0x1uhX7H0bnCg5rfRBL2AJJoG+pyYJvS2hjQn5Lv91FgFcwNzx349zzRnjZgTcC42YPcw73tQ
Am3hqBdIqONMeTvQgRIPdVwUlWGopYop75ikMKGwZHeURgu8CvUdLmN0LprVgw1MulM4yEN3IZHo
FDpFtMH46nk7dg0C89ZMO8J7DsZq+ijxyjrVWUdAEbsfQAyAEKXqGVhbIR38NUqRl6mhexPX6X7u
XKvkPrsRb7Pd8ctBM0X2yhIPRuY/RVrWc0yAbSnUBn8rpYoyapqgFyEZLpUz5Jzmvc/DDXeD6jvI
chwPGnZfzgwtfF3URrAEwhXjNTrcIl+XP8jqvEFGAtDuQjkBWb53xzLj3ju/NL80vSHe2T1kpbPc
A34qYzsM+3ECUOIup7d4lORo2lc0yVmniU2XKbxxL1qVFhZ22Ym8O9nm1OMup2/W1f+t73jMi7Pc
OCV5qLdbJLLU/IzoD/RyaofAnD3H4N6DREYn7NFXk0iAbp46l7fgVEVCA1mM+UxqvzlTZfu9NXFj
BwHuAQ1MbIkGIFtwd6DkUniHXrxhHiVA8L/nCEZzj4ZveU2YfWjyxFWqj58DHmDuFS85yzJu1t0v
OIqir6Kp61zZWe/YWPme3HfFndUumJwimlpYX11nZo5O4pyfaX/X2XzmL2zvpkGREPBBlgMo2CDM
fXyjwfCCTfNLCTxtW8mdlR11vCDHFnY/S0uT+EdHk3Q+gsPY42tWu0/oJfXltcG1iim0D2XCezG3
jP0CvlxM0xpsv2WkNjLLZmlr6kz7+z7d8R6IJqLeB4tH8hLxiqVSMuPK2r12mBJUQWnj/Qz0lpxT
543Rbfmy5z4EjPVCdSdhbVc593PPfNeWFRcuGEpU/M+N/TvBZG6wpJzi5wxxBgPD7kN/IbpXNnvK
m59cqeR/d2bIfl8mdC/XZ43bjuE5Kf6hL8EAqi1y8h5w0JC9muNCPgSNiuym5gfw1ZAIzejArIUX
uqKcW/nAw1Qc6102lmPFGUr6Z1vrtrIU0R0byYF4j8RfTLu1Fbo9Irl6s+xbnhmZ2wKaWd7y8FlP
LwRGXroo90GFTTjLFVj8DsQZkoVTVbtQduHFTPiLsxxvctgIIEXZ+XPKkPFHBGGrLM2aY20DBfLa
eL8etjPd3CYsML8OWcKWa+4TRdbkT4F2SGUjgMxQv7EK9iT/OtmKz3uBGkYs5A4MaGYQws9qQofX
ny8pVGmX1iSGUC1rrVjWUu9UZG998Vz4R1v0HGtOHcTJ9PGpKKUR6Lxf+J4CTElLyOmdX+rys3nI
rNyT3h4bzMkskCQJsHb5ze5/wvL0c/ypzVC2gHG9M787z+nqEE5ulIEwNsPPDEfxzj9PpAEAmCs7
oziqTZd3vOTYGBFKnAHKqAKpsQuJL2CGNG5cOvX1c6NxsRnatlvNptwZ6S+MJa4Nftph/FpnaEIQ
Vdw552AwgkUxdBfw1BamzNxVhrRW3G+v4jBKjZzghyXSls7ZPJlTXRf+rGP1xMCi5ovRiXUNPBZG
sMkkCyp/ogI0YpHXkhyMiu1e0KxlafyNpRibSonRGHKzI2MwZ5fHGVZDNTIbaol89liLhyXZeI6J
JzUdPnTw5CtRPgGwE9dbNz1vxIhOF3LA7y8cpZ6bbOsq1izFGMZW3NwZ5qpIOTZymh87ITKcG46i
7UC1Xjw63h9mRf7kH8Gw6Z7QDdhP9MgH0gfPu8aCAWoJZyVWN6//LFjO8fhYPoXxEYd4HnLOoV75
nOBch25F7/nYoFC3J5f/liJzEYRB8Nf0QIBu7l69VnDdUGMJ2R53DdCQarOCiXRgFbYBljApA3O8
YF+SnmdkCllmthZjsufmzgt/O6hrBmzzrBI3X8fyo+ORZRBoMrC/0prKZwqdcLORxeUCNWXaKGzz
ltNP4XAItqmkODna7FEsVbI0CFtHC0yS4ne4fUNrcreD8m67H8Z4Km3U5Z0RUBs7t4PgWipT6ua1
DH9RKzfORVkuHzjGYUdOXyfB7Or7xWcl2C2ubfweofxUudx51pv92Y/DaA8RU8ea60X/FswN570M
eA5FKI2Qd2tya0WhR+sYCkAEQCjb+joa6CoS8ISZeljxMaZe6SHQu3UdVMhCa31E2MwiAUSsp0UG
DnoDle/voiyUj3YoRnggCTkHvT8TUsd07Anm7gaq7QqPv/0PW9cmu22aAuZfYD0PfzK6wRV/5nPS
+9zyGoxeFFHquyKcQ2MkTe1VRQlQLz9jttAzqQpzIbTqKKnzeAlRZm/7dedymsVsXQUxxAdIjTxo
tjczttBABiu9D+csiOwv2hru96SZn7Dv5HRrbWkcuZs2iGAOkLbn/MynrqjWr3Hayo5uGjVHOOwS
tkNE6ffeVFfiGRX+9jlerJgNmAPtr306DkxxzZqkviwFVaX87fWes3JguxoUYHhszieHgPye/EAi
fjp0JVQFke2ADNEAztxqUjqs16SvEOwqM8e1rY2FltDbnHRTaD+f2g5jg4oCiqA3YvLB7MhBrXLg
29m6Dfo50DWVu7LVV2XzzztT29swMQfnTgFLIrWq1dxuKyd9aYFV/24oW35HYersYdOX0CA2iKSc
9gdI0I3A2gNX65RS/L4GDmOCq3dSbTVHt9BCt/sCgjl9umOiJoL0NBVCXITfBoudSW4a4x7i8R9e
6+R0wGvBvEWyRchBKSDuTqxBqMlkMMs6z3wMB9OwoyxReIdilxSyWT8lfdUb4lBt9uMUr0w5kIFc
AXewxGLYXlhKxd7i0bjjoKCVL8fUouSvIb+BlxIu0K1Zi61mVFC51z0gphzCvD5rV1AAL3BsdWFz
zQM6KE1MjYJrlAhKAf1HGGr9hge1dqYjS4v8ryR6SbxHZHAXYtL2Cav9c1ekRYrcw78Im1Us4u35
X160zRwGhv+VkBdiM37RzGDML0djkIJYKlnHZAjoL8oaxq8nPDraRRmovZ/SCcykRNR+D0ZdI+rC
di8oSR+6zrgHzhojIkHHbD2CpOtfLU4CBHA0MuxmpD621PSpZub2g94EHEu+4qNCUEg+y+UxaUSd
n+jKl2PkD96ItVeAw2QIG/O9LsitxsX3NoHRrjCIQH5oXYIj66u9fZz56UxsRwKYKXwmOzEyvD0C
VNMg59DI1OUtBErymn0TZK15dYsEeyfu2h/3nS4D6zIfYAAmPTusyDxXFhpsj/yaVl1L/K/9TW9o
EXojm5iTNb2oYxDwJK0XAc12K7eZMpvneMTPVpPgzuUBulbJyGCp5gH8PspTJGQqtTnhlofhT2Ll
d7kysPKFLVYQNpCHooV/aXphriWEb7xCkUvjYNgeA+0VaxlmQeP7ey2UB/SBfiXTOptWEu5n26qD
1OrnSv1dDft+6HZqSXMMJZyAWPTLjWcOjXU/c78SvO2M2kPkGR53mNaGME0IUsn9DN0xS6SUicgS
CdpN3ftFduGbMbfAC/iKKiExqOV2xzsyh19LgtSg6u38QWUKOlJ6ooWemsNMtkmM/OoerkPXQ6/X
BIpDXWOnxKJAtNQtU9rbcYRbGR8Wo8c/fMxq5XI0n0p2xaeeL4cxLdf/Xt7Yw0ndnfKjmXG0+JLb
fdqIqLbcddHY8+HDlvez6heBfLRCGTrtpzVddWUd7BAKoRCZO5KGEHzhoSpkzshNA/1RYTtxa7g6
wje75ZQGa70L/CtylzLbxnnDkm85TYM+K0C3fdIdeS4euHF/rimOdtWZlYZUxE5Zt7S0ZQtRlHO0
S3QDlVvM+VcNVSroDlWiFPsCIk/DxaWR/hQZkDYeAgokUgiEK21SZo00UsXv9Px2Xn11VjMC4T5d
k4r6xTqIa5S3ML9FPNA+/eBEoESYUi/RotzDQ0I9U0gloAn9nQtETnIxAuG3NzXfiicuvf8jnQHI
+niRQoH0fpbYfWHEPibENzKI2vrvAc+RMwG7rKSEsrQ4fMDw1BPnYrPO96ZlA7X9riugtz4vy8YO
6nq5YG7b+sNF8A/WzBR2QJAcLc3BlMi9DHILxJ3rUYR4kIbwZtZmEbiB1P9OEmx55Oyb0eD/wZaP
r1PKWZz3kgMpLDIdY/S16LMa9t2eDe9PAC7dVG88Ogrs4MQfqMRlZ2oPapUDDn7VEn2EG1Ci6N+/
NJJjxDVqOi8WM7de3LMqLKfvke6VF1qRhmlbu3mnLQ4BHPc0NFPKCiVHAJP5Zx60MjRXSPv3i5B+
HZlcbxuIKJc2hwCUq/zClP8kqJxOs5ZZ+mfbo7RnrLuDnxxr8kTj7F+f3iN86Kogl9MP1FSkaQhq
HUKiAlBHnU3mibEU9EvcpTPqdI+HF8hTaffPYeixSMk8CbfVz2QnL2lWR1yl4Cxs3VG2yYMX22Nu
y39QAZ2PbAOh+r3kzomETtlUtSDMnwUqlA9Dq+x8oVXEOvIAkUgawwfWd+c58PiW7H89EEU9tPD6
ghmDAfXUDbSSHtDoZGlFddjZHoOdGepNN++kbKHYjHGnvoZpLGCJWDno0pi/nacVAefMIBQ9VwAI
xMizF2LrotFl1tF6TvF8pnB5EoHMMrAN3iuKa7Bniy7G/OfaKlfaO74zMDqzUbclbYcYCusNJV5J
a5o97mQJ2OMma3yG61skpA8gL2Qdcy/dgB08kZAtfJ6xFEU51I0FzRwp7eoV5LYMr07cyXbOgCQM
WuRDLPpCfhwto+iRlsb3grvTsMr0sK1DOUMqJwKQkmB0Bssklkx06nm+YcF+AXbfzjnr5rP3ONLt
rjPEWYH+i2bOam0XxpB2aZbU3F7mDMKacgddtMus8qOzKTunugaA3/lNCCbZdAMnmh9K+dZ9InIK
6p4SxIIIjka+6cE5iGj0nBOGhp9r92FinoEF+H6p9VvjAGYO3cbjKPV5thL/OjSqHujOyPs2mroo
hEMYJNa+WlkEXctpnc0vSuNa1o5IqPA5GKST/gFgrNt1M4wqJyLHmTnc2u4GYlhXYOh9Y+jZEFYr
p1+MYw1N6lEBNKLud1+QWs7UQQL+GgWiXu83p/yBbWtR/FJODLZAEbklcSiYOOyfwnPuNaQOd+61
+Sd+U7Zf48Xe2TZns4B1TuLJoVDjIGcHEl2y6NF0mqINglr6KAVsFnJ1XxNvgdDUnkyC6Q6cFuD7
uzP2xijK9PCOruFdA1aI4cCc8xrOfq8IUISiY6/MY7YLU5oayFI+Lpa2afbAgH329Q1iD5BtmU1F
UbCz1ammsR3SChrDxNwstiMLTh6A3y89ZB5WnrERqPFzWqLCF0iGlhQAa2OHyKghHavtsX5bbx6B
Wn57+HmyTwooF5dpvDz6rpk9qruhyGwqZrCSux4BYex5wgJlAoJCjSg7no+f/0PeoH+JJx6uK/yf
AocROpP5kR5B4MZr32QkwgNyRVu+NdUqppzOPlaTRRFe9YgI5EC+9rb9gZFiGxR8XHqQNt5SFuWn
8w5rmM3k8r9AELCw4MoENu8flKvv8t32p/46D4Mca7M9VQiWTHdwhdzuq/jmSRwAHahQqpMVgFUE
QYvubx9oUB7mGqv8UmPqUZwuBVrg278h6AloKWd3iHBvxK04p0mxnVTvTddCLOxmDx8xPuacoAzS
DxW0FkdL3YT1TR1usaOtf+4TOmL05QnJhl4rFAMKrwX7nsvgBCEod/UrJ+hUAX8VYC2AqhJxmbTF
/yYDdd6EY5CoFDK1RjB99vFF7HYA1sW7vagTVRxoQhQ+XaQx6ZssXji5ovQMpreTqa0u3MKT3C4U
K1ppsGih8cgabq266chD3MNBTC/zmp8CE/tOkLvfF0v1Ca4hPgZyjJwu8B+p4wPm2Q21ZWaxn2li
er9pWrcSaGTXCpBnyseFf0fxcCq+baCIx9EUzPTP1hgxDUoXCSw94aPLVfG0h8HBSfH+oZd1fWhb
mfeJBFeDANwrNVZatq+mRDKA8Dwcz9ffaNzS1RXnvLt0vg7mhfLY0+sqyFRc5zuPAINnC5+Ou32i
80nMCV+6cLHqwm+uMTrkfCI30WwoYrLEkuR8HYKAo9/EihRGzhn9mOczAmKAsBXLsGA0ICmYaYJM
ldsTaeQUFwqlUQXmM3pSmK1NoTB0PHksykvL6qyHr1ejSpoZqT+QWUWUqTHapNMmSOCaxI2mbpUY
zfmRr7zGfaIcQKJlJ0v7agjZuoV/nOEemo1TtHvfHXH45zp7m5M4zRKL1wyR3sF6mMTiCyslFkxk
N4ocNOWu5QQp7X6juTkh5ggWi+wHRW7KvgTNuOF7TmFXmLJ0kARylYVcgGnzGZO+07fSzd7kqtY2
bMrVy7yYGPjDDyXT8vzb13vfUBOHg+vQJnO4vqvHW7/sjuS8ty7iTya5LPBap58dQocH+VCw8lvV
haic9UEHQggJkvcIlC0oAziinj8dQZGdJHjBdQL2q0TQmrJ/F7LIHTHaMHmmXC08Vpogl3MoN2d1
954wapPuRdQwKdztGnP1wugjA2Koru8XI0YE01OYiUlZhS6f3xGJ6cXXpTGzbsV6rT55VJqSm4OK
tGLKl51DAYAm/i9nfOZxKbGB9+5rnSc3paD3o+RUbN+ypgh5G96HYdckfJmaBhetg03HK91Vaptd
N5GqceTC3tlhd/YV7tnxYYfgoKe4ViyiJNk0C8ZSxv+6C8kPaYe+Cb+8n9mo2bBE4iG74N2bfZTK
c7fPS6DXVeyww0mMlDIRVUKhCV97e1WeBgiPyJDJZrxa6pMBzCnCdAlNbvaHK0HcuD9l/tQNIm6f
zu7i+VIhCSV+OJQwx8GjhuCOCoo1ndQyS7HD6+Tn5FGUOQt4iiLAfym/wbU+qp76Y+WpRsGA0ZWz
sqnPe8yDgHahZyJ6HbO4aCMnoDVHbRsbfADPlUHLAi7BmwWZsm5Im4BMgsodXI/YxAqprtZnleZM
TidpGqoSbvT5XGQxnzwwu6fcjOLt5Meg4q9Ev7rCYoPibqHfMFs6Ju3fHLxnKzSfOYvphv5SqMrL
MmbX7RzvRNn/ZDNzVhxa+9UBaYLWtCHW2V0gsesFQKyRjnV65nlaC4jB4PFCghXsxmTpk7Twehlk
b8BfUo0p+feOWYKcl07CSKQOa8bRytqc8QeGMhizJbezJb9utiGykCjK979t2Jrm8uAbnkO8RtzU
DIavNH9mIsHbU6kOYKuOlRLRRMCE96DiZM+K7xMQm6WZsTt8DyjQBTN9UzJa/NF1mT9X7gAyTKM3
eGH4bzO7coQP0dOUUcU8k7WoNFCKbdSoorWE7Jg6XXt3TxPPzFu3wu0N1byHuUUnnIch7dopj4Zg
4pGYEZAePtOjPnHPLnS8rElhi1yAW0V6zWevuPA6S3HJSNI1SWQ82JyO4vXUs+taK8MqWiAs+FAI
eyt5JTODhhA8ky/SyJ8TxZBcgCfNyW3oqIn6csPNn9X2iv5eF9VUkka+J+KWsHO+ABPAgAJyXg4j
vC7s6oYzXvqE4pW1XBCwQO7XtyVPemTydYG6eK+92uaGLd8uXyc2+yrzZzqPUxNYYRhw46Ox+7pA
2l3HQiwTztBqZazLHGAYnVVgAr5bfOM78zbWQVZigRi9L8WHQeZyb2IGGWSCqM8Ounn9iCbfV674
yndwzWd+LAUhU/z/NibQmnF9P/zoyTa28mn6Gi3VMAiI5mlwE0QCoILnUCPqQemEpCmMsaXlq1wY
nUpD+mPUgZmMfDAkK0gpzxM2BVszj7Cde+XNh0uJDDaRP40khzGwgLyd4LQ24O/dIwo0Fgya7QYc
UFnllGz1KEpH+/JzSBH99EvilRy/s8Dibo+eiICyFxncQVFOn64rVwBUCV5egTTsqGTbdaqpszxh
3sy+oS0BCndCIv8O0VCnEK65zWrFcxMxWGQhwJkS3MsuVhP3giChmVsZvg3qvZEToTf/M2J0h7I8
0rvsdntsS2bz5nKu3Se6DrMYIyL68uRB13mAZU0TSpIasX961n5iIKhbh2H5bCvE6/+70hm2bII3
2CxHxGENoY5fRU2a19vYK2DhmQS2vINx8T3ShOIx7j9qJCtFXxpdTOVZ/oVRea2XD1JVXjnpzmxB
iFYalKtTuhPAkO6nc7x4MHEBpwYUUQNqitd28krwU3Dcyzo7k30RzqUTJtlvri+hHxgXFQ/mLg/2
EA+55soRHBG5V8LV2YEh+OUzRl6Ykcwwa+b1dJj9/xN4Jw89UxosZ/ZG0T6HjvApnwfUyifxlMJ0
I9L+LkYmmaS78gPzgcW75lwRLUEOsR+zwc3CJjroY6jRvlSls1/jmRYx0GM5G7uW5dmvL4tN6Xxf
f2QS0ND1IffrvPGHwMZ6ndXz/v5/rZONmDUxsZ8n17bFv6E8tD/qPzoz7I/Xjmm0QNER4DN4qOW0
sJyWsErY1K6yOGQluU5JrjE4jFh+FevKZBrr5j1gucltSI+q66hocZPVZxSlrHZPA4Hf2ucag5M0
KcujURE0TukSoSTZ/r41OiGhZWaVS7ei8xA67wurp5UtAnlBbfi2yhLGsBxg0QSZW425xdc6UbuD
FgGdPeDy2Nfrcg9ue8kP3fS/a0djd242dPqgTGJIP8fsRsDOUln3YJXmCoodPos2u79r61Kx5SiZ
qQFcMr4/oSrCY2zpiGN9J1PZKCEak00qRjlY9Ro/7nMYi7sHbITdKP5WhcxXDQg3GQnvP6LR6DwW
TKF3CujyLdk3Tmj0g5AnKgX8ge13yEcFdRuqISoc2MaYQo3gB5iS82E9ZQTAr7q4+Uv+1M7IO4CP
CKMHrtlotN6DYy403V95QTLgR/Hbtf7rSfrd5CR4ZkXEajj438ddOirOPdLiVEqUeBMfedzaatZY
NveWiSBwedJJG15yBLGiP/zOMp9C3KS35nm9gHTXhxUKaGUxX4I7h0b4a/jykW38KhGk/5nmdqsN
+ormGQbp6tFCW6qvez3gdwce+K3tf0woOhsHZ0+CE8hQEgnx75AyBwoDgIU1HwCEP5VizXDuKWDx
7mQL6FemT1Uz1uBXOobpK51LuSzJ0LW2mETrzyH62hecA0s3uBLgcJB3S2KepGJfZ6G2rDUoTtcB
CSybRpbcuDJJmkUx7EJfTbvFTTqm3BQU8XlBHdTAxgCoOgTTk+7WM3vw7Xsynm7ICglqJakTDVfW
NwwFqR1HOMjTRcUgd6/laV37oMyn8tuyUdgB/4K10Miy+LtTDyjwcknExBdTHQupfpgtBjdp1GUZ
OIGUn8LaIH2ZaIa2tLE1K4/xYhdpGsr4cV2qJ/CcCun64C+XIjHwm+zsWRdzAPiZKLLhvS7JWHo6
vEp+cfCdTDBqu4NtCGPK2mMh7X4ykxia0aPbLx3ac003nPOzmoSabqvAh9sszyLX2aFcu8gRdwwV
iaEZ3ZzG+eGkFjM+4q8vR+ASYcO5qsSV6a16GAWe/VbGw6XBlHEmffXO4JuGPnwh7IM6/PkK/PbJ
5orwpdFks6pRYTMqiRGVFZom6+I66GHHi6rGrP7VQO/HOhiTmIvdCMFkxE75rczupNTasGjFAKJs
7eetvRnxaIgyrwy48Vb/FQE1jqHd31Ozl6+IyV9Etl3QN7PO0JnochW4ttWlEMDR5LfWLhD1VZeM
+ewQ1zr5gpvOW8rRZr+uPSaZBHJULSwppwhsW+DDPUVI8UKrjviAh8B7e9SxpSe2B6xwKR0WrhGY
tGBQP6aW/t2HwHpYtEKGEjlytas85IugcTU+zejJ7kYIh257rER7R/Znwd+rDxmJb968k1JMNzwr
5DiZrQ6B+ZvimtGqCVkO1SNU29uZyc8r7JxZQirBPnOmlUks6MlmsDSC+rwTxad5ggoMwwMKRR+F
avgHfi1/JhwBAJQVBUoDSuH1uLG9+07DvE+H3mNI0vJCge7NSPfhbktMmYVYGp0EivwgWEBt0uS1
S+wPIb02+9w6o9YsRqiBMVAcMD466S/FL4CxnXr2FtO1HXYnGhIQCfy5+7tWZtmGMzXplXCoAjYA
gQaEaNoGv63nhNBywFs7sDc9o2UGKl3jhM6YJFo25J0TuP1tEYxpWbSiHokSAPAB4h7+nAL+FmvT
t9Y20SffN/o6+BgPYYWVCFYjEsOSvOmJGz9/duPTAmcQZkvIuc+wHIo7We/urQavhAuy1G/dyZvi
6mI9k4l2I1FSXU3dZ5AGsMnCLAVBr7PU1jr9Q9s0WywDgof24LjFMMZ2kkzYjhYSSIpmV+j+uh6j
u/LStOoCRC/MfKO20sMxEFNsg9i0un+zXlg3UDX0tKP057aRJtBAOxYQAh8gzPUTaeAWkWKnaZ3Q
08V7YysuQSFL9XLgv0P4im7FXxHs08govETMryd2Bktq/B3Mm3q1exl7bRjdnJN4vTTx45Ox98WL
3Ak3GtB1chjukq+qfH/gL82qLFBga2c/Q9lxpLLz4FVPNoZBxl4QqPDhgDswy62yegORguTTslOb
8UAn8OYja+D7tnDPPMBI3eaSxnA/XPIHyth9vetSUNs0pwBB6XdjLEbZ0hxdS7WAfNuNkRKjM2zd
bGycuiwOwlypSv8b3wDvWgL8S6xuhJdEdFqYIoKLjAY1PnTpplPNA2QwlbhfCjkB6jXmN17im5fx
XCO1LWwkxEqskCvZcMeK11BOBcC8lm/lsTZfnCMLdIlcZASnF+xIIL7Vni6yiy4WaiIZ1M3GNJJt
eKfjd96AEs3jDxFvYZjymGmyCAVF/2ht9huzwW4ycN79hDMMiNmgIKfZJmZn9BeM9WwVfJ338LK8
P5wPsNst1yCNfSz4sb+LcxBEtZ8obq3pRKZGmqhs51f+go7uBoGjsL0nKusrjZD1C+8HGSn+E/Ty
RUCZnQkH5DOw1p92nQx8N6H5+CwCXTOQsV7pgaZoa+/+XVdkIyDfP3MY6z69EkgMVlpckMnBZ6uw
W+GM/LarCr8ftIMxumKkf317yaJySFIw3czJPiJgolHgkCKshskrZd+eGOTBEXRxJV029K9Ldls4
5p1ATpY7B/xJ0GDVpY0pUqsp4oiRMKfzkuVt2YOj4RWNLPRvAHZNi4uC71jPDFG8bLaPctsZnwlU
03yiJvYXZh+25P0adnuB9nlcxxb4BewFTMCqzdFo9a9XxfPBhDEUptPgRoxa+XCaD1P9SiAHRCHB
geU6P69O2kLMExDfxw6ntyvsGRC38mXfvaO6irgUzCTPYwRG0XYYSkpVg29B6nLuS11JhmYDItnP
wIawvXtW9aKGMYLIbQRRcxIQ1ZWlEPJC2CqU0ZD/UdAB61VswaaYunEdYL7X6OrtHHDSYYH6OnAo
3x2qqOe0GgjNoYsMXwV6Ux5egv0LFBLoA7B2ktElXPzRW3Rzjwu08CYRcGPy+HTYGZrXxpp08jzD
kAxfARZS2kSMu4jCHpV8WOaLwBkGf3ctEcXwqCX5dzVfsxR/ih6FE9aIiFXvao2syMao0BQAIyxB
f0UMB3DmZvn5VuL/Vxke+aFU6NE+0EGxMbyvM0GDu5ZO4Fzt672rrt6dyyVCkpzp/rSlaI4VBjGV
9u8rj2DU5ilK9A6oWONsVHQoH7OoW88PGLsSwSYQXO6RxEDghZLFxglSN0mkjCXlLTAsgf+8bvae
xIXvXp9y4hMl0RSlUHFyuFdRxmBt21i0toAP8w9Vt0DW9H20aT43+kvBIGP3cvQ1IUDEC0BS1PzP
4pq/bYRC48ZGD/hjgd3VOPcNDKPYPx+z4rTq9/kWYOF6uWXwoS9DYBa5R13jR3iwHTAZpsJylZb/
SyXMqmcD3VVw59WWzTSiIZeyGty8Q44i3Hzx07Gvo09zWdPOMAU8isimn6xv1juibJ48Y/yGNyZ5
7jyYBVAFnaKVNInlfYN2yZcigiiav5+g7vqfKNANvEKej2zP3CDWTT/ldzzkHx3VaqqUHP4DmjdY
7rcKi3QG5GclAm9Ohyd01xDefbIBRqQlKbG0IKfSk4umx+B0ZWVB+XAOsWWE91u6VL7Rr5c+7/je
xXgquEX3P6UfoTYXkHuOPpo8F6eLcFpYtQF84wPQgWyjgV6r7ObNhIppRxGKmOgpypJHu4pc5pRs
R/9JRGwvN5XB3b2VnMxNTd1dI/eAsyO3fUsxZ9+rrcagieCO/pd8db2j+MxtpFr0OzE+/EptAZqr
dY9+QUecBEbNcB4JLwbocHDDRJo2PAEBANDYDKhFKtclYviJh8R+iMoIQ2M6ZdbxKF3h2mnuvw9i
uzzhUxniIyxzwKnI2wNjt2LG4GY6HrsGxfyE/nksm3ZGhgq2X1istkd/KqnmXbw0zWSft01cTsX9
Um0w0OZxSz6i4m2GX9QHH+Ndy46LjiwAfnLfDvE62ZXJBZsLSdad5BOLGuuBiLL3+QevdZ0Ml/Ml
goAEZi4L8FTJgnrfbomDykTx9sIi9fIRom5paq0d8l/tyVJMEWtHcB6KfuSIBPCPzPX87OWM0gZR
x8DRUdEhUOx4AIssvNoWHjOhA432X2sWD204iiV23jYu9Gz8zEYB+rlqGWJKkv0hRfU7+1FwWMeC
Rxl9cicUq95XTYK/HlpMVyXeU1bjbGWJxwg/Yw9Xl3rZ+UThwmyGdXwTv1x8prEwG1yDQKHxDG1O
kURzvwv4tO91VkF/Kf07WoX4QoQWPYL6lRI9nLXypU4XkPleEROJTIAxVgjFN7ZECSjC6ZioQpi7
qAQKMjRX+YQMAKC+irQZOMj2MCfTsRkmhlplSWArbln6mI0wN1F78p8rtNIIhpuvzPt2E7eMSuHW
QiJ8QFg1iq4XxUDOKZBACFg+EYeA+MdeeKDgXSFCZsjlaRYzS7vabQPdVRt5SmlfB6ZJ1JZFNwmV
f1A51ccyQN8+jpA+3unq2mWB3w/qHwktdScZj8mMQ9TRnlbyekZRXfO0HIqfZ9BwztzsKS04HcrA
2qXzpyjiH0UDzlasTGEvegj8DX2FyL9x9OlCCyFndJZsjA9fKkRRcdnrXud+q0L3WyQCtLin/ZAS
hm8LCqxAGh+c/yPQfNJHPNaGgLqKeIb/hWJ2Pko5k18oj4rK1cLKfS9sznFfhx0UabSX8aZrROQs
G279F3gZ/AIoTrbscOo4/5SKnuZv+CPj1aBiA5xl2qVoJ1ZrDsqrzupLrTScZEYPaD4z6dvGKcme
T4S5xvam0S7mpgQgUdU89fUvumsOANcD6QIf7+CPBakWsR3mxUH3i7LPc4iDvV7eZbG2Pdd17hFE
xCM0xJUOSWQGopwD8VsKv/0/PjA75f0JRfaVx6gOy0YV8ORjIQqFShgtBFcZvLYRvSs0kmnwc7XB
YtefkWzeVA6GTUWdpVTgUv+aRJVHqipIVS8bgIMCOVWwnwe+4S6LXGtpmxypThL/BFkgrtVEjSPr
e/yAIuZlJ0yB9mryGdadPudUJWMza5AZflHPI4Yq03U7LhsH1BmXkz/8q6ETxl9m6bLTzttlupFS
7JQi/PLpXsdYqsFV3UKOebsjPnebLmBiLnxYHeBuUVrWcSsjfiSCEVLShofHpeCFc+xke7qAzpOH
Gvzg1MA4mjvH3RfqGaa6aXsUBBH590+E5lz82hS8taJBTIy1d/UIwN/2yHZiDVqNQFyU/i6lCE6F
Pk7164it8sSmugLc+89KVxtbPyd0/9j+BhjCe9YGXunCA3tpUnj4XMDTnhlA2WkSs6Ch3dWA4sRL
NMDsxEH0uZ9JJ9aP3weNncOOZ/YHfKILUz6J2GHhzLydO7sI57Hw3YDfiy0+Emkv6lG4MsFCooXI
1mo6SWir/ss7SfxrWzaLpt0cdtIo8yDPCtCjYYOpTjDR4TwUaNM9YiUOXg+T5f1PmXRTiFK6Od1v
NKJno38N2ebpt2ZMPiIHVz8vsso8CNx3hCk9C6OKS1OKDYD+VGzoLohOnqWFD+S6OoPSl5c/oSEC
24RsMOQxleDZcz7ZvfTQYbTGiXE6/gNyYKVF9CojRJ0MmmI1MNQt42q+XeVCPHtL6prI7BEjyi2H
aiTytyHkaBhmN/4ZDdadrYVdZ8rGiL0OeCpXY3FiPCEUp/fA38Av4oU6ZwHo6TRrarWgFYS1Guq4
TicPFU2wamjGIioGv/n9i5I7CU9Zwi5xvISPHDQbMLM3ro29l4gSOKPJekl1p9SieMKtHZrK3YDO
Rpuz+oGGJESMIyEeqIn/bkHK6Cgev3NaIpv6UO/Y0nZQ8jYcGaq9tj04zkOjMp24v+mnlDAxTFzn
U1ApAYjhPrpCZK/wkHiN6tBIFQW3kPq1vCek9GLrhJYFhmaxaJ+EJXctUkIe2ydtttX+7/ffKH9W
TD/WkNiXcSf2dHympOl4G7k4pObsypbT3k4sV/ZSx8a0nKPeSL6Pw4s18zqX2oXNJ9f+grtP/CRf
2qjJYQ2OH5RHFW2+g8S5ldFgmasqW+I+iHmy2Tfgy+XIsvPsjx51DOf0wgBXK6TQbFt1kT3oLB0Z
CEaPJ6bN96iEzQhNiuKHilM5PHfUQB5AAypfS3yAlHg0u6O4X4ekrPcOS9pxOb0Eci4PckhVLSkp
ILyq3G2KMCdS1oP4oy+vSiBIWkvukt2BTp6OpdpQ+FvhfW/NGbukJlqLDM+w7hEDgl/inN2yZe7R
H3avx3ReHIU6ZyJ+TAnEaBjmF8EBvzsMbguve7dz/WayI+iPb0fGvniwmTK17G4jLrOv/d3ht298
aREfL9IYQV/tU1ASHPj7FU4M2Xs1l2hQR/AZnKYy1PGLNCOEOwsntIFV0oaMUrvDxwudNR0xWkCD
NQfqMhbYS3O2o9laP5Tt9S/pNe87y28arzKRMe4iigmsiPBfhCOGqngIyk0qjVlCtll5LtQEavjh
eBXj6nbhiPn5mb4aTKYVyXflmv/sDKWUFwEFCicKNPnlRwaWiAkJY1nJbNBOc3PA5phUaypTGGfE
I7o/X2aklOVlOR/ELF8ti9DJI+tqJMrH297k0rErMajypq0jBcaBmNhXANieOzwv5fMuoi8rZtoW
uHXrJRmo/uzJOSymQYXEJ0Gf5tmepSFogODWW2I9zaUUxr3krLAJuGeV/ufPZEi3Hb3c3cMQFG5l
OssQdnIo/HQ9WevMo77CZKxDJ70EVc6dBmKorEtNkxKGd+tn4C/Qxi+7do0PvgjW88hIoCgMkuA3
PJ9VaAUefzhw27D67CxmGWY/oin6ug/MccxmGzEN6a0+eXJqC7vAXYET7LL7xnSxnY7NYi5QbFS5
aNRpuSfBK5h0vgTVkkjREnSbZp5bh/rCO3Py+qMuaFEjiflnhkcVxRMFiOaKk0deoRm/65+J0B+J
6v3pdQ6w4YFEByKwmI8aODEEJFh4YYFPl7TQPdUwwkIO/9dUUGw0vnZHeBX7gKBKKekdpam2l8dr
NEiktNKbF+zexBHYgPv27Fy7QTexdftacT11f0UKvMAncG3//uEc+WoNIbM231UPL82Yin9rbbaV
ahICxgdHJwyhooKh4MMRbILeVbPPbbfIDZezItOtvNFKW/f+dOSzVrxmpSIw9E01m9kd89D0fgBP
Q9A0VcpjDtzVaQQGCICG08pX5msMjqCgRzLm/O+fHDGo/dQ4hQ3t/tJkpt0guNl2CISYTh34XRGs
x+bhulE6DB6EjBIiCl8IxVozPIuON32ORskhcM3v+VbBH/C9Slh5lfLyHiqH0LBaG1KVoVWZ9vNZ
IUZqwfz3FsuxPvkgZ1bfIod3xVq/RyM+ebgEQ2JThIg5p+0LvqRp0/jZArkYz3cgCAfoZlnd1yqg
cdTo2/rvtJxXk4stnT+pjfdrDpynK8mNW+Cq/kzTKE216fTSZbEGHL690KKUCAQRc6AaRz7VPwyN
dmsagNWZwe9rpeKpxAoABs6uwb1ITTfPZSxcXMQR4KeKcZI2Gj/A80XdLUXpHnTI0gfZ00ZU197j
N4ggTw54w/pssjA31ZbQ67TZo5XRykWwswVPvqRC2JhoDb3eAvF50qXT1fY9sxPxJXHMOo+IASWk
yYQGFlwiJi+fMXHNBB8ho/fHkYLrNlFamMdCzRMYtZphXS9khmzVeMSd331CvX/0/TUiNwauk8AI
8DMMbaTc0vXOs+AqELUDzvs0ywz/SDJeUrW/MQ2dgD5fRbajp5ml8rKwgHGmt5Ckr69+F6vAwjfr
EkpY0FOy5X5a1a6FR2UedIVD4WN/1lYMXo/Ze1ZKHBWSoe8iq/8tPfL5Fh2TZa5t2M/GRCkZrYkl
GaPFMEFFNJ1lzpZfIDiqCeq60WcKmXU9krhfxiqbY3eMd6vg34Mh8FPCgOjriIsII6DhQy4jQePz
XbGsqeESm6dVB2stST/QkAyo0oEzVFrdMFsEbSH+gwAYighS7yftEKCppPrsmN3u1oT8H6pYCJFq
xd2ZpdTv22RY7QAslHv699D2ynxbMdspCItZ15FdUrdbsQ8wC+FWyhMzFCv7gYS/YIRy/uN7lVUU
2D/QSQw3LpknzjXwNsZYoCjA8rdt263uAUR+XompLpBe+5V8QL/j10Jf+ZrgnJB/YxHlrkGfnQaR
9HhNOkGft4aMEjZecBUV2s8RpurFccShLfIXJ9ZpcBxzGFb3FN4beBf4Rg3wlUXfMhWwrLwwuyEV
ZJMTLWgQvqe+VIVDRDYRzTVBQqB9diUwDtQWM29qd8NPbR4TKaRciBVDNfaf9aXjLI/7tZDpIcS2
gfMUrvbSZvhjjrNodCrbufncmKPSocV0r0Bnes81rBAomds1zJDYAwhIFMmkm4Bac5S0YvCR60Gi
siztcMgwp9mOxlwEyjcK1r7e6JNOYsVDufb33Vs2mtgUsbxUukQz8RvGKpg7XkGIBwEFQDMaazGN
HmfqSbhtmzDI8PQItRg47lKIOSWjzokWzbe6mcA/UW0M+t4ShAsU6fcmhVmQR9laO90Zca8b3Ozx
ExIXhjCvHfsPIaYbZ96EajEjPPlYoUNs9WP0GZ1vLnyFrhlAPNLINHSFd0SguI9Rez0dzrWcuE9m
lJfw9ZPLaCtsO50aRLawBVpNckadSGEtVEFDHW/np3WT6VaeZykM5F3Kb+d0vGKmlyc2h130sOG7
tb3a9BgerUWVloMTtImZJTr+CPgNofypHJq/UP4oAPbBI8RXFY3+hE/cc8KSSZI0QB41g7k3+AMw
oP8SP/Rk10s0Pg3yK1M+u8vUSsXtSnVx/xNhtVe2gK9rGNYECrLaJeHMkMTg9o67cLcxt8+I3MvU
Pv8u26o5pc9xYWO1afuADbuc+ALnVawi/Xp1siAjOeCdH1NBLSuKcZgO47Mkh1v29eCs9m4Svfj4
V3QANi6D8ZdMZl20zl8Hl1jOlGnLrAh/7xut3eyPJH9/IrAXypSsXNjTs68YeJ71qWTF3QRRgFqZ
L66wcc1Oxz+mGeRqhfHG3YtjlsM98qyef8M0DMy7se841Iu7yD5QFiiG4O06tu8ZAnibXgbGJbmE
EVoooK80ue0akSsrlmStHafQXDK0poTIWgMaU59gke2wD4ydiEcuY+phMnXkSBS4JHq07VHOz1um
4zo93NwL91nuDh7G+aVQZYP8I33b8tL8xO/E403UlK/UhIk+PIpJrO8N+ePq3zGaSlMS0QyU+gXN
mBrAVP7d3RArxrCvIfbplhPxho/yWEyCFhRMEmEq6maee2EIIu3+S02KjPdGG6NYNl7FlvuNsKHH
NL9MYKlIajeDWA4vDQwSUxeFubZRVfW1/bsaFcSuaipTHXfi6eMptvzfYigM23b+MpfIWFl/Dhah
KpCNq6PAMsBAGrTwJNtTfTh43ZMPVtjwDpC8GBqgG5gbHqF8ISaH+cgxnRR1zuzaPfOYiYvpg+TS
SCFxlAMNteWgpL6NkKz9MgUNtUJpmDi/OQ1lgABJw5J3nYUEl1zjNffwv3/B5scFlBwtKzSsBEz6
IfFpjGpYdY/1A1OOOUL+SwA2n7+sxexBt/Mmg+eXof229oK47rasg+li18nFkz+n8HYMgsSYWBn5
008FhwauoJevRmOYZ9z9kx9uqIYD6IU7bzIWUpKR6BhGGNnwyMnMYiMCxhhU6obF+42iPjWxepXe
TsKL5sS2cGLBJ48RYbz4uPgFM6MQCAJlMb94zvwqacb5awD5hNCaBJpGidDNlmvz42kRxaivN6ok
gQqXweYjQfDPUq2c0f3jD6WZj28AgSnr7lf2AtBm84J0vh3Q2l5SQGEAdpU/bmYS+MKSC1pxcAPI
pc6H1s9BxhBOlpm0IM9vlGgaL2kENVfBSrh6E2sqdlK3A6oQnMUHw47KmwIMv6xG//sngx/Y/yiZ
DxlsZh5tWrMbJY/kRB6cXcrp7ioRF5zHc72TYLN6urDAP7JqDQCw2SEnrUsv4XpqOVDOs/rrRPvI
3df5+a/NWOBd+bFxN14H3za0j9stOZmBISN7ej6l4jTB1bUmqyQkIwxCIBYcXGR44VQU0WoW8RPd
wQjXaOkCOfREpgM06T/NBeNGwqLzlgeoNCzCoRxeKH9045GyMCyyN9PM86YYfnuC1dtIYMtIpE0A
EQ8r+LijRnUuIPZhYKbmm8rwNxqQRVMdf78cQa4wbQh6y/G3FFEBvLetJ1MLYNVoPQxXE3EYjj2H
oTPQFqECaxJn1QjwahDFrprs/INJmOpOUuSEGSIPDmkXeeL92SS1dYNMtuZJOjb7LEKLxb1wF2B8
cIU2S1JQp74B9E2abEec6RBc76p5gQFnsOOOlS6jNoOgiCcdvrLLhH2Ux4o10uajsp6tDcwJOFZY
nrXoHRuro6ZUvvNMjdzAfYRf4BqMREPbooqK0hnudJco6fuBBQCaya42VqByeY7g3aWwyyJ5z0xn
pltDrEphyITYeMMjVS/Z0J2PODkq1VUHrpqUJnFPlfCdBIo5Pd9Qxvg0wBwwldUJ2o6oUWrSwgiH
+skXZcoxgSoScCnzMHkIsn7Xgj5DqweD3V6sGfRIxo3yLvI1y0qwPvioyDND3rIkYvbc5ROoz2r+
uiiTb8Dtqa3W/74VH+wW93//dP7g/gehjsNAc1LOhChedKZm4rc1/e0Aw5tgyLueSbEQgp8fhtd8
vzxPkncHGPKurgNNABirCIWbUEt0sozq8n0ssHAdJS9nK2hx89I7NzYM2+mXdnStogrRrYfOArRj
POAYy6hprPs+2RaPtKf1nekbXJho9bayBRXKc88ezMhQAyISxeOchJ9rIp78sJeZpokJBEVh1aCb
H0fiiYOxlZfuui61raE4j5gUL620TSA6mGFCGqCRj2krkLqFgWREmM/zvzb0LDCO3ipeF+1WdH+9
FxdwZp/Oy8SEwn5yIHrEaeO2yYw8IlK4XxtWyw2CD606MpuU0upWGB3LSPDgOM9hx995OwKgHCnp
omsPH72ndc63xp4NuPbA4YSRQCBIW0KkQZCznuATVNV7t9Lq8zkr66mWLNdqdUvK9S/AyLpGR7rH
27hchI1NwV5YmYPe27jsqRpbEm60IUL29rjbZRO4dBqwJMPixYRSbFWGlNPARvwaxtIKc37RJa+0
vD8DZmfC8st5GZRaOoV0vbTdD4K4A0Up2mP84hBD9K5Asp7fBDihvoNkFd0xdy+kAfoibknpT2Q+
3XdROPqj4WocFs8GHEfo3H7xVPjR2QF/v/kPEqFExHd+MMSaz++aLVjq62raiOeNJVT+owC9rmIl
mAFfa+zKuBs0giyNo0pzUJvHGH07GSPZbbiII6rsfiBpQPinc5ZIGa/PkwZ41KAE2MMnW9hsiSao
jibIPsikVc469B3jFszzIo3FBiR7wGNnm5yPBCO7A5pqidifp5g8cJvs/rNUndWI12lNIKnjaY+y
BmQhhHnmbJhch3uVXV3lGeiInlK7e59fPRsLXLTHPkcMX5/a6leVSwlOUKHKaMpHDR23fuKCt03I
AYq+DYXQfUiQ9NTDoPR6hJZnd3xVS2EifPYvVlhmcKN0YaqeaXYLU82WgIVeoWcKPOb5Vu7yhsNS
RBXvPEtfX/PHwwGw2h/EWt77F5XjLe3ci45zfVtyYuQz0IyjUTuBJX7bJOT4mwJgO5dgMN7lWKXE
dbw9s/MgQO0bjRxcFyNU6jHlx0RzxjO2Vx2snVdxkR7kxe8H5XKj96cTlspcslsDrLJzfW7Wkz7r
oecUGg3Tro+RP/CuMRgSMey4J/1sCsY+bAYCaEPuYgq4CXtbn5yY15BLmTpm4T7LUaAcIGlq2P/h
I7mvFrYqDuvWsimIydGI6ei0OfECcL5PP2Q3LgVIupFah0eW40+liyU31Ne6rkAd+lK4lfu/vW8b
dDosD417W+oLM8rwgwUoOAYbZe8YZ5F2+didMMs32O56ydF7tmXJsINsNRZye0TgPmAHqsDTPjkf
lMVxyOzInUbiGHXYNTS+7aYnghAz31Li+nDw9OXtbgT3AQclGvgdbibPPBaXi6Ja9w+9II4pqATD
UIRswrZK4M88N0GDqvBbrTJX52TddtI1G3rCoSTSIwMLIUIOPHWLTkheX8WIMc/91PGtoEaofefc
ewR9xkiAM9FRYp6EYNojb42+ecXRShkVjbvhA7wH2P8DkNa9Az5yS0kW0XXXU8iOOu5BBMKf4Kqf
tjaj25/fAcKWRMdSo6pOPJiaa5a18HVysf5UtoKK+gqhNddgG7aJBX6zNwey2ehXpfmGa9reb9/3
VKSsRTNarbjO216bwnr7vnxQuh7X09mAp68GpHQaz+5YqU4r1i4qpiPLzOnDmKondrbBKBU8jWJz
NYGVaVtCylO1dK0Wiml+dmWDBjRo9sxYlCGEpDhjVHUL3OFlnNemq3rF4JBrB4E14BcHRNIc9Y6Q
f3A9aTgeHifNtuwEkEqlEtz69v7Ccf5MffL4zANd5wUjo1oMnPz9hA3x94HA/jN+wWnyFNigbaYJ
7pAK1+IZutNWsEiRMW0sYksOVh0C7XbmfIBLX842A7rxF2PE4qi1ASnBlUc44Nk39RKt7vJ2iSHx
mR3zIUkGetvISdH5rPnWKsiHjpjWntHU58fqz6hKknrAUBSGkqi3CDOWeLKlEcyNzO712AlLCpMz
9dJTrVxQVbrlMOgoYl5r74bMNKFxZZDsFjZHRs9RJc/uFIzIhENLBR7zGLJmWKM+uP5l0kn4vGmX
M2CLRJ7O+K529qPdL9YVKTARjyKDJQS3KacatyTz8xBzK2lxNXGy8B8+3+XNV5jjlUHOtcOBMZm8
PlL9SEv5aIdPVwKRJSywgKkacbZE2/iIqfQwYMFj115Wx96/3XBGSbr1YR402PWopW56vWPH8txm
T3edimrsIoUFXFJJbWthXc+1yZFLHBgbP1Q0RQQ5SYsfXHlHN6vLVCN5vFV/nOGn7zrLBe43XEay
UinPq7vl+BC/f2idFtfIvkJHshe3l++mRSgDtRPSVZIlxQd3fJxW9bcPpZb1LOEr1CTYpDqzgEiB
V2ihj6cjDr5DF2yvbM02SSM/k8VGwj06A3a/8kO195AvDUzWwo6d2YML6dK4uahYtaYHGchqqOHQ
//H0KKDh4psqHzaTsWbmaNNl1ClujV4LU9RIesHq0cMjIPnhxoH0dw0I5PsiBeqc7DkQG5DF0RVy
P2yxqxDjWFl5CMGTE3oWQxb1vSPJRjow9jHUyiwg/u+G1ePNA6rAKxDn0dEDHgczUGNYbHq0ov45
wEO88Fgj2jBjl2pQMH7r3gq9jT4U9yXA3xM2eNTGydpwnugny04bZwwkwSDJVIagorIL5JLYrdb5
XCasFbSuoQwGr1Sf7eqDMtcjnNVIItiMV8gafMTFn0G00KtPUJ7iou6oi325VibohNJsIFDmcX7K
0Dit/17FO64LBW6ZDziPiEZu5ZGjqCVKioKNYOmtqK2m40qnkq55jI20qAsnhGnyGJWh0B8Qrb+j
yGTUgdBHnyyzED1oAs1BwWH5tvCn3n6dA0SGwheKIUeRS/Cq8mlMpGtB9KORs0QAvPh9Avlsfq4B
C9Ximh6AHDXWncTKlsTyKgfhZmwe7GfbTzS4XlEiSKpaXtY7RvFzWsU0llqIJU9VnUwXk/XCNbd7
mDgIUO0r8MMtEtcECpwR0LQd+n5Rl76zZw05dEdrygZqoQjdwppJxoTq4i/h9+TbqN0DbfCndFlT
AAWG5xC9CCAiwk9H2x+OB77uLTLam+uV0J9naHw0GmRyu95S0M7RnnvR89Cz7oxjLIDdORQQ+yxU
q1WkVNNZvfRJdgEgE2KcXaaNacxmU5Hn1TIEOBSof5yvEIbOJB1LX5cy6e05kpYc31510WV1OE+V
SSCHV3NOJTM0sT6rb40Q0Lb6xlNMN6GKKmUSD+fChxQsEutOxpNv8DockT2qCIeHaJqZPZ6EKBrQ
wyhqWH7SW4G5uGgxA/leDmXWZifdPOB1Fv5R4fsTATP4EacP2APBd7093S9Oczy4rq9PARu0vkEv
PrGpTHauyWCnG7VawLF057oosWZAezxTrPE7k2wPl9oDBTxLGLO3DYi9avL6Pr1DLfXb7qKpjl3W
Zujk8+/mXlrdbcCAHXF/2vw5ojpwmB02BwvHn6yJnMWMO6V9zZOOyOKXdrj72ys2vhPtOyY62HdI
HB5dtNaxIrAZ/afCbYXGOy+GyvZb6PZ42eux+9JYSHHF8jPxJeJ1E3TEhML5/kbAOfMmEcmd8xPR
UBmlpVlWZKILx1oSu7x+moHGstmcsmYw+jefT7JjVG4z3itu9RE0Myug39Ml0rYzGjbf/BRBJmc1
kPd2C0xZe0KFR8QciiI3jsN2Akip2zAasBvNzSpW4Mcrg6osWrN7KL1GLyVs0PzVxWcCKdKyWDZd
cPnUgGFUXhMogVKDf+qVDlA4koUt0vH45sKJr+LtG0i1nCJeCgjUIoL5QL/5nLTS/9Hn3ZhyDCGM
RqrYfX/m6vJhcE68AZ264237/uSKliLxQ0VXey/NQ+aJnVupivVK8vxE84Q6ntnVa+gSp2Jz0Oq7
QOVJE0zYmLg1pI9HZrcL0VJiIcwuKJJneZQevPghiSu5FG13jtkuPuHmgZoTw1YLNdLkDL6cTK3V
s4d8CS70iy1SlMYwj/uJexxwYuK0cx/yNV5IHHn0WjybmjXlfBS1PgE0jblEIpK/d08pDR5a9wF3
6gETwAb58+xgoVVGLZBmZFsXDO6czUTB43MT8Fg3samLim8tAzJtHzwESWERQo+Wxjv+GpFSJDIQ
+6jo3L+HlqF6Twy0Umh++YOysJVZn3ahI13YOYYCUCBN16/kQW1wOyoXoZfpC9hJBQhObpKzP6yf
bkZ8bKRgvsgSbhsZZxnqpO0r2zC/oUOEAPQiWTNY7t2TBC+O5w7nfP4ZN7jMo+Q9d6mS+aDbMKT2
yA4lmBTRw5UL5PtFLoab55oeWMvHVHLbQLpHsSczc7Hkm1cCHBQBuZAv5YnIm79m5KhCSwI7zNVJ
/Lg5wn4v+2ZKWt65n04q/6sbpIrjGWW/G+0WVUF5Xb1o3Mu55r0k7/0HYhaIdYufKus8HOYDB7Ez
T/szpr3qgKjcgqUlqGhlaOudAIut8NSlptjTbcZbdcMWl1mVOm/ofQ1KK9ATgTeBgydVqJUkZMKG
8u/+a+/FTGJW6LqULRlFf8vqYEcTZPizWA0LoBph4cnjpcvqY1w9L7e8ohTskXHV+gU8IkyCPDnP
pRioGEA3C4JaMw8WZlAdtygA9HKinYtRhQz9ydVZ1+/KQpO1a4DIKOvLANSmFmuBZy38cwMPnqwU
EmyeWgi0WCaX1C3MxZmMKAcu8AWYuQRFeq4g3E9ZHOHeis9heH59as+JHi0XjhSnxUHYUrTWSQxr
gkVl07vkookpraRvjkXUwb7lBm2UHA0AR7NG0nfNqTicjeQCWhyvlwJdCj8YeMH28XzmduaDYXNU
FVd6wO3ynVBAj+6QmNAwY/g4EYiikTJXvAbAp9npiM+IQKJQaLw7DL1ze2t5/VarvB3fuR8VraeN
nm3O8fBwANAAqoI0KhM3tDEUrDT7sH6cM/I9LBXQuTjOdMATwG8KE0bovM5ejU+htgE2vh4g5yJH
MyzQVXPixGrUpm+AlEcb5SG2vG6mdTn9RNu78uDgWatmn95PFzVmnd2uUzpjKCD5nuK3BL5kJjlV
V0oYjg2xgHZOHjwwFWNzCEVamY0zz7YkiCvdke0dED4uSCKIccvczkdOo8re568PMVOd3i1GFQ6c
PcTkSsVPAI4CS8e0dQBr7TgADI5rdhYM4Bj7fhI9I/pxSGaiQ5AfoD2YKBGvDtp9sW6PDMFrPXBF
2axwtz28oEFLSCmGNvPsl1OGnjQaO2YKwcvaP7fjorgk31l1v1XrVlOVzTUZ3Fq8rxXxxnrtDr9T
uJ8IqO/jolwbHbA5e7L95IKY69K9i1MwaSFfOeOXry75V+w4Eh67z9I23f/SGhCelXF6jA5thBuN
VSTs7pA0HHFNmDRXrnuEopSOKgol0l8NHp4xY9WQKM8dTmqDLuHV038OjuAegRLywd3SR+30mQ5f
9OczbpgWqPT+4N8o/+7/89AqjxDfYnV/ZtcnodQ2IQp4MHBCr/907PW9xeKE8F2YSs0NX+aHeqrU
twSMz0CMIS4Fg9yLRcPPuzhzPJ51mXRjIWWP8UMFfTAiYHMoBm8ZG4Z2drRVxozePK/qrb85rUIW
kzArN6sHTir/WyAUadwXovX5yeljd0WwcluRDrXmaYW4VXlzm22+yYsMMkKGvHeP+7xLy/EOVnhR
WfCjAJiilvtX9cB2fCosALRZA9gLJL3o9z0IuCbbjRgK4ytbHTCSPZ1qGVktzeAS9gD6bkhbYq6F
K+9oWBWcac5tx5ECb5pWOKMxnT0cVTlQtc9hbLjMJa3W+5xn5eWcwkIQkzGWQd0lbTHDlBMaFAzR
P8lJ3UE6WE1KxbUDyhDLQk26y2q3x/vUi2h1svgZ2ToiE2gGPfmPemvA5Ta/ewW/REBYlii6gnCb
USW5dHiBa1We6ZuiNydiiqSZ6+SYy9IXs24+tl46eH2hbMMG/KzUTbq7hAgaMven0i57ohTUDZnO
IeEsWa3PTvRvs7NpSMqTe8lXdR7lwzf8wXYqFBKw2R6KxPJj+4VK4Ipnx5wh52GQXk0sBTvZgSVq
2DyFtRzKZvs18NpoaGreeVoJSVwU8hVcRGy7YRciciPHNHKWO408gD7tDnjUlVrWdzW/nNx9S8RY
L33sfiZQyyMjf6A/WbOywAwSh1yxMt4ROcoeu1plnYJNPN37cgU1df6OaqPGJ2tikBVH4jTZWfr4
KJHWFb/omnv1Lj3/nrHLOoJXhknE97DDKRpyXeu4HUuZcSq0FXZ/vcy5KsH5S+y7KQ5GQMCSpNay
I6hMyH63nygSD2RlUWXIe6J9KBwzvYOTpeckIAyMGEvexNZaYbXbpO4eenAaOGRQuQddCRk1opCp
KECk2iitMyJfail1HxC+jPc+P11Zue9yNY3NGiWQzTEGov1Alg/3En4AFBvNivN7dIMSItaqqRgZ
lz44QytqvXVfotiasPDPWHc6/upgpY6PP4S+03LnUZQP2ZJ9PHKiC6/FdQKc0FkznzYTKHsHgvjg
JGffcWbEMX7eiWoZdBUY05EIl6yybf8lkwXhMFkqZqbUygGKag6AHRpFdkK9OaqZqDlAyBxC03Sb
53aqJWeK/0f5+W+Od1cRv0KXZjtHEP0D6hhcMY17Q97a5VjEY6v4T6JaNqZ65m7w1NfDbK+hnjnl
D61j7Jt2Xr0oU5Gq0BIsDupAKohz0QjIF8kWtWJARNSbXYQhV499Ii5pFo38so1OO/Vd2LhRqsUi
ViD/dgzpFXiAxtJzMZ8HNvx7HQPGSltMUiowYfP5Z7VT42AwvRMfajCGjr8JZmiXYpcUt6lmRJk6
EPUlHx34zT4jqLO+97EXjWSO+hWOdEerd9puXTBmCYgsPSejPyjn/ZJve1LHunX5pXJeSt/tq/8E
nTrH2VT+Lx9yvB5GuL7ScdN9+Hilw3FnET9FkHhuY7YPPNolJ9ksuVmJSBc4QTXeE0epi+VTcxz/
hG2HeSTFvO7ysFDketdxp9lfhuu0ASRHKntU4N02gDpVpbzduh/9fpNoV0EZwcWtsjE+fWHcJOyD
fMVBhYOlBdBIx2eA+cMaOyw5htLJUP3w1PxqhLj+8d3Ph2umSmm1wpH58mlljI67JMDcw1Q1zmEy
QLt5CuxRB2arMm8sG3/nivMprI4aa42ZR7yFDGATSAO8YVZXg/Zsn93n/J4QPOyErBQDKE3DGaVX
STFtOSQJfKPzW+MUeBQlwr1j+nvmZv/cVehUm90QYs8zx2hDM5UgLg8EzfxHkGYuQ+Nk+eKkQ/vH
l/95NnPMOoi8O1dzqAE1wxjzPttXINJu36SE50XkiiqBqTypJHxKIxtRBdyhZ8X84feencVcbTG1
Vfe5Qkou/UAqWtS8WQr0zEJhaK9r4NZ12eeL+LJq55mOjCFiqX/iUVRE77LxS6Q/mGf4Emf2XW2o
fQh9kaDH/Ljch71XEfNCXWUQbEAd5zmsg5j22HHhlFXymJINq/Htzc79vBHUhkAnitgNzSl4KeaN
cC+uZWkWtzeyvTS0P0a909v0ZmUt6xj+iJY3oCiMmsVcs5MLvKbYizhBImmffZm39vsUq1ytLU77
y8FHDgU6ljdaql6IQX9Flho3m7+vRyHdyxm+fh4gUDqIByuLSk9vMNQqPZIM6d45mKU3bZVZxdWY
VYYMNJQfaE+NLEqQVGGXuFK6azgIoKKpZEKXr0AoAHD+GmIutfqfTomaciRa44lsAB5cUAkbX6qe
RrnZY93wV6epivZacwnnklCS7GmvRLD+siwvCrALyHNggt6CQx06bRD7Fv2/5Y8pcTFMUPbpKV8L
+6cXLLG6c422m6FvnnBSz+DEtT0KqVCxl0P5VQONokaj2pvxYSMNr4ec0dfyEHUX6S5Y8MgPbuKx
hiR/YKOgU+9R1ZpsfpW29JgWzxvLxn/gDe0eaJEZLPGf1bHK0yRcd1PO0x5BBJFuy8nmmavW2DBx
pefKvOuqRqpFN5h1jovK9O0Ii6CGkUOyfpfCzK9dSlQP0R091yp1lkb15GKo+TN3NFxOnJ4aLLYy
83D9O1czJt+OJnj638z1gcz185KJ2RbVi7Us6osZdnZtEiuuL7Fa0UH9PalUgdRpADNVvz0aMtW7
pzRhHlbnConr1x0e3S228kIL2w3OUxqaoA18GYWhY9BY0M5d4XRM2v/3PaJqu0AH4KLK2jhA/KYG
FMbvOF1Lkf86lBzVtAVQf6skEirMhHr/9RXgMkdE9LcU981iOG2Y19/uYW8AW6sXxCBWJcXTUUbj
2WbsSofi0qC5lJ15YuE+B5k9bJoe2TxJnUQMjS0cZpZAEmirwIPOQ0DucoHKtCtzMQ25FpXHU2R4
ktv/y9VQh7bNDTrr0I+/lSgR+lDBivxCG6oGbgZBhkH03wL5cdHZ0n4Fp2VqVduKAq0Xnwr1Q0qc
i0wRtpIqANfC/Rm2wyQshQ8bbLbxvab3bL3DUJjcG2go4S0xtJxBfDB4hOlCKO0E91UfA3AZLhro
M3uwXFatr/csK/N2CVU1blpjxvGo8anRNDYywL98Qqv0vwS9ePYASTKVXQpBw5mEbsJNC+/ujBLV
F1tg+cYCdGiGHGVC2cWRMG1mMS+tur7Rsvz9SiMuPdF55Fu4qrt1pua+Ypb/QAniBy+XQWXv0OMN
K0ysN0PwLqEkbMnHULfrB4wdvqhbb71alO273QH0DtpYVay3tyh65rUOccP8hegdspSjHU5pEYuN
Ult/0Po4MycCXU/yjCTApnXChJTe3WiIe2swGfrPa0kHGWLvjCOy8uOZ6VAy+6BHmyORIcNBLvGo
CPwIxRjGdCv2Dkr1xoEKDR5REpYE7N3iGa9qHIxquzULjEV1jCtU04+NLhqL6yy5rfXODcWx8zBK
5Puu/5su7mZB5J+QELTi6XnDz4gL/+SIvEGolkhw5DhcdZI4I5XerYoFgNfLIWKvP9JVE9a7xnxP
G5G2pyHdFmv6g9MNKFx+Bn8ddqqha/7B3g7FFPhaWhgK8ThBx/XHRvGieGVh+VXcLmgLRoq/sPej
PPYegUpB2yZg5olDZCePqXGWw0Sg0RsePmoCQN9a3+REA+17jCWlbr40xRrP6LWyo9O5UH4gLiM+
FGUDoj4LiFjH1/yc7H2Gu+/Tm2/Ri9566CYF8sZBIzLd/KDhD97syWAdkCMyoSq879Dpma8ZXHO2
f4wuzjuWvZorMOv8rOnC+otxbUf5QPk+wojK2Ow9qBIZk1+bN02tUEt3xIukxxLPNiWsF0PRCAAO
RK1Pep/Ju1csRnVLuI47xJFSohdVKmMn6C5gunYwpfDcOJSvI5fw6TBogMEZfaRRsj/fhAw5tRas
2gnLZu8Lp5wNU3Mx4g7el1EO/5cMI3PbSVugjQnndS2K5LxOgnwZZS9g3eppxk8lilTkMZzse5TC
pqDFFfLyagHJ6Y2yGHp6tjXPndVO9rST6zaK8sBQPhThDC66IVnz7jo6xra7ZDoSNC6qTwViNrVd
ScBrSAB1E7CXnsoSMbRvDqXMid3o9jAOxwimG97DYz+toQiSUk1+skH6PdtbEes8b0JjE5lnZJAt
iBJBcVxnsWPB4I/ySA59hXpnaKyUqjVCK33xD0He4iUz7k9mnSD1ZzhYhqKddq3+Lyo5ir7riyxp
LXvaIzpFwrvVDAzhgWPwSvnKSAhJpmaYYG5jC13ap6RA44schkA5T5chxNpwLj+RE/zWAaJBtZun
tmMZo7V6J1MWrCRnYT1aQYQtWTohkYXbz4rXthCxWf4L/y1IRGoCQbqOBr1mb2Kwcgcca6gN2MVQ
SwQ3ZbxxeSf8BO5N/qGb5v99F2c164ZKs5UoPIEJRCbM5uiwp8N2OnrWPjjPGC4S7kx7OPMmRbgp
jv52T3DCZEoG+iN7iiOV+l+RvxqLhjy+f2Qiv4ZSv4RiV37iEhL84NgwZ5Qc9Vnsd513MGwLwBOz
8EJUI/zRbzuzoDwRDK19KcDCnPIxuqxiliZgfwHj015em4HJntw9iJZQfVh/gv75r+/rZ8JPnmJb
4XQNd1i2YfMVhyL/TPk+aeoaOn2FERxVSJsZYqrrMyWVWr7fcPLuWdOkmCnHDgdEvwjkTj7yzded
v2u9GoYoVeWv+FHWrA7muqKEsPmSNvC2FWU1fQIK46cOfB2+gKyEmTqS/cnnHMwGNFdINQnL984R
u81Tu78o1XcVGIHa2VxHpdWhsW36R41pi1ISUnSXBjuycaiL2X4U4XQn+HcWHqb/e8cWV2aXvp69
FwYHUFkJG9teeWPCTDKB042lx+Rf1i+grdpR4E959M2nY1x+2fbUpPVWtJ2kUsxJU/ataYLzkIlp
gXjFo4hxcBlBRGJhHGq1IglV33SqMf0RAxkJa39P+BV2x2SP0/5qilOoGYE+EkV1V6s6KK2JMvr5
lZXjLxXWvmMD6abw6UPd/MGjyhbEtiTX9BDfQbCQOQ6R0fcbWG23N4HxDbP/4eSLNA0/vmHbDPOm
oZIxRUqit6L6ntgfCMtPz/50rgKaKOzbjEJpGTsaJvAFA9AIq8qWrcvT4kyExZjJXl6ZjPBuMwXW
bP7HeOOJBS/xK5Pzel1t+nJvF27FXqi4VdtH26MLRZ9KzEZ/Y5FtYUWsSB0R6zqEgcdX8wrzJK5t
C81bSBn8DIioUGD4kX0vwFbT6txrl6J7WghnO47237yW0TlTxhFv7UDZDV9Xkh4HDRLBSSqSmqfD
IfxroG2Xb/Dsme7wiFJVXItOTp7TG1+AoAkO3KNqL2CDym3PAy6P4gbQ4w2GvY+hwXCAFWXl7FBV
thETq0esFOz9JrCKNINezJB5N8u/vI3xHilTtyw3q/u97e4o16QQ5U7LpO6b84uETjbJA5zBNJDU
e64D2UOvsKkUP8V0Z58dU30RQoibAQStpYXjDDw/HAV1T/KCOVFjcpGepLAzi0t/Llo+SNZZ5sIk
930jyh+aDy29nmFARETVuAe5j8HjItfts/dNf4ZKTsL5IFLWnGg3b6DfV1RRtAQqvOegVWGaoTnQ
z2wlLs6hM1F8/y6XKQhLKJQMJ4T1tL4dng2RBu75wBr1WjN/wwXNvYysFa8JPoyBHLAPo6mgJT73
X2TRlvAv8QAFEhAqvxpuzS1eDkCj+pbn4m+mytL/NvJVr6q87prtzQMj/sAGt0oBOhyJ6dsm5nXI
nULQOp2/ghMSteftOtXaR2R6f0HgXZC6odzkHUZj5AlwavaL45wMIW9Bl5tQsH675aT7QvS1TQG+
jX790/XepsxQjGW/ru3VQWtNpBtgfgaGv1YkrpAIcXsi7wmDU3k5FaWXiUhApskLFTrIgFzeQAcQ
w3IMFvXakFt4QOu3gLkDj5uGbuGrFff24JfH8iim8UJbgYEV+gGkUBWsDrrQ+yTQR86D2QtZ1DZE
djzaXkfGLGYa74k4O2lpCiZXt9p+l9845jdQcjdR5pL+eKyxZBOEwEsWGTZqKHtDXlu9+nY8/L+w
mH8DxrMNUsku+bhz9qQoYSZOqKAmbNTAsIJ/lqp6z4zp2zvcH6GDOpIpZ3uFZs/5K4YolmYO8xAg
JxDXWQzdJboBjmlMYjDSmCJT5+QYQbnE8fyZWui7Y9Ppi3P6V2ToWHnLGHWx3ZWCtVjelxifyS8I
stC35pZO1uDU+rYBgiXcWEkZTt1+p3B3oqo2QLMDmIdMI5qR4woCWOxzSRyfCMdOJZoENy/MvP55
AYH9y+LGcJsTXnaxuz42d/UeGcsacSx96T6gcjQjRPdpL12a0Zd+/Z4Ra23ktjDuq93Oe+iOB3qw
hqxkvn8LIfxOtpLOwpT3aqIcU7mVwrr614d1/7WawMkvPL6cxVQin3RZvWRXGpr5R45Q/PQGc+0y
mDgMSeAIA7F67tmpJzbVQc6QElvZKC35O6/q7FeCsU7i79znVh2/intKQGzLS61FoXWsHAOyBlzB
uR3H7wZvF0cEq5kuWYeLMSqWo0jdQB1yPuByUMeIQSd0a7WfhmvIpqyRb1hhsMCQ+uHWtVqlQpD5
KQblFs+Sun1rXdHmb1RCRR7Hh+JynQOu8/uGekuwefw+FjdSEdD5mRvXIPIoBBSGEvlmN1OmUSpY
glsq5e1A5yzvLLOnlWKJ9yylRUtn3d4Dde9o3Yaon5riZ21PK8NdXIYhRIMwdnb/vfogtrV0GfHD
n+TSeHL+welL1JP5dpNDayRqoPhYgwmXVEN33GqHAuZSISEgkGIIIfrh2z4itzLD+V9TV42iCHR2
XxSMByxA6B7JWxkQtpSdbTVbzbsbZhtY8CO4wCzHBgbXJJDgyKEnESeeblWGRD1zWtbG451/+pmR
inOyIP+6HdAaY5ZJ3RvnCa4Vwqfx9qoM2dKp9Dlux+RLmleW/Ba7W7uHPf1QHrvvfKh21FZGnWUV
lQingnt1R0W6EfWhul6B1vVi8cnb+QuYIqj+/cZ+1TNYH+kufV/9yZ55B98fNyEJgk3ue7DpWPcy
rQcS0zxDOCuqPQQ8cxBtGt0yh8vAoOdJYPlkd9BrXdB/1IRdC2zzNDQpsI8RNM6hyR0KeZAcGnZy
bgvl7G/0J9Y/9Cpdz0sH2S1gXO88TPEXOXkoV44DFmAym/ir74S7rplUneXdQzCsN/CVx2HGDURR
CzNLVP/bfXz/GcRwGgXnJdF/HBdJeAC8cJ3+LXdrRudiq0tR6R69ZcmQ0kmcABTpXNBCjOJWBSeB
hRbcXFe8Zy7mQnN6VIlhJm2ldz8zM968PBLkV/a/JFIcmLrdLnohcQ4VFImZkQEa5EETrkIjY8Dc
L4fDM1WkdVw/CEiqq1YmgFqm4ztZMXxGtlyGzDnkU4ffVvMWL1+buw3aQQYmSp3cEIHNZildAe/C
FjxUT8xLoGTNR+4dNgtTIyrWQwQ6Gu0Sbm0iMilHOgDhf6AFuvDA+t82MK8VxEKw0mDm/xePLxWm
x4UsvgiTSHWKHd1P0I9PcN7V04eMa9zf4b/t8FPtruBhTyhXjX8eUXvHH/Qduu4KBg1itaIlSPQ1
JCJxeDOhhGmJBgmQKvJnZPCMzz5Iu119fVrmFXrnXg4cOAKzFCnLV5EFLDioWdv96lwHDgdzVKH3
HmSJpV1JHJnoIcR3ZbxUzQnX8gfYDVtlNCNzx5BAEC7O4cCHUe4IGAMm6337g8kO+wJXvXxTzCST
pAvt/U5X/6kjA2rFGTosThMOECg/p/pHSVCa7mW8GuIbc60k0hM1l+mQrByq9rkV4f1VeyF9rKrT
KptYK3gQUJrnagE8In+/e/VRhgUsusBLxFyyTLqUE9C9qmO2D7WXkPVt61jXERdMCEuyeoPVV12j
wNQF/9Vax7njJ7wttj8Je2X6KoNJV9EjdCayVhWfxuD6V6SOOj6lKRQC8kBW9W4SF/uaBgRRqRlS
CTSmEt2mRa06/1I2SmrXyZ/laifkAw0RKX6WZGlq2qGRXwYP72UyeuPRkIm+g0JKX5igh4PihjkC
Vcek5+F8JYRgumBjgTt3qlYNR5ESaMbmatkqQalmP5cSwy0ehs1p1PV0hVfZE5g1ODQzfy1foHtw
rzAuSzS7XUg0l5CRjChZZD0CTfOz8jRAQWL9yoddNjDeQWkn/3a0SZ1kladNQ2ELyRj6BP3MAtoz
MiBfCuXLHwMJI8Gb9Atjk9YcsLGIown3EgfcKo2bUPa6pUdEnxORDj5bh2606A2AhTmCr5gmpZXI
1BqH+eV3eRqztHzbyLP2aPfbJwIg0z5n/rtJjH0zB8t4A7IT+IzkGlMHA61bg+pJUCZv8TlPP1Gn
N4zZysYdHDrTb7oIdka0C+hRs+BZiTRpVOywfiAbHtKEkaIFNcYEKfNFcjPzU4s85MumtvuZ/S0m
FJDdVHyoQdvn+Q/2YvpqNhIhzzwf7LpbnDVQr9bno6Vu5CDzvvNTQq7B/5VWZ44O0QsB9aQUPFQp
Kb6mCGH9tY7hhJzVBsocBQczydSNWPoTt3OxZf+znPEMESCXPTtrZlBZqLso9ybJm20K6VPyJwQT
yLHIrb5TETsjrRTfxsKBOrtFpBU6y5EeVnIfK9YH6XHakw/0r04VQaYwWiJ07nFacImT8+fiI2rx
dNRX13jI2xlMTn/FldbSzF3cWPEYlS799b6HW05jCeFmbgEd87MQl771VYvHUgmCrC8Oui6qk3kk
HJDhX6XsAX+51nzKafVg8ZpZhIof4cpz8Nj9BoLgCQYMcpeJnB83WCNEDqIr3ib0XR4OA9anxMC9
ySSlStd9v3ul8RrYOZDc8Dd+Rj684YS59uNNlsiVQmkbGJ9Zx5FRPwwQAwAOkGo5HU2HGZ4YOTns
jKgnEpkpVc2IZLx5goaVqXSJJzwNPSTX24P5Qwllw4xrIxApSDjadCEthRg78hdQfYWDWcS/UMr9
cg95lJFSl3RCV5dBORpAeXg6blPsfWL4tzFvIyCc9GqhPtWypi7Y293AVrZCX2cXyjRMBJxZW/U/
B1SBKnyNuCCstElW3qE/JL059q9Ri19Qn2TSukQh3DnDf9CBv8gyNfeBZhpnLIdEPZY5qSS8xzaJ
dBKtF+t+lf6EPJUdlWZBlBx3Hmn+ulcvX6TXJMmSAUDRNKKSXt7o9iJ7mUbBmyanGTLSY/uoNiRC
ziCo0I0WZXuXVwawQzBDK7NI1cRHnlCHaAOEhvXhI9jchFI5rMAu7T4DgCCx2eZ1huSnxEhA3cxs
fA6kwBYBf9EeOKT7yMelQOw5a0g3R7BR44gK9PUTdBxDxpKVkauDQysetcuXlnncbXYzTPjcfwRk
EBXeSeWf27h2/vwkKsEJE94gooDKkl5XePAztAVggqPJnSYaT+SgbhxeJ7bPFiF6rvAEa4xY2tEP
HvlgNe60J4Y72t0eDZCq4RLnOUuU2qGSxaafoczKl+/z+aMDhzuOAkyebSqh9ffdy+hPyqWQySwk
RBQp/pvS89W1YlBM1h1Srd0/ghno+VEqSdaShHkD7mZCjaZIpR+X9MscmxXj9fmG2rD1Alxyqbqk
CJ5BlSRsfiKCXw2PWwZJMe01/a4Ug9tVnJS2ya1JRDQwZ+8C27wQhX5W/42QUzLOK1s5w0guSs/5
7Q5dg0a8uffBV6XwmBwj1cU7q12vTeiq4ZoaV7xDqweD6oDPyZvz0SYuW+iuZDX5vbYYd4BqoNef
klNNIPXbTNopuvxwXoXhGaTbsTwdNuAv/eIkrFT3i6WHRMVOjqpQTHkzRU1iXxIiDGcL1nhlcklC
nrBETiqzE+ARw8exrMJZ9Gx2vg4tSwmrZgCaps6zVpH7ecGukCQucZFTmeCHJHedHbemEy0D2jwI
N9CHJrk259ehZZGHlcGynGi1leZbCcEBRCdk/rwPYrkFw9z1YZ00qlIC8bYFJlPUirossaMwH8dj
CmhTs1wE2GMeN6dHDDFEdXuSu8PyZ9cgAXRhTIny8Zb8NNY59TMdiOGE/mdVMs7lCiK71CD5DNRC
WmGspsb/xkvx+rHI/hl6muzA7f5LAfJeSi0gyc1VPbi0eFPRhVgb2egLDiJEMBl40CvyFty+6nGG
9lNjMjRMO0FhuDGtiiLyDTopd6+b8rRwXTZEcRNH+VcYL9eAXSQZZhkM9FdGwGjl8SMnA5tYg/p5
K4D+EZR5d6OQVXJYn4F5e4NUKdiU6w38yQBRCpVtNvOS2g7l5w5Anpz9RU1bbQsB0Hr6D9Nb4P6N
ZEm4rOISguTf65uYibrEC+kXUJReVYXWJKcN1o0/ahju0v6aau7LPiF+g6VF1hx6TQ2z+zASqhPw
HUz/RpcsfJgZrpy6AOWfrdSonrvi0ZJfu7NMcwtooXN77joq+WArscYSYQsZd6WXhWPVsgqXm6co
Ta7/cfUyKn1+k/n0V+d9rbaGJ+f780cUYM8Ul7hoyXV+gRH+PWRdToSnWf++B/FlYJJMh7QBf4cI
HNbMMUxDvyscoE/u2C/jcWzYbR1Tm1Ja9RRd4+/FeTTfxJ2Z8TpD2IfCbF+s4wnQZsrDz9NWOZXS
GiXZ9K7Prxd8T3JiH0dIEXEM+5Y/wEN1eP+ZnGIr0sEcr0eV06/Ts6RMwK4IAvWotdiB5xzv2et+
FCvKS2FzlXJf0ZZJnXUGVfTUHA8716JNThGMEgEt2np9WqafBCoJWuMs8aVWg/RF4hwH/GD1vPWW
hNild5LBBDy7yRI20TyQPALeKtNBqwER1vdBfIbM25244tdKNhIFCEFzFerIxRpQA6VuluYt+qUJ
7fGqMKUa5i0avWRiDk5kGOa2VT2MGvfTiNemRbFPI3S2YuFWyaIkeJ2FNcc09HKRPHqEESEyB9Po
fidXWt62xk3ZTIZUOlmau3Bphn2lNdksr2XQVZj1aKSRPXGJMSGUI4uEL6HEJxuUInxUtEkj95P4
Ocx92HhCpIJrJHUDGfX08nRZBz1mDNIKyCAlryxcQoRubAg0PzzU6XnToMSbTmLn1xuxhmiJmE8O
mCnguocvFsDkD3dk0ZSpYgtJmAlE5Ms9EVz7Uq6koEfD0lq67m0Zn+oeurzy/ZpLZFZaNVbF48i3
fHSyBQveCI5BssiPIF9FbI97mvS18WSvQYZ7+Epuo0tTUYa94ZZLgTBTTcFyCIpvbjU1/hO9Ix9f
Gf0O+trMqHuLb2MRawIkNYz6fLy0/Ei7NcQkXwiHWbCvrTpPEC3wuLN7vybqb4e+RQ5J4LJPjA3r
wvg+KusQd1ivUD8seTNcIK3QVb/ueZClce5I/xRdFKhE2bS3/UCNIpkMlhMHIMXm2vM5AZ2ug0jM
sHQE1/lOxjyr3sLc6BuyHmoR/IFgxJIApkwERP/rvuPnlGzXS07oHFiwVyGntHDDWRMvfNEV7Nkm
inW5Fzv/D4QZifBjvhA61/DSV0jy5x3IZJGU5HpYnrd21oRckI2zThysP2BevW3jkB7cz41/ojV3
U+FZ+4YEgfbRKMcCPRewJlXLGvi1ieSByDjLaHtsRGnAGvBvgD6e6YjzF9Ad0t2U/qUWQICLBPDO
QLNzxohRioXQgVOzpbS5Y82FGn5i5QHDZrc4NcO2cNQLXskcui4d+oeHXOntITy9PpVti2XLSXbN
TCHN0PUP33NNOlFLTbTvS0DqdIG1x1dBNFa4CzE6JOUqULiHZ7UEzX2y1V1yuyF1cycfLrE8yVgZ
8umMZVROQ79xmsedb1q4udQRsanzag7juaZ8sxdMT+7JJ70s2WtAXopmSi+WE3S4I7cxiIcFCJQp
Cao6PatqbvuGn+DLBryQoAiPJC6tzJ7muCxVzL9H3U52GzQV73wSbgU3tVRAO0xZ3Kyeh3E2fPFB
WwYKSAx7io+8/k467j2fbHTSaBBxrAhtK6HDkij+pWx5HDd21GOBF5tnenc4tuG4A2yGSJ48pkGX
JWbWeMouI1tcWYQaFz6KvizVe7yh+2m4xGUFIJcxgaYphInETHlj8p1n6BDN9Z77qBrhXkF9Z/0W
wlDkjiriM+dZQADZxnGc28uejdKMbWbO3xdIC6RxFGQtrzB4W0MJc0Uo+N3QawrdQp0cgIO3CL1Z
1fyrG65BmuwFSDdfAItKQK4gIdRgd/MKSh1xss5WsgD+MnCwVpYz84gp+YyKZvudbpxmXH6RPPIg
TxGvUZ/jZKnbqY8wS971m3s4w62z3oUYVvwdXAJp9RtjVtm5dT26+KdE9ljJ3bZ8RWmFXT/AYH5i
KQuDdog32Y8IrGOQsPZZRtZ+cyTUU/kmUCRbGsVCQorDinwhLDg6tlkYmCNzHhwE6/wc2PTgHf4z
T/HUEyPPBSTapaFAVNY1lWbUu+NBLalwEsexkbkOJXnxCQbAUQTwqs7UE00Zbmn+zwHVNOhFCRkD
TXQwa7wcBkJGc4KNrDO1CynoyYS5Cowrxcb2F/irkmFWFgZIRUFikJp5e2CuNqyYr4RZ322AP0RU
IcgKVhEFONufLrnuy+SwgL8g4Y/5HfiA15TJF7Rd+3hzVVDH4SMehdkFVElq2fQIwwRivnhGLvMG
CWDcK4fGV543OQjkr11OsExE1u+30RAwQ0Ll1fe1lRkvpcDtrILDEdpDtnfUxIxdQ4qbiDuXai0l
xEX67AyjtQzFw3iLHfKeqFvS2V3yncDOzDJa68oXeSrPEy/tWEDn4qE/NUb5wMuR8RoE+JCASamD
gQEhO3Vj3aXTKaTbTybG5x0EQq//Ixl4Fx07k6eB+gpLNXElqGcAI3Q1jLKHtJJswNoJk6fxYjup
tXi12ZJUhMCCb2/hGeuiBpXPW3UljBZqHDBxsKvlgE1SomSvEFx3lw9OypW/+byxUs0UDJUFWSoX
GujmLiNTWdvQY/cfdMYL72u3f4IoLbq5fzRft/+q34zrK34IfeZrxM/3p52+EM0kryKPgAlWK+Cd
BgGDk/sMsUMgEgrknJAcXitlTG1eHwSZB2NziJsRT4z6WhXHP0wZSiMdh4i73u6X0Ue8v7muJ+EN
0LOfNoAZM2TX/nfc3xKGXvbcbhbNBWReCxerF9N+tEYByxQS94VJoQbjypIjtsl+o7IEqJpg5J6X
9IqWHapq7a/KAabVR7z4APx/+aU3tgO5N5Y/5C0+icXR6xLqIxl9rnfKn+ewXxcavq7a4BUrkM5G
9rJcqq9B5m1qKE2R8eTbzV8j72mMZrTparvxwnaNN7g6MUILELyfkZRyLseoJdlz0Lj266ZMMp9T
f/wwvn8WmgcLio/AbkyIAvDq8QZDHIlwPEIc+Xp+U78lq4DC9auqJQkkFAEM51KKCz3fygnxEIBV
RRjHNsvWThRxZVJ5tIxP361ZaZnAXHuRVDojmfAEh5WMr0hkjRHU+hXUHtandbkeIcTmn7qeXQvn
uOJmG9c+AMY3WHXwoi/Alyv6HFLlQeKEbzeEGuuACSiNsNmWINLIFWkT2IkJynT2MsD/PiVT5ah0
ic5uVSny5jw+87rLfVGQ3vKL6cyPTlEX0EC5f0QU3sEjgRsWcXF/LfFAP0UVK4Fgu6pU41q7IcfZ
vpRRI9p5fEu0HERc9ci01PYdqE1CRJFUulxmF0qUShAQyDFY1Tabck/p3xCfGs183CyhlV88HGGC
31fDsWQyIOaFrPe+TSXwETeIGsJq935bsHUNBn70ae9Rp7sSrWdknGughgI8PKRe2XfhqRjzznHj
ciBqACrUh53FQNSZTigEK3gMElfDQ4imPDPW00fT7+FCCAZIMupYwpItDTE/EVtpko1MQe0nDFka
tzqSIwKadFioIHOUOs37j9xsnT24/f6S6WdYRFr1neaSe6FNifTkSi+gbkGY21G6ngT6R+Us7QJO
vUhannKFC/DzPwNYMMLHc3OJl/ypa+R6arNc9E8QZf26uQqdEKjeMYTqMLyY40++s05Wu1X+nrvT
DzQBk+jBdVept4SKDz8sOzBw8ZyhtyRMytxr5/yISEEUJze8rqe/DYUAOgjoFGChqtPjNSyhYyZO
ddgO87xD6LA1YO3xLLqeDR3tveZ/kCYiAKpHwjn7a1DkHo9H0k9zC6lwQVT/eZBW6emhKZqBsleU
FB1T5IC4bFHzY6Z6X0a1/ASa6apbJSK8W3x6JOEGaKK3CmlFQ603FS8xz/Dx8Sg71Vd3gnUxMRm3
fqVTs5R5plf4DVe4Hia+k2/9+ZWhzvpmPr/WrpY/7vCwyy9iYvvVC+oO8Xtc0BDF96ixeHY5bi+L
8dlLK/Xk6syEB+v1zRJkXUhSusxpIvJT+psRBrn6j6U/jDTgO43vmllwGZM+KuszrcKJOrkwXuiR
yhPJI8HYUHLtmq1LbuslkNyr0PuiJu/E8TDJI/x1TPMiTczu7Bsw2MiTfzCMuvo1S1HPnrGBIydM
ZGG37CI/2G1FmIaHcxUy1jaJ8gAlUGh1hGTwZkxuj0gCjqk0AYnP+k42hnlfGtDAel1sA80PdaCg
M4EeT25qPL1aWbBKsBJMMpzTgvspJrwYVyuWhyv6SdPPgQsgENjjtaj/cCvFvp26aWrMKB2b56AW
4uM7GpbMihIi3GdB8DVOSmmXgGd83LDlcK6m6NYaEpCdoN4xfAiKZ13luPtcEGwRVxyct6JmI3FM
0q6qrMkkB9j/QibLFaZGA9/eIi1dy+Y3vZhAuApznXALyFlZYVgNBFm3Ug3Uq3UQxPXuH74V4kEB
jzRRN75Z0eIHFbF5YJTqMSaBQrE4NEIcvqeH+CuV4kSpVrtq5CIqYcdrOKKr4tF1J8rRkH0PZC+b
dxkRL7XKVmvoDtoq81x1qV4QVm9iwP3+hGjEET7Ooa9gz556N0xNcm8aYqiNBbhDEMbfEShz4s+C
vFsb0DuTAnhoRKmo24JOlN4o7yh1z7K4DFzk8qL6F9ki4WgbIkEhN6MY6pDNTbH4/bcghYZOgpO0
xn6dy88S9rlzYW9vVWcQIkGctJDP8e8ZgZbAwDQcD7pdK0RxycooKBrcGmWN2DliBTYgT1uuFdKf
sq4i4JNo8brf2BSUEMLAK7kXy+c4NMkCZnCGnX7zrY7O1hP5INhBFOHbGr7edu1B71nnihebGpkt
OhU+XQPcu421boDGG4206kTHobEqwPnAXsuTzr6AL2tH3TPbZfgKAjxIjY6W1nqP0MZXqOWKqnOo
QOA2lz3/NOlQXDfjOnRhGenC+Ed8UU+UiJvh83484BNnF6t0sIQnMZMbY4y3PY/nojnLU9rfa0k8
aHQGXGS+BK4yxIiFmTK6Q15T8vHs0N3ERVR65dnNJ/hk+Z7ln/th13KdR27t6KSsKM2nO0XZeTTx
JP128rcB/D4vesSFUnaq6ndKI8pfTwbFdpyGhsnppfVTKp5kcD0Mjr7SfXXW0q5uVI9JKKvoCVEi
C4YIl/HzTTOVQn1JuhOWtGS/hbuUuqXtAYyBY0rckO5SK/NEayLdp33Tkp4iM+oq5DpAx/hwFJg9
QIaUrvto656rNcPO1oAurpmG6BmtL4v+kyPMXvs/ROtvwMSvXpkPQxHj+o4yoC2poapxqr7Vj2NI
F5bypG9D9IKDI+0P1l2RzI1PdGhNW+9OZqFzy9+gtXTvs/RnmjBY8fNXM8j6UaYbswFu+QkIrLA9
U4STFXq9Lot5FGhmJey3bg+/UfcDOxF5Z+0bWfUff7liJzVf0OEeZzvL4JkECHhl2QgIJLxrsiFK
Z36k1BiXa3tdP6EEIedB5Q/nHiX5zSKoLoFMvCzq/K1iIWAh+aO8cZAcJQqgfreVu3nFgMF6iLQz
fvJS5e7NU5rR7uypsqloncbeBY5Y7NALtwMSA/4Un9xsjDhb6yCENcpAaIWnpQks5OEzJBoc0dLu
4zB70R6VVe38t6qzH+QNoolIxnlZBNzSC4O6FjRe3K08oX57DmOZXPWw92zxnLChNKZWRSCDjMkz
ZWaqeMfJucWbHf/4U4+ozFFaVjGvgts/zqjWqBQClEbEWjl4DopMdkONJmOAugh7d1eGqTawwuRd
LBQ5jPknztzcoGGs36TFafsNNX/9cJ9o4AD7DrwysjTGEVg6KPNDMNM7HhMBUpsSeWkFNKu16TiO
7syeSlYF6kUvMzXIrNqoH0aFlCRpKvslcwADj9IOp3SeQvBMrVqyxOGdgH90zg2ipzPS76z2PA85
r91Kuo904+XEbByTkg4tQD1U+XaU7RvhXSNJr0YeCCskaXROIa0xs6wVWLUMZ3krBonOgw+dsFpD
pCfLyfnGVMkfHAVDn3gBpJWFyBznr1LDoW5JL5hf7oRO3QkJyoYwmgxJ0N3bTZ2iUr2bUsxApQVH
jJ1mOWfxG4VjkVhJZdkaITuolmRFryj6xuttsQHJ72eh0Ot1YaonY4l0sHnYaaEeGqsAw08dx/4U
LRzOXiqi+cn5USt75MDX72Un/up0UP5O+BApha0xvBQ/kAbyHlHtHpJ+9FcpezDpFzgRUNbWgrzp
W0oYurI6zqv1efKVzPKml1srZnEC+mpko+/9ku32+v2ufcaqdQVTyF2k8u/vJyQS0ZE1jZ7FLrDZ
wd1k6qCDYDXG2qKdT692p1bEhbcdSuB9NuBRtqZHkcgRBw5luV2dpitYaYUfU5s3OngxWUj1GRCh
JCskEaANoqEy7rUxnc6yfZvYvFqGKKAcJ7Mpf4DE85lxHRtUVz3LVNwXPPhoFG0GWdWquKuYBV2y
BTPzbxYXu7Mim1HAZ9c/D1+pb8EhZiaBUQlEno1TT4+vmf8Fxt+RbtashM+2tJjLlu2HFOE34cHo
VVE8nWLPipVTvD5peHyt/MJM7AfhL8mRipS7eNPyjS3goLz/+xWo5PAnPtAl7iUZF/w8j3MPHU5q
uykVWJ5ltxkyMcnKT/+MnulnSo9kY200gzHqxPTpMMtef2f+iGAPijNo5PpK37x1AUcou3r25fkF
EjumZU9BqQDgOcF/8deBJA2NEYhE77W1h8Wa11ueE7qlJkSny0bOrAjjhllzvtL991EWpvXPb1sH
KikLpcehSgk8AGepnwMx4KbNy0QTjjbmlJF6lryGNrNmxLHVV80ZWayv8KtbmkRdZqMyjs95Krs+
hTGc/z+xmJGR05KKEKzU6Y8MmWh6MoqgKlutRxhRpB+LJlc5VH6au4m5NKtl9XY4okwxyRekuejP
G3CBBvQ6VVQ1/2+B9bkfUWaa01x9hOyHFXhhlfe3x/r7cS1TxP1ylyg0YsvcVRCZnFe3UP38bTTY
UW0XKuvisEcvW56Zg99LZ9GhxDUvfQKEHuzsqBVbOeG3CIj7euObYcBNp6MRNXKpl0NJ+c6pPtRJ
Jr8GSZgnCgWAVzkADlqIC64FrYvYDDF4w6Aur3xdrTQG1+5PNDgLHqEY06s0iCRihMi5wuVDBypP
zY07kaw/jilQV1dT04Ws9ZT46+2cjhUKWFh1h6Kwe1udyodtj+N/1/eXk9hBfk+DWdPjL/XsNya2
EAHtqRrzp5byHV5i/8AJXr69J5gmmz9nn2f+5lgrnOTk0ns+ym3N0IW8vMZOGP4jqvDrSZ46T4vq
gFcZXsddlHsHdaUkAD0EDVbJvo+DjK5ejLSS+ZXI3WCNS0k9uqQFRWs9aCdC4q2KgC0yaFSRje9b
rOQtDLLs7Rxb1K4sWKCmE6vG9vKcA4VmB+wTXxP0m+Hcv1GOp8Na8iFXcWBcCXVR2o0MamPAXRRf
MozZq4kFZLCdszwaUADKHxfZnb+4hGuFyGs12UnaQRegUNiToAYGbJFJrWuygegVot/N4dgEh5kE
W8HK9ssZuumLVraNKDWLTPVo9iMEPuuFjALi3Xs6Ogj63i28TsdmnQCjhNYTGz0KUCIl2GrRpSD8
d6KHcJcSAVUt2015LT6A/mkJFHHLLEtQXsbOIcjOiSZUWw0fnVu4rAEnF5y4+S/1Etzg4C8gUpMQ
+Bnl7RykTFAOF4cdXop5SODk/Q1uolZytjbQXTHYkFuO1YjF4DUhTAYZ2OUGn7B1//k3/98tJRkL
L1hPpXZaMIuBEHb1yJBjyIAByjooSu6HSlJjYd2TlqKPzl9aRt97VpMfcP4PAY6RbXmGfgu0kCYx
sN4yP3DHAunK8X9FlMs1sGOPX2CwhAfznKoD+n5UI1hIcUxaxORARcoD6cz9HqhOIRVnSgp8C3qK
2PlgYhS7Uolxlpm6Gf1noBHoaw6odYMrDadTPh2ciqo7h7HBdQVYGakeqFzHckQW5HuSZgEhlIqI
gXFTZe09/VmL+KDc1S3CCWfegxkSPl0NBchOtVMqoET4yMv9Z0xYLN1OnCysufDf2uhlkVs6ohUR
EAH7/HLn8C9ksBQS+sSLV3FKaXSbcnnEtOEFm7l8VDP/66uyDefVL53sutjvXvIF86SwPaxeBM5Q
Ul5C3URTzr/DhWrHuQZ5N9VpM60kmXQBlszmaTDl6P2eE9DPuO9OTUEo98aLmKR5wUWBVODh0GHn
Ay6Y3ui3eDDKvX8NlBiMcqKfTU29E4goHqP1F3dhkMjTqoBpox985ZLYHIkSgHoaUTLCMuGBz65d
EydodZ8Ca/iYWsCzO01DjsUhNMQRpeaZuI9obCswG18uNOz35wzMlwKCYqbhXgXByixlnwTNTY6D
ndoO8og4Ht5tB2AlqjPSsOd5ICvq0WIsVJAj6zcdI9CyK2IocoYm9rERL0PhPxbgOWn6cOTwrotx
QfCS4rlqWe0UGULPAToh0Ky/MicivpLN97gx1uyvDH1d3OJM0921nKmDwyVlRRhBMv/x+6po8poF
XBnTCTl5pLANhyo5MzIt139B5gmGMrrUMnHsUg4Mn65SM4CYyM+KKHq77iDozdji0gAftjtYpnYy
6s5OiyP+pFS9ycsc3UqrzfisRYzZrFswf8whIDJaBTSiSeEXzcKJgwNaCXyeLgZxPsBMIM2tPQZ8
OdwlLcE6G2yIDzdTzVHxq3IrEdEZG+Zd+CZu/u6q8w19DK9PLnSd4ETRoV+CM0QMICKTN3e71cXB
rGPDS8qoIfmr/eDINT81bCzDZCPbi8EXYLFJR4sINBojt53NZwpnOs1CBimk3+40q2yxWbUW2MJd
cQB07q+2rcjcgw3Bf0zoYQ0WEke6JF7dlOUSiNbKMkbRwTB6rIxCyCkyPxcR6zbVCcoMgkyjJH/K
XaDi+CZZfr0R7HKfrRerKciTmWXnxc2oskY+myxQc7BqMwqWCzqgOShw/ON5z5NxHfXrY94DMZpL
OmlywQTWLZW8wjUGqp0xo0UOoFItE+ymJHgM2ABFelgb14eOSUuAbxGw0pBJ4JwnTrSUnraPWL3r
aNT4yhmrBDrnapQXcN0NvZS/MNh8NnzuAG4qEQd14NvDNzbsd/SjAtbL/QrXXhk1tGbsBGJwinx7
ukLiIvlmZ2niV4UCZrfAf0SpGh94R+2IvbGIeA1FKZlDx5nhX+L6exq9bR7FyCrMpZTsusigrhox
pMj3U49C/RT9DRqRfZB3ISa3RV5nJnVB/l57bqZlMkaw6uLjFtjXp5fQi6KTpsyq5zfXDdd4geYW
En1NRUst6a6qZwtFLHn8ZXHN8B96GxJH3ywrULK01TLgFp6326O4pkRdooVmJJxnLNh/QZz9Z5vE
T8KdjU5AqOs3JfA6ZRBNJbBktI0qaolcYVHMg93lRxPoGlS/FOcXQXlOA7mzsQmh8++sJ57HcYFN
M6PgD+wWJtV8vsb45TvXZ3flQ/9Ew6WOCaCAmfiuzZp57c+EFmsehI2N4FBo6dS3S7WmFWfwCZz1
CVbxpFwOwtdSQH73lddbk6atRCxST2JzUAwWiJHT2f/bOg/+xQOmj3HdXZ6LLY8YBcwPWWT+42bd
nF5X8ThwVAyVmX+LP+HlqvIZjbG9twlGiiJNC0zowc2nag7jkWYGd0PPPsyGzwA8gQaOttIOmiRC
fiNUJDJElQm6QQ+SroNaEO8swk35yDiNfnZ9oj+n4oiPfZCmywyeQPrJeRsYERore6p4wQcKEMFI
AubryVOzNRBE3SUrXsZajCRPgqDunNoij2q6B6xh0bg4WHGZBuxkylAExeDvSf8RTpNVi+jDrAhw
kbLrAY+kds3YZGbzswIj4S9F0LTKwe5MDsU5gLR4keILdNHGsKYitXTSAtKeqoRtt/tROh7EhtqO
FJYc8V+e4+X8pyPJQ1pLRU5rgB74B5RYpqGUpjMROsddONlC6jjEygFShGL3SZWGh1JNcw4qWp7K
flJ7431h4csp5tkPHkNNlQL/YgaW09wQNymOfsEncCbFwWrvNwc+flYNHqB5qFqayEmAttHWEh9I
oMRAI+FQH4DiHrEmyI3MWWd9/ic+AZSWYYhJWn8zNxLMPlNhaWe3vWYss6kqfvKMUMBcVPJr2/jG
Ly9sJi1RNuo1yjP0OBtJlv4RYO58rcxiT696fchfeqxkLNIHJ//gXhnDoKUk44Lr7q8xSA7jvlP1
NQhIz00n8Nms8PZPi2DpcESH71k2UK/AMHh3vg/2cb58jvbAVUg2CG9RivkBlQVhXZLt6lOWM132
sQJBTWrCkq10wMxmN9K6XvwLwKYaHe20fXKkIJQYrt/ddGSLwn1I9VkvGvqassjcdEsDbEQLNBGA
o5lNt8NAoHfgbgkse/pfjufWCOMFmj22wJhp57Yr8h4sBRIMJU02pH7QuZIQOWE1gA4d1ZXxdGPs
K7EgLkVD7Ox8iyq4814AcEj+qqeMhdfNbbmVCb2hXkeW2EhwGDYAA6qUFSpcop6T9paAHfLYIH9l
C93tpJFAnGITpehibkqfHqdZR6x3dXrxmzQMe2qgkuvAB2Sp098jG23j37K7yYJ/nEps5YgQvb6r
PtmceNazHMMaACyriSDrjRgVlUuPOvw1sCy5uwk8YaOM2B6ROJ+uJtW8vnQGeixPzGaDWs45nvH6
BwpH2VQUZVN2Byn6nQAXn3PprMdSNcG3k3wILBZjzhBCWPkp/IUsGlJoO6My+KlEfBMqfBoNbpZs
JKDoLo49pjGFUS8yi1d5tZnFpXZNcITK2RwwGaHdwU8IPCzV88j4FZ3HyMgXFGhAnNp8Iii9onaH
DnMfwn8EO8WcgeDXYiAuC+ztpvj32SWWyBJf1Ogltwh8ADB3ntYlhh1qDUOe9+9yPwC4GK/iD6NB
Ln3LztW1wOfHlXBUqOyOSPYfHliNId8AF41YhxWEBlBreB+jM+R2d+GL+f2xXr785+LV7AXk/k2v
dDjrt4B3Wx6vii8gkfFKqf0Ji8Z0i1B1gFjvzTj+P7VfqSIT74djrSvqUaYDzaDelMOAQiRTrcRZ
loMqZiX2jqzsdhLRw3yYfDM22jLiyOPVPyiRx2XeXZTg3onZhV4KNrM6U/akm77+HpaHcmX8/24q
a4ZYjDISzJWRaIgWTRpjWCktaxT+DlV0+dmDbbmgm7bbN5d+LfdenbBw7mTqBcRIVXWrdwJUjsQT
67CJJrzXlcrCTVL43y8yjTxETGvsEjYIgzmMX17aT6tEZ8RNbJW0RZ6GF3WXas+XNGKrHAspGdAY
64c0WEB/5Dd+jeLpXDcjRCXvCwfGg1VPqk+Fa1r8q81QFGk5l4amymk3t4xBZHGRPyQ94odJs6wY
PvNdTh/oqsUVVZGwleK0yVv/ssYhMh1Nn9Vi9PVS2LwuPP6YfEG1KRer3vZqh2I1KpNiI7Rb4I1a
j7rDw7dzLuzvDH1pixHKnEC/Z5GDQGTO/HHunuL3qp+Lcn8dYY5tder8CCX6WbJA2xFQZZ7Nhbe8
01oW6IIyHH7pV6nclHBhNU4DcTBmg+gcQQZb/FiugKUQ9sI9O2tIoKPWFAmxkmKufI759IVPgHB1
JrP1YXMhGcuuHfv2LmB8BZzT917LbJDVkMySUIta1Cl0w2z2XpxpVtLyPBNMdBWa8xa1NSVUQtD2
uAxDsWXPGqd8GpqRo1iQL5d0XpGFUzgPW4nM8GGAZHLPXoUzLhpwVnConQYw7KxyEsIoxpCav3UN
mjrBLCN+xMyEd9fbQFiWeKoF9a0f2rST63iAvkIy+35blBPStx9iMZ6lPvPP26saFYb52vN3zDe1
Yqr1cKKbNEKwmVPQpj4epprouPy0TKeHThbIfPIPtcIRRLyPXx692TD35cro7IKJ+ItPFjwKAfCk
g+oCtsTHxlt3+FTpkDeAL/KFKToCs2ZbS0oxilqA5E7a3hpofg/LDIDIeA7O1/OXI6ZkbB0UYzTN
2j6DwUITNCiKtbM07EXrVoanoYcnGu/RJT3kXY0jy1tX6HeSz/qr5q5N5c2LpUkO+K019eiVYz7S
+oIEsVqSdammzOdOTgwPLftQiikN4sjgw1nys6NiTUpw6ysuBIK9TCnUsbbfcD2hpVPdW9hVWCeN
mCPt4Rfzu5ZgqacGMJwd+aXS2VsQ9/hO9zJdPipLra3nfTiSDwtPjnyzaWKQHYkHWLX9HcJH6QJo
Ckd9pW7jCXLDDc6zvY2J5OFfLnLH9QaVPpttq0DNSisKkcSiCEVKf7BwY4c5jIt3+AWqiwzcOd98
O1dda0f/hdHpXC22RlmJ0Y1GH90ZjZ1Gy809nNkjzaLfDKep0xXaEA6MBEdgvvx0nRWaOedYjMUP
kYqHeEiBSkW5Lh9fjbunbZqaN0fepdNdEwPg1smEoCjqqCzHIJ/TMsR7822RruHiveoBqqv4Tohk
LY8zM2a7pLXLRkKgPNOvBm2N1xUVJZVFYp34FeLma5D9TvcrfkRWi9RKJfew0mCnDl1DKHSwccNj
gPnd93M8t/pXDR5/NZOaCjEVMLd9IAF657ryNH2gLdASZ40xvND5RzSsI89jhtfmaPM8A4wHTCJv
L/csNfmqH3W7LOoJkYbF99L6Ubc1ydZd9SwdA50azBowx3duDNfvToXrArSvzd05L8yolR3pkR02
mOOwlu7SVqzj19jH5ZFvMqesWa1K1QjTtbd5WDn6puJV1BB+hXvhStpK1tV+j7PnA7huuTEmsPzE
AedsoSNQZ4y8yQdhBgtnTjoqWcwxLjvXckN4KwMgR8eLZzhPU5V3tpEWggzxXxSc9hlcqNdxVm/J
hYHxuLUY3th6GzjwO949zXeq8J1R5ukFVw90USes7AqM9ENuamcuy++3LGt//EfP4pawJKZmTdCY
7xTElbmftDv3ZVKyaMQMaIXU9tajNNIH3AmneGFx9OWAIFWxPofZ7rVKYcKkQ/bpvl/oufvRCVBp
KUM8BtZiWDZd/Bpp4T7NWWESMzs2EsQiHlu3ILe7DmcX4AFWh9D6xxt0LkDR9T/Y+F4cabcZVVT1
LAagkjG3Jn67Ncyf4xV6yBeQ/FL1tLHQzw+3Y5ctEDxtycLKzkEHBXErl4t6SISU6i8UEdkXj1mg
uqHaIqG2OEPJnNG7C1MaTH+hJXTj+ywr5qyiV1a4VUe2YXKjl7+DI5+QvRTj6/U7BRxFqWtDYT8s
vUQ7YUklxntnfIaUUSQW4I9sPTwjbshMRbvfdyBArQp3lHWvO4DyPBcUZCjXNdQzOmJa+gf3fimt
h5jeJLfuJFW253fKnHAKAHgkBiAulCKBZbRkgM2MYjXDc2MHCDKX9+TaVULvsrj7ZDlEZ58KLlOO
TO7P1ki3Kq8UTV9DZISBPackAnKEVWKQs57HoqMeUl/9H9igi5r6Gm8rO8oNt58xUegWg6WH6LrH
HtQFEvDL1xYowbtTYl5Ck6bV0AjW10seMxtxzrLJyLSmHQUA8DjrRw4VqfwCUgMObCpvDzrotuNB
ZEPGvZQ0MCoFf3YbZBZUJzoVrsh945ne189mb4dj9M3WEqZBHmV9bMBmmWhEZVB9GdeFsedIlgv1
JBcaIkcef45mtGFCG0WtjOP4qYUnObQZztZ/Sb7T+TjJ5vU3dX6ZWjEyFTdo+kbLE7FoaOyg/g6c
frnHTyBDGh7dJgiKCx7/aAwaVloLVvltGvgUyGGji71c6Uy9P3L9wB8vjGNHEgvN59fX8uBm+dEp
vU5KqnocnRD7qNCY0KK+qI39tw+TifaI49mjcLD3CcQ2FHk1+X6NkyRmyYZSAD3ibNRr+E8xY4ZL
e6hLBGvny7STIFL7iYg5QBA6sKPQjG7DfmNLNmwftSEEVCcqLnBU0BozuUwiKOhCUhalgey+Nmbk
Gm+6oMDLJeqQx/7h7z12csJXeoTMQiSCNyN5612RIsh/oeata/eyL8CBnLqhUCeWzQ+2pRzBoSC3
+vhbBIrmco38SREEOb3KQMCKsu3mZg+mmzuM+U7fZFphiIUVEe5zJIKqWTqdf8JuQy+LuYraluCt
e/wr4XfmVhjp54Hy+e9jkz89ikVk9SnT1XXoXlqbUoRuTFuG+zcxM1hDQoI8QJDGxUzGMdYWvMh7
lupcaGOr6/UcsQFjePzcG1zGLRR3SdSxlnevWvW42EBMNj9bKSEkcQNGj4wEmTTw0Tl4A3Z6Ze3v
1TQ0qmNsRa1ADTtdcKJykBAHaWiETssazGM+YgsZ8PZuSo9zSdSG+s55wQs2Cyy7fjBXy1vsYRI+
o2raEug2CtXFzpNDbRDi3OTuvgnRL5+ZImMasxiFKOhm/+LSAE9hRXbQ8AkP6w5bsXjeyfBf/Fu5
2KuW3mXArZhwDRGb8TnC8KhBUuZJ5Frsc4nY6XIqSXyxU5fNHeyNjR9fKUjdWdRiV6bicBw6pEWa
5//xke7yeWz/2uy96Pq6kfvSDs8XZxtehtudNu884pvbaN4oXspNKKTsNs0drf2tuRtIrUAlNEwO
cLctG3FtkTZHpo9BP4xfnHePNVBdvDzHVZdnLi+zNUF99OBbj/O9NKOze7T6+GI6dxc/Q+2I0EFW
PZUvXAOWIHkngC7e1l0y8Glbc7bkpxEZMnXEiYrgntqNOnGUcv8XGoHlZaKcJkl3z51SHzc6NNuZ
T25Rd6g9LAUoDakujjOmC8+eJ5ZvzJBBlm/WWzlmrewsJ6ub1w7Ir3SRcDEFMFCDLXakESKTjqMe
HnHNMur79wSCNAApFkKepPl2imBBNc0gDgw8DpD3XwwP3otc2k/0Z3hO1YVgOQjaUlQEJ7Rqjp+w
cnEShGkmR5E+x9/AhNTsSCzTZz6YldRwOsKBMXQ5BFWhXcb6XsQxtl0BngUqjjFv+LOaRD/hEO/G
rTZaenjx5w6o3DtJBL1JUKP/QXuAcMcv03/Tis4XaIq4B0bpRqvodLkLFnX5eAFTOIx+FEoObsCn
wACp63wRzgo0u0QdHU8W1/bzzDykFnOAjlzIzZ1A6etfWvZZQ6uwjjZ/VSH290FMOCCSPJt1WfE9
4JPd02C1H0cyhIk5pQUz9z8b4nPzhgd9P9QsPh6RLHqt4PBvXIqFsnSpVLWZrzKG2RgBPNQcmnzL
P5jGyeHZk6aGcXMf1Tvnb4U9n5JIRdmC5E/OTjeIwc0LQgQLr+tMf4C6vmCQxVellOGofZWE8zOv
0p+TygUVlAm6Fuo5Q0KA1/4YETmPMSHitfeWxYreQKBztlVL+CAgKfLZ2D4sOkMBH85oakQYr1zT
MNxUXCASBq9QXPTRTXc7Yf8fstF+NJPOu35iezXYXOBXvkpcyYHXwbanNmIPqx8p1HHcrKQg9I5W
AwZq/+oGBPZV1A/UNcjIZicgZXs2Q/BCLUyE0zHmbBcsGk/3M9gLkMSkzR4oMxEJq0xLa67fDLkx
Tx8tD172wBnWGrTzHtWp+u6UidAd+cLHNNc4KRWu+3n7yHwLLXo78i3O+Mm33yaojB5HrmKl0Te9
o6w4ZM5SbiuZdhmdBVdZXHrcnYUOVhSAC4BTtxmLqm0wC+h5yOavpxR0EGGdOKePToHitH+/8L3O
Y2Gm9p0IXxpVHTnmllf7bO9/91ovOnDx7o025j4KFW/GMsWIacCYYAEhE8A09J3MPGe97mkC3VCp
wVXvY81KIuL+AuZtwNdKZi39+R2XfVgTPkjxgpbWb72HXaqhyb91FO5q1f5dMfqq6g+V7VzUeFYU
59QfSlHsAjpn3Ykjh4bwHwIylMRj2D/45YqnA88YzC5nyFWt+vnHXH88rZhbZ/eIk91H7UNgDFD2
Qc0XJXRjCFhBSjaJyF8XP2Q0+GucK7tDRO0rxabdL5GSNI6hDjAzARhKGRt76Tl1VhqnbRhhs9Lk
opyuyuL7kWW2oOEvZZ0Gz7cpZITG4q+xsPa7L+KOzxnpdHWKbSsrGVaWVwep3sbHvYyFUV2+Daf5
CnvwFxuwssMXT8JBBDKMRTPigN9+12CGGs2Ns9r2Rfk55gb92h5RsXafx63oH1kKHzX723lt0AK7
hhiBJlPGB0l1La4T773Gea4dcfPirQbY5H2iqwNbb+r0XPRdRd1zVsyiMOCXIyRK2Y2n912riFbH
w+3UnJWeP7beBnuM39j6PzpRoKV14U3NVRlWIHfpvY0FVArAESM2wkrIuIJbQRUeMn2NKlPWZJwM
a+2jV3dQ+ayNIbCIOAWFPPxNWY+Mdh/cXdRnMqxJY3XM2+j3W0pDipoYXWRbTjuOWfWSQEsRoPR/
VuqdJA/46NDM479t+4r05HN1HiiQwrC7zPIxbixxh4AptasyGRk8PtRCbiDNhfPLAbuSszQW/faq
drL53omUH0Ovry9kvMalF8EfJy/X3hXRMifZ894VeRX/JBLP8OQzm9DFLD9FEikQitqfStGZAH3j
bK3P0vTof4fl6GDi9gyO5NDXPW+TTEOciChnBwHoTh7CAGbQrBQwUy2CrE7x3iWPs1NjZdqFh7oL
dy5kL/eV03TVB1NN4S0C4RT8s91NvMalAFeQzx3v183cTFFdd65Pv8h1i80dTIlERuuqvDxFciuW
e7jkkYqjsqcdatE4Rbf7pzbcOAQa9DGNJLa/EJqDBS7c/+cvl1mSBcFoJ8DQnFOUqLnlqTq2WKlo
OL929usNiADU0BUxu9IAF5mQAIya5dRHY0POccHwcTn7jiB4rVi4ALzL98caJK79v5wSnGutI/iq
hyEHw1J+alCzY84phCH2BUq1awyOxNF5INVVZstG6Vx/dwlWz/pP5WSJwbN49i5ZzET8K2SQOl8t
xXZrb+2TgbVhwTFjUr3EP1UjKiPmCeiXX4zShrZmmA96wc3aMMS2GuLxRwzO3V1oI+qwZQoQ6H68
WytfPFIK1i5R8grh7tvruk9AJ8RAf0nZ9VB5PGJHArFNITGX9giq5LoL2/7XyjRAW0AhxIsbfdOx
UShVwvVDkweRTBwRWNt9nGNUwFqh1n8WXKLFIjZAdCew8odG3qSNGiddCS3am74LvfcvpNAEPTE4
mCCJB9ID0km17oFZkXgxEsCS7NrwOefd430oSDPe6czg8hgFuGaB3ZAf2wUYxd2FFSFo74iwQpU9
/znAzkaqKklMjWBiUa+uN0LjK8k9m3dh9ngOquPBSp/NlVGcZDkGOB3Sqp9DGa9LEPlE2pbRl3GW
CyXF5zr74Gjq6ji8uIwjkCX5A89IiqsTm3LAAIp4V3HnzuL3psi4DOXypN4wj+6rbZUmCybCgjvO
0gsiAOpfkK5loF6amc7wJvnN+rmqz+SmsXK3msEl7PodvilsNgq5C4fSDZQWNptCv24dVrkkUNXG
CHE2rIuBkeRJWMNDSKekQkRFTtlp0rMRz1lgf8kwJLYuEgSuo0Sw2TYwM4E1j3SxKmCusURNBUcR
F2MmdbHDvzVdkSQV0YaErD1RrsJV2k1Ym5fk1YDvdEA+NhnUzPukOh9W01XICDm1qVW9NFOAAl9m
XuqKNz0PDmMgOCZNutUS/Gl2S0LdRWB2cViZPtfu6EuXeELV8qUFw5v3j4J/vY+xpaIIGmKhnqS2
HjOgDELjU0XyF8WNxQqZ68krNvBOJwo1oD+w0tT8huAc4rG4dP2yj5c5eo7+xQ8/2jZOC1goaqUS
Ihm+sFRTCmlgAXp3sfJnkdwPHLJXI9d27e+4GcAY6iqdp3U2SHmvrXLLHJt8yqhka5IPctwnNpj1
jaBK/kacXXJZCO0JhGa4pOwMOKbi8feJ/Zz5gsIgRLa9syQMmoTJKjtIR4LB6Fl3dTT7yOEvfEEv
VbkqiW6ppISmWBgqc45U/mJcL00vBSJpqBVJLf9m1wwvxoLB/LxxYdTHG5Hj7FpexmcyhhMJa5Ug
RQK371nCc+zMmEpJPnOxIByb+dWHQ88gaeoo2PnLWGk2+98y7SCQQqwQvp9pmZa4zs0edPQynd23
oAvIg4heesOkzt9QDFFwGB7ctouv07f+bm4bwosWS2VaD9gA/het/eV2v2L3vN1nv4iS+qs3LYgF
S8BDzJc+8enGI3L1TIai4CnQR9oBHbcYC+0eqTSAiI53/Ol/2s/aRuzxjBw5gYX7i2l57FSbJJAh
NL0fk6MS3a9AAf8yIa6b2+UHLXTYUIu2MPVWIbcyDW20g9jNXfPZxt7RAjO2+mvntrHInSRwKLIY
1TuABZ0i1pjxzLCuLUrKs7nmppiaNTKljeKxbmEhQwgHM2sj3wuSpAG5CiIfJlAQ+4KpnvKjNPjc
jRaO6IOwmHG1BsXCOFVhkkiLGpQXE/LsshH6ltTeiqc8zjwCKG/6ExSEfHDToqYOzBo8IeL1pgQX
C7kdLRAAA3AJ96EGAXe153HqUTwQNuQ4Jsv7UgEGZYuV6OIvYyMiN3yejLw+8nEiv2pcBYHCcbf5
TDugFiRevP/njQS7PnSgDwGePShUUNzkI04NdhNSla0Mm0JzpUnPXAPZNiD5/D+T6kVtjJmSNg/D
5pxykc2fFQbbrTg7m0rXRooI/tIdtTnEGKHBpiA5HwnBtv7L112AL2vFCr+BLuKJXGMCwXKSougX
nmAuSLbktkkRFGOGTdExrBzgvgux2f+CNZG6ktvJywDQEwZDgIPf3eZrdoR8VrPg5xoaGGf0CXFZ
yHvrgp7JedlMZ3deovCtlFiVofE3AHVm7eBv0ZzNC5i0L0SyeFPTc3a1NgOR2xPt/PYKWHU4z3eZ
4MEr6xTLNyD79zJKL2m4/mw2zJqugvCY8Kv2/G9vCa2Fzj81wNcQp1oyM8DuZ41fAdJhSEjjPVTZ
xCbwN+JFS6vlQooQVcjJWRkaTnTw9lybXZBOQusIuQk+j76NfjOjv1XfYIdzfqZoS4c7qyiVFeky
9AmZa9SsF/NlODzJeCjhqoI6ZPfJnbLiMX9Hw7BtPvT0SI1QzL0LgokbNagIyZo8ojTmdae/8avq
kZfk1J1puN5L6JO11rYs0RsWiLWQsH6YC0oALwMaemUil69Dj8mq0ageZr5zzW4hgoYwWfVwFl91
GUa+XaQsuolnuB0zflI05Z8OU90WbznKUxZtddtnAxMgAOkr/ePnY425LZ/D8BFfvsSZo1vwLykZ
yUy0CyIdxvEfAkbtyyI977AdCP0aK9xbQuTMzLEsZJSwwaR9j9FcwGVrerOrdgDRsifK4GNGhTtI
WBxiRgv3eJfMvPaoFNw95enIrLVmLFMtXKFc/VjZvLeyUI14fqntOQQlo8l4jc7U6GZ6v0CgNF+s
fXnGwIFDHNwO/IuYA9v9F1qOFdtnR9zM8W3hzdGnzobeGw2/BpVtArZcr984Jpb2udpG7F6Iqv9H
w7Ji5CpFH6ItuIyYoVXSNOhgpcZTthbPQ7mf6mqC0lvdfTqJdd0nC+HhKzEFCzmZIR8d8El3EzXW
CAeeNoImzrfU3uedsWjov/6lnRISgOJcT1iQ15WteK/8g7gYHoJ56sugchWuAuTZoy4GYLu6aVDX
hgmBvKR/CY6UwZvt4qvb5E8M3rXL+kVZ1yYisUQznp6B0PHy+uAWKLhbUwSmjgnUBfMnAMNDCmFp
XGifMtupM8+PuMXVGPJWkxvSElQVRvAtP7bnqtLltbSgq492gWQ8SU+R/6Qtj3Bb9vx3tUrFWuMk
06QfiYC5ttE0moFgXjH+koC9HT212L/j0R8mLm254fbG2/JyJ9h2ZpsCwYHiiLoJDIlBSfzq83aX
/vZOMNO8lysFO04cC04DbZ21Djq0uSm9aPJpKg+mer7f8CuM5TH5ameAAHFGYneEsqRT8Hqaqeml
uWMOvHb9WnnXS09n4d6AHH210g0b5+i83w3bk7NfVMGj9kQ+8opq0y74ucE/vLgBzu9C2eorsymI
Z17DaJ5sY06hmKhQJ0nUjqsvAN0VaCx15A4mq3RAPKejHiui5xuNz+T6Lv3/C6jgG9L7uBnl+Ni+
oeBQrh40nvChIybm6hCekKChsAN5jr7FzOLIoG36XRZGUXdC5nB/C1RYNxYeuQcxyjL57xiUXPVY
YvAL+xNa0i2CfRDBaFkYyFKqXECJDa3JcSOsbFPTuhwzSjnwGmci8o93wEjWa3JWXkwgbOB0b+C+
pVHbiM2J1uYpyw48TcA9QveULvPyJBHbMmT6KxdDDS4E7QmyI3s7Ddb3FTpwjgkg01ymeWb4IDNX
r6yZVZVBjKlKcWbDMS5q/w9q6Xw0Utnz+beL2lOXR/Q4gqC3hvWI5K2uAf4Cw7YJzUBIZUOZcaTQ
vSkvPz4TnRSDLKgrD52UvAyTvM5/KubWi0QJlhX1H4ZZf95JqWmdKAf8MGMKluldp1HD9x4qaRCV
mEJeeuVs0Qm9VDeujjvWdbh18rpl3NmLsB1hG9ryQj30ohlo3z5gSCLkGU7mHqHC+PDCskrpLlTW
qMYjef76icVs0Tu8DUw1LLw792kpC5W9aOXmLSo7IMhkBi8/EgrZOr5SH0FhXDaNWXtaFudneLor
I7UjIX33TGoLLbCAokgLflj1Pe2sTuUTdsb5xbEJhycXkTC9y6aDKjugFqVK5UcVBUZAq6AC/aZS
cYJPjxIBZvc7cBqV58R/MJjB1vw/0fp40QnI4oOrivOqMVR+0RntlS1mKXqQNRzg7s+SDIekOExT
vzrfzVaAImtExW/S4wh5Q8Qe+4EpX+Wq7Kas3/vVhAi8sAyK/KZuDPLPkFEj5HP4PLblaF0+xy9m
ladIHcxx9QD2LFf43NQkgnxn4Z8Lu5rHKZS9oNv/yuwn9j9Z92LEQYwBqpbupVfp9LEQKKjbM8j1
/hU/LWdoeii+4HuHVmOkqomTSWgPre94Lpr4ksTz+nreL6PC8zmHrvWF/VL1gWJ/KetZsMXeeUGt
NSg39vUqQ621i33+3mFQTAyui9hoRcno2VE23/5R7zaVa+jdhZxQDmnCxiIGLNXzRdKDzDCpIVlq
wKPtQq2WgLA2TgRoOjqUJZMY4gDTHFHy4XMdE2/EKWW3E487wWDamMEBRaCT8DFIUPMd1tqxqIj1
2oxvpnlovm6/ReNkdu8uXyTVrAADeIV5eAcgYybtaok3MCrbvrtSjHrK88h0OlhW2f8Ft/SlohYY
4V29z0wD/i9fxy02g35s//aNsmHfCZdPOZZdZ1pv2TLERpNu3hkEC8iJxiKzIdsUDMrYk2iiJnTY
wzRyqdT1G/LUUdJW6hWrbg0v+fvDCl/RyPKWRfYC1wBoDbda2Nrvg6hDV1SaunP17DNnLmRVChU8
bpBhrop5sV+O2GrAGJgHplVbKRtdcB01AepD1CK0pHhuYGMzxsnQTwM6JCnsSt1hQ4WmTn1RT48c
bjacw9a+Yte6ei+XI3JbkhZaxGcdA4M8HDq/pWb6C6rMU4U4av52vOEUOC2BVfL4tWYIDYKinVbI
GpK3T1xuxA+n2cEVK5S2dURYs8F3AUzO+6OK+5nwVO+3qTMnOSTYYky1ICrfca/4DZC3uTg16HeM
r7fj9jtfL2zO+Lxi8MCqwabrqNHT3d9Fa1wNLCmizCOpbI1RdGEe8yHXvjZOnaO+571sU2/Oovml
O5XetJY8/FS+ToFIAbrm3b5ywSyR9DtWwAk+81ndCTZNGn+5OuzkL6STrPyJlDBG0PRVLTlu8rzk
XC7JuGOnqjQVfnuDv9iSlmbyVLi08oR6BjoauoBFFX98DpkUQTlfxtrz9SBpRJ03PS4fH5g6sbo/
vYrt4ZbL45njwDmFap42T6m3OJ/VCfu2DIO3jPLkrq3VK+wJVSzwTF8GvgePDiU2ALYG1V8oPEgq
BDwAe76bIoGMECZspSbKsEobwaiiBBZEK6dvS7BkXL/EiCIngk2Cbk+dZqigDu4Wv9iZFMZt82+E
becc634mmFmyThUtXRGfhO0OjF4NMfgh79vSnSJOj08yWs6raUkZeiqBiLW6iLC9dc15rudpcVVF
/qUMHcHmaJKmSxFLbxzNPy9tojqWFW/3tOHI17LPzoJZt8QiZjN8YtXPdcGgE3ouidsHHe8oWvwk
8K/vu+UHkm4r5NOnGU1jGdvM41vRNhs1ebQGpVWbr9O0iRev6eSWvayXScUjFqpiQ40Vn5gsCXGS
2Ptwb2LT+zlDy7sY+mdW8pfrXMJC8dhHAOJ7mon3REF9GlJ7SF95R/qULZ2424XhnYb1ScHgiPuy
BDMJeXkqk95wrjK7a/ha+roqhgNlycPJ3vSXyS1/XjQ3rspe4twhz/ODt354TddzbLQFpRNCVY51
oTvfsoYlmqbly7curMbUrvYAc8HhbHcZwGB1Jqew4I4nbh2Xi2GUDQMXRfZJ1I0tslSKw5SKibUi
hr7l+KRCxSnuvGd+jgmKCMPB6W6xRQZmAijMlV3JAwWXa0drsWa5YFJxXcoOcky4UugdbdwB1mwe
ZQnvcjjNefEnKeVAruI5G5RBOEj1rX9Qef/qNzT6zfKRft2QZIzpETNbUQWhOoYIo6enOMpd7/Xh
ODI0EL40Rw0EtbGGgyulH746MHlcsZmPWq5EJ13kOYgeBYsU7RceZMr6mDDszjZK3ix6nM1Id8GC
MHY5YIf9ylRm0YubJj5SZ3wypAOJHzNdSVDBgBKrw780rjqRjNJFwzJIPx48btSVzfozsVyWnr84
WSSMMehllA3G0+cUSc/heghUiFBhmdPWob/mlCo9j/Jay2c7Qtcdq1cbewu0szPbIr7PWaF3vtub
XnPBTLdRvnHC1xXyN/ItDhXaPu4loCSAjy0gSt6wMKnRLzHzzrxTt6bhX2PEf/Z8A4UB+PDv8iGt
e0o8ihPLeBR5BxnY2yewpD7MjIbwj0xcqaxebO1NRDo1Ws1YBCz5wPGmyRGRTQexw6M85nMtzh4p
4DkTvEbIlevPjrigbMlfdwZZ3DoSrDqBOz60Pq62MAa4g7QjP1NUH5CEq4moykrunbjnJNOkT05J
Mm2p5wrslXtOhGQHC9GOGtae8zRIIc2oHWatpbSLRvr+hIZw6ibOALnkqLYy1boBNC7X2o/y28jH
kGXeVhSGa+ImhQeummwl12HQ5D5BnnYY0VJv0mRZ9XsMLPF+YkEUSGrWjFXXf14NoHN4DA0XAJ8Q
KWqyveZhsWkEp/krIu7heove+bhpWHNLjlAktkoOy/Vtn9H3GCUPgFWLMNPiR4hI/4BLawwRz+xG
B7/rC05fzVYGOXUQ4GD7AwBn0zcPyPWaFMoyzm3dmNHpV+K+WXgM8rVCr32jhAMw7WhAOMMPloq7
ruYi0Hk/Q2uFrbWxiZQTFdiYCAmOvDix94urm7z2/eE1LufhXuQ4FyoKRBG8r7bBtMmM5vDhgGU6
QWvPpNvgLPK8Yz85p/mWpI5dbyT+AOwkDjPQsKDSjZGBPALB/kSscxM4CN9Nl1Pw5kXdJHjhEPvN
H6i4J9mIzYd2SEzWekPTfL3mb9KACFCnJaZInsL5raRGCqAQ+D/NBnb3+G9P6H+t5T89G1izjYXC
AkWG/Eu17SbDvQ1l3gVmoSP7wu+st/KFE6SCy/dFqsNOu/SWyfMKOf7ZPqgfP9kh43cVmEzASmxg
fXfI/64z3vdvLHbTCArdY7P6eMXAba84aZNeAAax1LT2XXaDo/QRsZre+V8Z/xDIji99ez9h0OaC
qahd+vhL09XJuXjYNGqjKaKKfcyoSMSDgbJG5UXRknYl2+Cq3MiJAA4F4XBYrRSnuMoCkzQcg/tN
CsDCX/e2cKYGlgopd1b/puTVNs3vROVEs9logc1OGrAGSvrH/3Ys14U32tHhqvuCoNgbem53iQmu
m1HbKLSbUeowverPe6Izv3a+YQmSKS2+BRI6kTQVxIa5g3OMKKq+B6QkYqitYQTmiO7uFERoSMiQ
O9K/8JRn40r4F2Vz47bDYJHy5CmUBwNURR+QY3aAR+CJynKcQ0UrSjwstzSOyUQtjkC7f9Lya5mC
S6rPif3+HLkCEPBMoYiVDlPxFGSUFQ9C9c8/Ep42/JmqbODFn3OUm2rATfsAA13kzJ0jaAxtz5BL
wRN0LWydHyYxnEgKWDV46Ed7Mu0H+g7J4HqYktPINNloqHBkQ1Q8j7tAU144L34HI8XN5LVDBwkr
ZWHZcvXClfin2QvPhqslqMvvfQieAA3uANcwzMzJQfIvfCPaBYtT00c5zvzCC98RBimWqBEGMQZJ
m/ys67ihLirQ6vjH6Q9qsqKOR2r+gYaunopzDg50lH7SRrJEfmW3a3jpRJrn1O35j0oaR/4TDgFU
O3XGj6NxpuHLgeOrKBjeFQyNEtxHlEMTtRR9r3gGyfwry0rTkjgZSsWO/Iw/xBvAtF/wpxk9kS6o
+xRm97fFQ7uC2IEzvPCI2Ggn22DPRhriJcjQIBb4ZYv6zjlW09MavSoZJhzbqkm+O2/gNKuQZGPo
tx6S/N02xFfXQe348d9jea/8LWljcR78MlNBLA5NFThZkYjf3Ww6spkKfI04afR3skdGPbknhwOM
XAIf9h/GQJnNpjQ3j8lNaBTh+1gFBjKuqY1Vjtj1Iw4QT56W6eJeYkZVM+kDWoTQFQvMmQPGau+6
Q7hMkDoeSz3xOj4bqfog3e7EiVcMcD0iE3m38EZf7io0mSeYMBVs383QCV5KCY+M1ztI8fa3mp1x
Mm9a0jZHyGD9WtNNmredKDRcyWZ2Dp+2ishGHpjqJ6anjflsOG9eWrf0gQ+byw+UZvL30+ZFcaET
GEsX/4DbN9qEMs3mq6kRn8nygho0YU7+hiYdHRfvi1xWO2Ef15pQHw4oDSNfpc1bTCFY3292Bm8n
G0bSiIWfY0zjuMuPGr5oI+RUZxyoGsoLYLSOeVCQi+1MLz27VtexE93VqBh3QMJ0Jm9Y+aN8Ax4V
oJzs4CEnUvBr7KAIYACO4UEhuvlB8RgBoNgBCqipqwNxtl5sWH5p4VSE0Lth7PVjkOtEKVYtREH3
QwEJb1zcBT/Iu53BWeqt7kjFIPDe4y4fhgPR6rDH3erqX47nY14R/b+kytaFx+XxHZCohmGYvIMB
2SJaCyuM0zQtr7lz+Bbiy6Bu36puwKUoAAjw6ikuSc4LzB7vGOP5FpvOe/SswKVDM66YxqSZWxEh
AOU8W/DyHj9UjSW9Ezde1Pqj4h2rtfTfFhAm6oYtUilivXFXyILedplM+a9eQpoUl8ZW4BX+gR0A
t2DhcUML2p9q/vfe/xjGecAn9rYX1s1BqPxRvY+Xdw9klgz4lxoaw4dkO5dnsbeH9MQpUs5jcV2H
l3UsmhVK/Q88/Mb7buF8EDcoCH46Im1mAv9hQBMyXnuetvH2bc2S1a4b5DaqjMVwkQlZAx5wGQG5
NJzFlh0j6MhOo2EUqJOw+xD5cgZTH77SmzfJTYJ3nkKqzprGGVn/rYXYDit4QSINr2G95nRs3M9+
5IaurdbvKwz4UPE4Da7NvXdNv1xlAn/wYvlTZUFmLM8zW2WzcSOJhdGIklYFH8tM61785cSkzweS
pBsLnvQA1aovT44Vc/i5eLZRNAmjxcV9KzPgLIFANutOiSn20od48GINQVBvIhVpmO6UTy7g4yAt
zxEpN7R6JMbATrvB6dgSSqe5fvfEeiHDuENwrdcVhyHzZy1z2fWFa6aKlwfTkXIa65RRv3Y1AzQb
TLgjPirTSlcoLg0fx5GZhpaisIrUDrj0XseZOo6RH4DTU4IcDEGz+VYHeZ11w4hTU0EPy0mohYlk
+v5O5qcS4lqxl1d5oyDJqmsKihETIsSFbI2kfos/45X2/q1T1acOYO6qZMw64+msLFN+PAXWECnZ
fdswLsqrl3cKsZPW2soIrh5D1ZdQTgCrKWzzs9QrmvVN1fs5QpfgPrAD7UYVyeOCyGu0aVxUrtw9
U+H1RBan9tBupXIqQsIeEzP/9sabGZaT+EDWetuQpxhirEScDIO/ACz6D1TaUhXecMsd949TLnZ+
gh+vbQjjtF+a5WVkxfMI2WqGNHWC/vdnpIPlTOv0yRGSbL11F9M47KNIemsywuwB43yJqwOAGcVw
ajSMBf02vRVaQChQSlsQqr8TjuW/adnKOFO4w9U1P30KX/mGToLi/4tC/S2tyIyGkALbYbHeCJcl
P+HdlDwxVnkKsDKVbPLW3v4ehndxHW8GPBd2+xAvyOGlLZ5yjQND1+LRcc7LzWBo2Wnwe9Pz3/WB
l09FKeCeoSxW3rYDmArdPzSgB5Cc5PZzCi3EUEOyOq8l7JBfU3HU4zAcUFQYF5Ot66jwZXbVtCSS
Bbn4u49yrbSWHfNpOlQEWQHphw1lFpQx8Yb4X/ONBOilakIUhnbyXrPD00Uq6GM4RPNbD495w/77
6RtSidH7fz7czJf6yuAFOWmHGGOMQdSn2k7iPlq15ROMqntmvKrSU87rnsvbk1N3FkPOt0gHd03k
OM5Ri5Bk+xlN555DFMP87I0yrCeQidfSBEBd0uJitr0OEF4x+kfDZuYw4/wBtwvK7QMBEuxwBWBh
rj0YR51artGGBXm79GJqTa0MX3S38pjk8kQVk8vkzoatCbYr3xCzh2AnIZx3/S1KCdEfcrxfNtOy
0Fd0db8dsrvUDNSFdz1/43ssDRWhOrw1r70bQCv0Wqv4kFRZaqsZgLaNBg3QQ3Wt7AuDAsl7RW8N
JakxJieEFpcQFbfycP8nbkTQtIFRP6I9Awntwc+eVpqrH+CbcHxpBgwK+fPkL1GqaMtsDDb65Y/R
vkfEs1cMHe2wXUmxthnI7Tz946FnIqOC6UF6qwrPJzUNWx6aFME5U/BMR9cDypV6tFAHEDDVgbBK
4rXdQ4DbyN6XQIXomK1G3lHq3CMoa+DAMGQbSARXD5Ex2xcPlgVzcVS3/Ozx9rO2Tay6c93Op3Mj
UGb11cPaxbGXi14xPvLWN9uWJmp5os0Cz4PQyEAGE5b+yhaAImEBZE6bdXv4gGRMT9s4xNw2XKSo
CNePCviv0WBXyTmKLF1VgUVXCiLJCP0531+zgcUZNmQGi0h/ZDVYRTv57QCYXUqnDgzIIX2594RQ
Frw0dQYH+g7YfVNTM/Q5Au5LVfXYcv4DupijvDpACi3U7gffrJBOb6nAuPQLfRxQvrMWRdCWbmAw
/Dh0sd1WtNGEgaHepUqjrhig/JozwqtyCUH7wTi8DdhUR/S6w7SxJ4qpTuGfeDPV00bT8+yqs0Ec
qtVgCr/9FwwhytqdQME4zCPUqPQEoZY7YS5EKmjCAB6qmGcGXFqB2BSSRjIlTTFlsAjYBDslYLpx
7B+42x+xX1oA9V5z7La2h+YgcPyVdtlo4plR1zZYYoyIoYhpqQH95QE0gC7L+z+nRCftQiTbYVtf
5S4QOTFcwLnMg4G+qtwZlTQ/vgxl4Nde4m863drnVJFOdJSv3BG6LHaVxX29u/5hKKJAsU2R8dPr
p0J21X704KzIHQqbyXlCNhxwGTOW4iOP2woo7UmgQLTAz8DnvEzxNyTqbVMLtb0QUy5YxsSovg3r
/TTBWQToKG+0IL7RtxK7dRBIsXXTCfBeQhJYLc6z1TYHmjtEs3A66Ehi1VwKEOfPuRnoyJDjpp0M
tZxzIsqFCN/jZdf2BjDdv2KGfSY4Nh8l9a3tKDKh3mNZqmZFPLVyXCnM6fbskZRwRtos3KnoOhzw
pd6dAl1vcsjMJS0gpeia66sgNulPUDzXH/8pybdaZ/7vtTgtMC+sQnx+NKimng+UjDP8Pwom57zS
mKrmX0PVNUYwfY+0JjRpUiELmeVMUrZ8OPEy+7pBVhrMDtCcCzVN7Q6rjG6F2hcjz5Yp+qQhvoTb
IsHG2fhvTEInAer21+cM0CnIHx5M4Q3K97gN025HlVxiEdhOG8RMVkiQCEHno3Dp3DsZVWKFWeNH
iSVi/mZLVH1skm7DF5ZrYD3BkKL1dFEmRg5Id0mzBZ/id3wyIv6vU7DP2WZ86DM52ruOu2DgFycE
Z/iKxquA9AHW7AffQmFhmSWreR8IkMDkPW3bUw6TfypsVBCXZtun5+TrLhVnR9Bimqmdk/dR7U2+
e0vxvaWWrClAB640p1d+Hcmyup4Dzh2YaNfzRVSA1a80/UGlv4M7wJhDBrMgcoNLeJ3mJK3nW3cN
/HjNQmxYrS/SEjG4jTHpsTtbBP0Dr8s0wO8KM0fepZkffwdAXfFudssXIC7uvjfZUNTqA95O6wfe
gEXRUDlXA8+Dzqozek2mppFf5igeT7RpfQ/gievovBPVBTnJFGIuE1sZwzdj3CLaupy2ySc4pNYQ
ZuLfvrbNC4EBnAKg1/HHqjQEcvZAEJsEXsTaPIv4s57lDxC73sg8S/bSHHkAMSZ8LHmzMCyvyO3o
T+ghXj8yZy1abGbxmz3/VjaTaWG0ONloz65Youtf/nSIhvs3e5b1JgTfoawafifZKjCahIG4JLZx
6Z4fz/KYY1apr5mPYS325BIUrxe+FVpawoPSZ8GD11ZLHf6f+n5Grtq+FY3s5tUDqNEwzPr2U9Og
8bJVlkoSZyMyx3TWc/DhEsE8KThXiBBd8xXvVutwp8nQadb/surgxdk1pLImZ3XCbWhH89I/R90y
HQeJAwC8tEYrIFZaqWhGhaFsssSWC/r5pvCk3Alf7Lo5+HX35M+fmbZE8q5uriyA11TsiruVfFr0
vZef6RXwjHQVCf0YaZl93h9zFNmNCh+K27T5xPzsk+U28azWgaTEflkcVDYQ7/Fc9dlGsT/G6RGk
y4AUQkbyB955THZvrBDwmYw9KOqWVkAp4hK2OtiuRPn5d1VQy/0G7lfAGl874El2/V53gTyRrFAx
0uUZcrG9tj4Xv9NrBehELzDRms+KF0yV4JDENduNZWFkDTU8nocbJJ63LygkdQ9r/TJM5Tr2H1Df
JuaQAisJd4ERLTSTCJCVUL7FZOBXnefI273iMjePEUl0aoezptUXwBfu/KiRAwI1qThqnYqX5QVq
m02eWxCOLkvbQT+5IKqwe1fYudqcmHiDD+curjS+9IH1sMRa42xd9SXd7TjIN8XKgxL08A4woYTD
8t83UV31IHph4QB5mrDC/2uf6PLoUDrBDQZb5GUxfbyah6R7IVGKC0WShJCxs7yLevdOXcTDubbG
FBaEVvYhmBJKwHMm3+eBsfGgJF036XRW9QS/bRvEQO9uHQO9eamEWXtkh3q9Xrw2vw8LpBlt36U2
cXy2DUgx7LCamcZLnXc0Qt9mdike70MDAhlCGeOK4QE612Yq76EMmp5VrCxIGo7GNhs51CduxlAL
fV89jjCpIbcnMqXI3BrvSzU9qUtSpiWFre+hoAG3RrHREFOOmQ0EChWx2wVWek9aJyRN/TTd0vQZ
thzFabmsv3nwyZ/cBBC5jJZAYcCSY/raDSkKevn/2U0AbUXOuBBfGvZaDBe9u9ZxXnXh1PejhhcG
KHZkY/ELV2MCt7kCiGx6Cu6rdnxw9WAeWVm1IJYUYcXzXFYNZZ4GLWjHEPv8NYUcFmYfY+v6CyWX
6GE82xcEDeZ9sVteQmiPMP4RMFo5nmQPzgja69l6jMYpGW+bZS74dYKBekdSh2z96DaAcvcz1J/f
QbfGGvHw/JT/R71HaPY3whlUKdI+nFlWXVPL6sRaXdaXwj7MfDtb7rpQ0ppXGaJlzQDr98d6MjNQ
YrrriZTq4Rtb+kd7X+aAv6m2D6XCb4nYv5JYq9l7Q7RqvQ6PQAFzN5rhj8Hk5hFjZpI+RVsHGTZ8
Fst5MKHcVte3gFUGuE2zWp6GK+SwTwRkHu/awnEqmoTRI/t7nmgGVsyJOulcWneNVk8raXtaqIJk
eORC494kLe7QuXB9LKI48Xo3NGcESsCR9Qx+/ksmEYAL8pZ65Gke9ugzKbev72nUludlFjgsQlUM
oIcDvvLPrWQWipicyJv07Tp+qIrNv8H6nJmkVxkiKgHpSvHxHC8slsYX7zVDopSDf2cYp8ChVXfY
y3red2TncP5AlwWdWOnwRsk9btnb0c5Jri4CY3ZF+lo9I6Z+mSqD+fR9vhAC77NlXNWHI31dsXYk
BthJLmH7BlE0+UHjguOOLPFn0oZj7Nf70j1qyXia5E67q9nAy5z+kDNbk4g10VYzbLjKX4/6ufJ7
z2VEHIW3bQBbniH/huDWetXYihwztN9FBsdIm7730XSMvwooQZDO9mh6nIQauWsC/zUhwJIXp/Hc
TbGu0tq7pgtOf9vWgNSZfO4X4oqxiePeJrriA+syIAsQzyRwpbPj3oNUqYXr5FZay/e62nnVl3Xf
m8Qr1gwjDGS8fDEKhT9qpbz1NqgSaSBbvh9hmxbVLi6Vo7/akUL43WC2Hu58tfpsLwrT4nPf9FdS
bOzka4mjdFt0iKQKeWIG6v6TSk4vke96PABkFpDpSMbN2PXUj5WIFsNqkdBJrQgqA9Vc4h40EDiR
WuqVfmhkDtV4LeHZqJMO+GDzhd/6VvPQojbQdZ8A/WCYODYeQJYvHtR06fbGGkupExRzgZcj7mQI
3s5bIH7DEdhZuAh5aWm2YfkOb8Hhy2LSQv6ZmFCbdTizRK3VrRPUUvjEeeeKSebnM8Bzb6MgKOmI
w1h0HpuI83ODKaKk4C+oLRF1mDh7b3+Ee7FaO7Bi8WM51TeA+bwN5K7XjH+XA/oRZd2L5zwPN5SL
VndQOz5ojM6QUmGN0uLLVGpKLUd2ALiapPwtwyWYJSoqV7Fvz9ogkdBqyhuLihKx/jUc3ws2Z8Kx
Whs6GtJArHCg4CH1fS0IyU2s3LogzAaGWJBYs1O7Z4uLSCi0b9JvnDaspfK+jdrmIc6qFi8UOpx0
WylJr7cdXpbGN91BNVn4xDohLp03ldG0kUysvrT4UPdHaxI11RXGYagoxsoxYjZDxWegh8/NQbkG
7RpI2YW4RodDBm15dhtgo1Xu50FcwmOeliIjqBJHHcdmlilNpS3YnEkBRkog49D5IMW/EkeRQWYg
c4UIKH1jlKE18o/9KoZZezTXhTbkcUwkvs4HjVszUDcXBPC3aXozk1b5Pq8pUAg37Nxn11BxQBqs
6H1zBvfsQyH0VqpUBNAZD3kmll1BubFGCcxUA8Co4OuYPD/gDKruqTferp1W7L41zWiYpJWh50U/
HRuZGCsGPe7Rd+wHlgaoIlNFlhygQDQsncX6VIT89jT9+wqPuwR7wrdqUDzCgDZKOZuEE18QJmYu
MNrVWFzMQFamymIPnXU1whwdsd6OcQPhy8EZToSLDEhI4Rq0FGbdDZvH4Id7ha8uVNUoP1LVAJRB
nuzuutx9aye2V9RpjP6n6chULcEC55jwy3bOWbWpPkLJ8MlcfrdX6DN78w1BxR2dfeMfVV026ggn
34RrUPwNJwoNKtKuNyC9g4BdJFLtnNtyWcQo/UrDqEMmIZdZ8ToKa5+LYdet5hzATyiDs56B8Dhj
m9SppiS2LnAvBPFVae8fIgc6uv79jF7AsmPLoJIrv6n3+mYJp4KS24zZFEXt4gN7Z9NYPAVeLKWC
PA6fEwOTUx2DpiYewJquh76yH7vbs1Jw0MSYIUzOoNRNCIMb7bH09dGMdWIQ28lkZu7rIGrVLqHD
DNhqwH/mLwnEQGrTxEqCCsZ5ILdHvfe3RHQ3I8kS9eMC3F0wbteEolW9jKCX+/1j7F9cEy9m5tVt
IbdjMLAoFnOcoTOF4WrlM3T/QD9lCDqGgOyZoFy6iz+mSn5rPmQ2SiH0V+T26OpMuSJ71WEAdKmE
vrCZoUY50oddvV0eHpModtrUw8eKOmvMeAQuRN6ZAVVBlZW+sKsw4EIz55vdz7h2GyvFWz8JeDjf
x8YbM9XFjUWF3IpDHPDnXEGImyZtC3vjbxaLDDHxt7RVhgfMll+Tus10XQsuRn/Y8GkYNJueICfw
0ZPgfrxSiBjeFupvzHUoYkotd0Qa/cW5gyXfxLeoPw9aGAYYEeW1WDKQhJ3XgI7BjXY45gnqW/Cb
BH2LpxfEDdKJqj7udRrSPcrfMgpoWpEDiI/y33r7Ug/dwdI1fj8IfDGnG7C6DWgRxccaGLl+zr4R
MiTlD5VwBuzCzBynpokcxmwElswF2Yvh6O5r/rjDoN6pCIrVhpglMBGaTa7UHnZeB5GYA08dhxje
H1q8/1rFwbFTFqdFEOlNI4Znz5R0MFaYMs+OnJ3+wTIE73SeSLemPEHNr/FcRGGtAT8FW4rllYp5
+xFe7RPl4y6OP7VlxHpJXSwktX10/yTjvuuSTLZK1PNlKl3XhHK6aapXWIC9Z4kPyfrTX5SzZwTH
oAR/m3ICZ0auWKg2jFXosYlb5zHL/pMoM/6wMg9ffoDjRjSQvJ91FyPTugH8Q6H/kN5jf8f8jMtq
t5fGH6AM9U4SW5VUNU1C7sECzkVOqY8TIaK31VcKzhrbfUSFGF8cN36IwJVjjPUZXY5lfQ6emGPB
7yNpN4G3P1/qc8kc3gV7Aedpz7/H8ZeUPRLwo5OGuCOYWycGrhJbYkQRwMR8CsauHGGfCAeX0sxB
9BNLXBtwGm8rQz3PcZfWjTao0HYc6Y8pR3I8dPQ96z/uTJI9MW2jgdT1xzTLNCzHvO+o06ob1bd5
9EVLrJGumCQFhVqtaW0MLWtHjlzOYIOovcGGTiAGqF4NN3fphNNbSrAIzvuJvJdT6rP9gDAqZ4ie
nfxvyTnZepzCQXCcRNw+7XqzB0yPxN+dW9jgrbi0f+nKDiwgQOl3RwEqaUaFeX6g2k7GTIr23DrS
o7WYGkAtFbBBOhVsdc57yPrdmZD7eMYtCXjEFk7SnbIbrlDqbcqTtJjCi55lQViIUhj4kuNPl/T/
sm+pBxiawOcsSH6nejjSrZjWEMvYESsV9oy6Xafbup/GfrHCYf+1ZyaqCJreaTfLnv9kEQmBsr0U
O/2gFpoN9WICTPqDlrJTk2qCGqR/WAGmdJARqGF+kYoC+ouVmEe6wJ3RxO1SPDK6406MjKHRbacf
+UYEP9wCSg9rOBhJ61LH+pHbhob+M93fhxCz3gI4g9tlQdaG9W0ZcweWe4ynu2bAcwtEmAzn1SXu
PGSem0aB1Q4Afsd7ckY2GK+GV3Y5gc2d0eXfm7O9dBBa5C7+4eqjyH+2Wm3JcW2Q5BdTKKA9+mig
mDvWOyMVWTYOlgx99M5xvFCCrR4kEbCtUfCSU0UKiBAVaypd+HpUNqGUErg+0YyHdXLGdB4iFpYQ
rfLnB5iPAZ2MjVYMyZc5d/fa1c+zVgLGSW/qa8mYmOEBY758FnBJKu4pVWlmm7OdFlw0k5Ah7S9z
FzdZVc0vV/G6kTWiwZIo7NgoMeMXvZElpzo1/7FgAbfspzUG5mCCPjROpUVi1sBuGbPHARbN0ZLF
Jg+32EK8XS60+DWYW0Ob8NweCA5f3fTfOxZZYs6O64YlWJmVR1sNqVVIJKtZ3K3AC3GVtkiU2RhL
xtp824X0u28RrUYZ2fn16KO9+Kh8FR5W98L1pneWCZnura2mx7v00GdIND9dNlDxGXXefIgKj0d7
EWzPcrzufFWH4NH3ZPV1d289vNRPGdeP9GAIWc8Ildl72kOlnJ72TH9INaI7vNDhA/XzexBgiTPL
QHbPdmKEQiowMEMZAO1WOhOjwLds1duZryx9DhHrksBMjQyKWCdHL0wCixhVjzM2BTpCTQGw/3Rv
wLELPEM8sqfziKpmr7TnDb6qsvqLs/1OqoOhLsPQqd99xpHivneJL7Z6XmdexukXd5vN06VFS8Z1
4W6546siT4YIe42bYUeDC4foAk1Vg011pcSAyuC88zcZZamOxw/5j+qLCPaa1xsujjJ6xxBmb0kB
qzPUw4++MiFckIqYokVLJFZ7cf4WKK+GC9cA1MTM/nVq0A3Es3haTGsZiKkidfywUSBSAdkNg5pb
DDZqM4mAc4Z77ahA/5Y6iMCnEBQcsPw6Y/H+j1qBnv+QEz6QLzR43s2FLjlX75QWDCQRg42QFhK5
Qskjyx+WefkDcioGTKd8BqJJgZpfjfna3F6Vl22Ou0DO8hM5JYXbw28iosqMROWwSehkawaZoirJ
++dUxB7KWT9LVTfYNgx8WXlnSzeXcOjeqmhX3dGnxjas0iwugsYyiveDCvhuqEtBGhdU8fgYfhyZ
GkZ3y/xh/i1Sn/6uKz+udtdGNLQoLeiWdXxoNlTm4ABKRwOONGdRsqrnfbUDePfBl7uxfCdpaw3P
00X4hqow1cjyWQsdLozTfs5G3VCOtCaYqvqn8ruuheZwIgDoY8/XJUeXXbbDMDDH5/EHHl7yTsm1
khzj8n49V0fvcllNm5IwnBZA3rUpA2tqe4bGKtutcRMnUBf7heSuFlaIaxQcbRcn7vRK0Hzou3OT
fSlIlrqngwrl+CHjiZ2VfrKUL9lUVGGLZaIIabC+vjlrGSOvAfJrD4rDS6tcZsmfXoIr4iiYBKSE
QF2yFxLUTZ9vEHIZzze5O26DBB4RXicdYjElIqehhBCan+wZ6s2laWJs5SvzZl0Q1WUlkl2XbaEJ
S+qjh4z1tipE9wFn48lSTbwlZx3YGoKoDrXbFK+MVKMncttyyheUbGjRohTPo+ax0VhBG3ykldz/
jg3zSur0/hqln4H8wneDGHiB1RaTXSvcKY6T4MAKsEZP9Fc9KkL/k6IL20p1iWskPRBWD6ZQ8KVB
RPdW9rVFhI8ePufYu5dcgA1l0oAWAi7o5mZ6LW18jNRywPL9jbl3J7fmwetArVgxedhn3+8i8QSa
LSWWidkVO3ncZE87s+SXSDGAgvcIIQw+IZc+zJw2zYP3dU5LLkRDsD1AJr/t6GxAUottyBN1bvNU
30Eea9lZI75Q2CjIL/L8OAtqyK1YWLmO4mU/MYDBhiAOZgtC8f5xsxlfvR/Ni5s+WpsSqqItPquF
VQQ7cpeuMSdBUoYFJkG4T665rc8PbHtIJdJuM6oAhVj3a2lFUsLcV3WZpeJ0cxZAvf1tV3qBy6fh
8ipY62IKRnziUaPfm69bjMbsL9MkZTlfh7GhCj3igRYNkPObpH1QVdiIg2vzmemJdHyV3pxybdUX
TifYGYnPUD/a/hEDmA9yTJzPjptvVkWDJyJyO6NtcMbau0wi9DgcYQ7XG35V7+cfaEsntN2TvGft
1s6W335CJ8NObdZgaJcvl/sONavWUkRxxyp38f32wCAXd90qUaxcMn6B8nO/BE9RLILz70V+W6Gj
SVpw5ZB3R+GcZvljPcQgQ11LDov9t6DyMre8npCGCeLhAn8uvTGbdMHTq/YMT1veHkjfa943l8t/
9Pvqjix53xf0rpVUji0Qq9HsOxD1ff2vf83M39O63FPgs23Y+UODbRN/k1cyfIod+H5g2D9qgzTy
6cBU9wytYGltlB9a31oGmlhY1gczlQGfMi1va4ZrtEX7MEu3UXEdXcsWEoztGGXbtoipqWzADQDO
4/aGtEvTTJejYeMEeQXoySteYiLo+hb6kqDzvT97NTCeqUoDR2ZSniltZqK2rKLWXze/1Ke/t4WY
8ObW/leCS/g43QRPPIlV8VC4tKOYpM1KdpTzJjUg713ffpkzGB/NtEW0oYs8hUf1wqS/CRBFhjg8
guWRNdXiGpkqksYlJpCW7YS5W5oRxEQmDChGrhBsY2IkKNZ5KWILZs1DBkdN5PQoIIrQtYoIfWvc
smt3RXUPOttO5j3DYATkOqB6LfuD05HlB0EXeg3cjesXa2Z9NuwZktAPf3XFJALt9RQhmQMe8zzT
DKr3j5a7s/21PHArd2gj+NV0miiPIQ1IbBMZYd3SqZQdmTfvH29I750gTWoEU6nXck2VK+OrDDZT
Pm1R6Y8+8FlpNgI95yg5PxjzflBDdyYchDzZ9Vqo1RvIX4l1Um53TsWTXGteqA6xVipu0TTBf7cW
olzWQOlDiYBkK0LMIkZR6Ryw1YmK6XrMGjFv4cFw4Kdqin3cAl2PKjlvfPYy7uSsPkJn8Gdh7pBm
feZb8b1vBfU5jnp5pTftMIx4JmdHiHyiHqllxU2IMve3V9hgNTXP8hkY15KlArn/i4dCWlh4yzAT
p+VNkNQdcSNW1woWf0PVFy0Vnte+KDcrjpRVio15PGu19WR3562zUT98FnI5aq7Ms3Il58CC26TS
qpypHhhPIlPO+PBL9eTBWiJ6bvkRCW1z/5HRFz/RuF15om/r4vKyfmYpBomYUJDne6pnbaTY3qTn
F8xwoqLlWzU8AVwn65yQbzhjdQiHPHp1qvWDe0c+KhHtQJAlLvUL1nrCAojde9e3c5jLlR4PsuPm
Xk6+6beMavv7KLuuCkQ4Zh1Oord3AyQTLhS4RLBxvFhMw2+ksOkle8pYRgQagWEpq2jYWVTQYVK9
OMz86tUgHLMQPjrZQYw0vPXSe705PJRxr2oOKggTvrSCC5zo4KAtsD50wFxaKz3xGgGcoCX8hX2w
mqfK5EJuguxDbDXh3zpl5usQ75K30TOU+NmFN9plQOpBhw5PVu/vNzcIQ9QdyvcOUSkPMpDQzKD1
tg5bDRqw5YFySXEW0WZL0n7XrOLrYZMTEZLHJNn0MtyKoesbanOUOpdwBfSlFHHON36H9Eod/7vb
ixp1N67wCWCVNuK4fJzZINPQtI8lz45OYfJ9eKJ8VQavtpoM10wlpWXdr1xq44eRVs9uqCgelxCa
fJ1CHuB+UWYKgfyqA4ExnqgsFAw++VnjsUSfiQs5bvGTj6dqMBtaMwPDv+r+JYIC7JcujoyBbK7K
RXzqoox9jCObbEIHtSX7deGj+2ELUX5d/CGNXXRbJwIh1wJ8tcrwZrid95hBPQ8aKMKiCbFsI0xx
CrHRyWfDrkh1DRliGcDP11yuq2MLEpdZiRn8fzxUJ8cHC5vkrdXjytYYF9bytuiOIQfuwypXJXc8
VFxbs5gNGgvW8qg7GUPtA9I0UwBK5s9ps01p76LdsLuU3x1XHjLSv8+oortugykQGqEilmd1908C
0KXkspHrfdeoe87B8MwW0S9MEUTFNWKNo5/qSA24JXwY6QCMZkhwvkyXyjWhRZYxG86L/KswW2DM
R2E46rEapFA2ZuHeCndGAo93420AfbRxgNz383vA9cJXvhO6Wg/g7vsu+BDnmbjSa+lY6gUShq1O
fHYHm0nrFP1nCZcl019DgysJ6MUWJ8/M1Jt0s9Pa9IaoZaZ1pil23bbFkqMfuDDjXcXlF5jIxv2K
Ck1LwoPHFIhjFQu04GrqNLbiU38eUlxyG3Gx7G1qaQ0HX+M8GEh/7/A4yCH2n4tZgJaqqZ9zSWlK
LhsWzyX+wUcKqcR8vxdkhrkSt4Ga/Y9kcYC0AGs/2ggCkE4Va3aNxnOdDM1TjDk9+BhQnTThinor
oNkdIxCdA1oZ81qm2QQZFhg587zsTrs7d5MaHgCaH9hMUtr0N/b4VTBx64aFx6wPviTovNWJC1Li
F4d8ulsXV066rSMWG2PxYbpH3HvsyjMo+b+OZP2zvNjl9w3QRr/1taOXn0CSBKBbsrAplZZF9RSd
DzU2cUVAn1JPQ4GONyT9mBTAY8HXxqbgug504kBHSxJNul+I7BByyYqc/R0low+RoqHAlh1O7Spf
JPrPGzH9FwBXE2lri15FkOxBtU2Eiw89uL/kBEulS6MsEuK7mmSrqGGiBBx7ZAdSkGcph9CiFLO1
ra2QVKCdnru61J5k9qVV2wp294lj94buD/MP5QoDJja/PeNxBxn1uEeIRpg7+aIkJzfZSSt7Tdtz
sKAizpR+y7XN9v9gTk35AQOiHO2MbiYry85QSBvaQusaAZDhQUVlgoycG28EhwTYs+6/QK/jvTxL
NJJo6v82EF5q+YjFoLHMKZIyEc30Xz3UfGKLdCPETGgPnH42+IwgzSrzHAEufQeL+izCSipuFJx2
fi9K/XtHg0qkkLAJjeiSlZyPiOgySoylBNH3Yja14CefMedjy/J+x4tZLfzQ8X+qEfjWv+yf0Hox
PYhOz89zzDDqSMJ0LBDQHm2xGxwahBmYdD9RFnWawrPYCO+7RqyiPPur1KGjdjf5r6B0CieqDqdw
VvjFQMBwM2bahq5n72kw0sAkbzOr5aXrMroEy2ASUIV6hMYE6zvtqFkGtG80ieqqflvhH7zybwEm
eQthaOEc1FZMFsoWzeGmdXJQpsd+vDMvZVRPZCIrghge3H4e+VvgTeQ+JSTDfwRzLq+tJz5+nm6z
zDkbNwB4fS8Bgc5lBE8/w7yIPuQzN/pGmYWQR6N0HRm+HKspTdyx0kCtm92jeqJuJiMZqADXsQpm
8twzTzEcEnYWIWnWJ3hNmBuUySRmFTSL38CeWYqmMHlG9L4MKivHlcI2FeDXZ9ZGQOFEGX8Kxr/I
A/K+Dtzv9VPdyxEhCydDrqxzopDSoGi6FOsXQACVgof6Rbs3cbXGIZ7feg9upIrum37e+mFLyaNd
0e79Skzp5uIw8zIdie9iqeghho73pbMiU8L/6zvDghzpbZtr02WmvMBlRhOswg7TSKBSbd8pleLs
b+qKopmVO7PrMc0mr7SZnFwk291drjvlwUqZBQ1gH9pp1wC1FLzwj+sCW2KyZ4A6AuPnfApMIkab
OOXeyc+pVJejlRFKEuKca4RNQ9sQ7A0CWZhFx0AhOYFhdYDQPHj7dB+hmUVS1ZbF88X2suSx3wUD
4avDUaV6d8OP6kyU3mDoDL2js1qCctmGjp66ss3pBKQQcep7rEIGo2hkguktJMnPyEj0NvboG9dY
XCsSvRRu/G+XdpuK7BrGlsiRlW9IHpV9Kq0trzpJD4WqR0lH8FXKYY7HWxHubt+SguiXBlc8uhpD
vxQbce3lyeR7twqPCu0UWdl3tBZqzd7gATHihjDsQ7xZ3dGUZlc/QZKXKz4XcvessMIO+umDAlHq
JPP6jqx9L/oZ+/Srv8CKkPjMIbBQIlo9c/btmihvVaDBkurOr9cPLCqyiOd1tsY8wxwgU1sa0Z4/
ifM2FFOZV1VXAVI1M7aCk+Zru+REZ3ITR3pOBCbIPoxPz5f9MIfZ32U4ZmkZpY32WhqMr0ucrvLb
qymsjvdhrs30+T0/AWXRRt6JLwi21M5hKTFr7nYAQfSFe3JIGK8PNrqgSpZGo1nakkVxFZclSGUc
1AkZyC+Wp4lKTFIqFyqp4EL/lnbq+pCQAdc7emxrStNR0fiiWIqDgD1c0enbuJ7iYq/2yO+ZTEci
p2OttE7PrSU8tNq08DcfeWRIPDHQqcLerdbj+Z6MJu7YDXL+33+OA6J0ZemZsc8zrqJujmdIcUnt
Zb9B02B/ho6NzcZzaBDu//lJdxA4UXlL2/T07ngNp+sap8UisJv+5Y8giHhnpGGSCPqldavFqVTd
NE+TKvB+L8Pi51dV5gNsT0ToaK59JoJLBrgzZepXwwL/rkhouv2tA8+qAOECNHqCJEn2FtIo+bkB
6VKl16nt31bsLCr18Avh+0aSnRr9uNSqees2HorjF/2i+6OFa34qvrdZwkJwmXPanYcd5dPuPLEX
d38XetrpwlJXAUYJmsVjU4rDagaWm9V+pLPT9d9XcYxk9oKCPb6/SsL5VRR+Ac4JnYHU+q+OXkZN
a7hX0/pKaNlQy0FJPYsWIqMHvjouEGiEEq9/Qz505mttf771Qjjn1x58ZsbS799N3wRP0GJlOuli
W/38J8fFhW5QziaFHhC6jPfU518gVnOOaWYviHC/6CKp7gxNM/2UOi8nOB0Uw3vpQFuI6UwwXBkb
Dp56dtmZL/tLRJNcejsPGE/uE4MkklYs8dsGxn6ORj9ZRhe4LgFKF+2wMh5Hdj5xpJPIIJANnOhK
Yd4SvSUeX1xKk+EoehobSouDLv1C9vupVaNRYO68Zd15RnEFTcKTAzQNxpeSgJbxR8lCTYMLPvwA
f0fTxQKRfA4rsFGdZicffO1Dxf5xqU1XV7SVWuXBWRwVAJwpASZiDuaDqO6U1CdBPwxN/NjjpVVD
mCRhbKbvngh555a+LnYTzMfSaGDLKWeY4duNLfKjhy5PB/kzC8aE6QkFj5CxUamVI9WcTizSADdd
HocNCh986qXbikyg6k+0cX8r3NOFkli2U6gJhCQKrLGN9hbMwDVyPp4GxHokumceJtHWydGZlVt6
ziFTx9loVrOSN36b5O90w+rnsfoC2VbdXdJgNERmZN8Ey3CSS7VW0a42uwnqxtGXVa/1K5rno/hC
DzbFdHDqWGVkRbzGLmSyFoLsKdUHibddStYrmhf+Eg6+jkuFv72NkUraFpEd6z72OGq7G4JyHoAF
UtXpj8G0AJNav6maWIU1s2/eQPoOpXe8AGFIAVqY60PYlmXGoT9qJQ/k5Ol09Zu1hYvhPFt+549S
rRJMK4Qtn+reqV4Webs7bExo8PxHMmlMlsVF/P1Za7SncK8p7K9nwljG9dGBqZhz+7Vr5q14L8VW
1DnFXKGuNnfeH7fE/bvBr1iHjT+X79ZwLoIqMK0TdAaj4OeDFWa9MKh9attVgA7li5xsY4P8Fg7c
FA970rFKLUg5AJ2Oaf/7YFMSUcGUYhAcIyHhPkMg6tNxiSjK2A+GVCPwvZPkYi/PL0wh2fcq1aRq
A9aqdN8c3OgelwuuJlWc95HVRQMKBxpwQb9fmuxR/v5W95X89HcQ/SFxPw48h9KDqCL+8ePhMtu8
cFKkHbFk/lszXLRfZkMqCXJpougqirgVrdcJO2eHG8YcyEQLXPwC98RABoMPtW+URL7/k5IKzKjY
XA1XCnxYZ2z36GcHi/vRhncaIaWCqOorf9upp57Ay/6Vro7m6YEMZQuCnzRG6E/pANvPj4RoepTS
+Y83hGfp04GKMbO+M3V6tIDeUGT+jnDwU3TAKwUVI3aIM421penfAqGKPv8dx0h4B6OYZsbcIeXj
QK5ZRmx5H3c9G9eXdOZt/iK/am612LYu9O26j7wZSqww5bn8ekjKoW5TRih9BX5ounlGg0r6tdbI
29dEKW3Oqn6UJvpZ/YEaE1ABXhde8jX7wuqm8msLBwUnj9yQRiucyvoVOUQ5iTz2jLrR6JdfHWjZ
46+CTdlh11jpYMNThqSeW7phsxV08zvcfeL8KujAZ/cfp+vqIqoX77M8LeNQTmMNMmjaiBPFmzXL
a2hsXVaWUtQ9+G5FSRY+IwIODa0ImHc9/jQdmCOGDWfHYjTDQJW2XrpE70pxdOmQTyHEUa12rf0z
0J4oNQARRhFksruVe3HbRLtyY7yKh1vWP/f27GhncS0oazeNtSAQ8yhOiDCeYw6XKHHLBXGhMpO4
J9rebsOn+IIpb85ZxQfyygpqiycpWi+dQkI3c9rVeykAPsq/flHjSy36eJp9Y7w5VaurZHkkVQ0E
i1/wlkbLhOCH9HehGb6HCa3pW4Po3/liowykM/x7fRCCoRa/OFrXy5zeiZDcR9TWv5DIyiAnAC5B
PN0S+rlydtso6hd/U+MYigdGfKHeVsXO32KcFkR4ERptVoJkDvYfCQP35o4R+lc3VuzBXYqf6moA
7VuvhxD5XIfo4npNqTqiTiUslBqBZOUn88h3Zr2P5xp+ysICZH1cQaIdReYUYJY15Cqt+Daf5Xup
6pvc6JL4UaCvYuTYnL4VGlfnAcaCzwksi4SOkH7KJb96SYgU1TZ+B8J5MSearR2B0e1OjJB7+qI6
U8reoxGqVIOf0//moMhYIdRUvioTSWQOFoIv3Atv1v1uHzFMjhZGWwAn1OkLJKpwa6FY9SBYGN+c
jF6ZEzkLUydybH4Nte30tAT/iVkKHwQKYAaqaZFlgfduYH1xJqjV9eel/cBMpBVXY+FFInZpiZKF
FgDsl4xPCMOXJ74YUQGaHK8tL9YsBkxQNu9ksC8lCa5AhVDA1GuQ3j2O4Ht1o+7RQRjU5YmJgchQ
7VwCUC+K/Qp46VSPav90V7uAcWH01eIO8txRlYjXYSunLq5/DzDdcioiejYmYWbOz8u6wQ0rku+8
XGh5Vom0KCkh24Os2IfEtA2PmdzSjy/cxj4zVvwFYY2ClwZxweQqu0T8ScSGljJ2ohgGCnjPIZNF
h0kKDmWbMXG2dV+VEpth2A/IyJyHRWlIWO3kh6R70DHEt0h7EENl6gkCXEiGRPUj690B0URkKTBW
/BjF7yvfK8KMWn7QeDZgi2c+3zkoumswVlCkrw8JQkuQAFcSJi8LDQKEaswSgUVReCbuU4liXrLV
UFgD1sRCDGWyvMBB5Q7+LZ95yrDtDFqHNc4qeq1njHQzws5cI/m3tRZkk4JYmiWrj4DV/ipf1G4Q
sLUZTYOUy/XKN1JrXzuZsVnpAHJ+zn41e9y5tvNJ5+3fUWs9gD0CkdXcgHcVu9M87gxQkYEzD+dn
/1H7rT9R2xrfOxgNBcVlFRBl/tRLLbms2ZYHZVGpXKB54OZufMrI2h0QS9i01dkQ1Bb919eYuemV
P6EAtBXCdPJpZ9t5nNhgvvwr6UAKUsC/pqMBunwyB683zUFLbzY5mv3d4AdvJwBM6IQom88XcCdn
tMjzEenykVt6x/gg4HWTX/hFy5JXZHc47X9n442oHk5msX6otSWQu1rL5DFxj5DRF/08nIhkKQMl
OtGF+2xOBgvzkHkia8w03QxPuwQCVOg9lZblkDSni2OD4HPxcRuCpue1tBXHtiPgjuxHt36KeZyL
RM6MXajcrIAluvBEI44lPJ64DLipuh1msSqmEfQoH6UyV9CjTym0PJ1uViyvq7OluC9RIPgCvYTH
JyMPfrSWH81HEGV7ZAkzXTNyMR4MU6VOt8xDuHDtAQjzc7vZ0d/oYNzgqxM/2lD/nmD/dd11jOFW
x38q60X7NV2muopulBX7zT/4n6Q+39J7UwW66rXf5Qlr1KIJblhLKUeYRgRVh2BTiYlSuNOv9O3d
IniBGVL6GCB42dV27+8jIRc6cIj0w956t+tj0dnyTJu9eigQS4vn6GVocsv9iOiuIe9Mnr4fcE7W
x3dIlf3FFaBfdckz32o1/g72QpyN2eod/MmOqn1Yi0xRpuVbulPRIBF3mr5q0r2FMBvcQEPODpj9
jKA+wj4t7gpXoMYILPXl2NsM+KPqIOsrB5NfSweWJG/A24+Sr8Clt5qCMxx2Oplm9sUDLqpuypIu
gO9u65Ca3vni9LxsxcKoDJHpjR6Hi26GM9HIx7KtQhPIzkeBpOhX6UUM6UInTdh8upJUyCe6LhJx
fyrzfFkvaUDMR8rilvOTfs7/saA/JznJwz96eElrMTrrAdFNamgNRpyU3vDMndeElWetMW0EM7jL
6qt7lnWcIt7j9vgjt4wXKEbAY0W8BLGdoIDzqwLcmV8eev1encaxQW0/F50mxkbuDQ5cZsHcpWjC
SPZRZH1HR41lP2Wi4CtDC/71lX9vXau9LNflQWH7DCTI2Udp6cium2nGmYsa5yAt8cmQA0lHZQY+
Y0oupPbx6U882j+bk9erXq08EZOSIBfwQYogrJD2gpLJazRbRQg+ZXhzBBqrXqJ+VHMekrz/moLy
z2WRZlTTp3e9BT3KjmDZqWB3chD9ItTO0ztWKJG21npkjNmSH7divNymJ2Pv988EgHYBqnI4Bg/w
KhxNV4p2bffqkWum8YXAKIvIfhxJXV/Tlwb30IhujKo21UFTo7wpDyxarRFSOYdQTu1OGT6U5OHA
FM4JhZK+9iv5AYh0Smi78gq+Wlr/NtQ80/0nOlI6V7E4E0Rl0p/OH3C7WKdjkLS20ks6l3rYpwCQ
vVGZlf9kwPbTsNuT2dyPDD3mt1l+uIkAVs54nd++ZG+RdA6d8doT8eaV27Ybrhsk+MF9uSEFqQDr
6Rl3X+toIwT2YuUaaIPI1ieFscAxQS1Pt5UJRtLy29d0MKFI8tj7afMamitXDGL3f6BCoFH4Aoei
lMkuxIzvCRMCa3Lnj0o0rIIf0ZQwODWDBEVi2VdiezHQmUg6N0npGZ3oORpz+u27cd1UuprKqYWh
mhAMBcgO2E4GCR893yU39dHrDIeXnah9kRhg7GMZjEivDJa4RgXnOb+kQffqMd++Lz9NaM8Ol3lr
m3+97HLwWAY2SNgdqs1GJZGryqffpdzREw1HlXeJSIQN3vL1rNSRX3FTFPx/Va3KbO0qJLR4ZoBr
ag9F9uLx+WqLhVe/hryZj1AkFq5KenrHEUznJhLA2OygTiQdYp6lrDKUCJeNPfshQEKhW1fI9SjL
nEZYzCDHCA6lU27c4I1LF56Du6K4joSArcA7NLAOIt+Dugfezm7u26JVJMdjH09uwz6PjWDMBM2V
O29SZDdtREImRLYSJ88D227sH4gNGgFQHhFHHzIFRRTbaSC+2y41z/LQReACX0NH/wlJgrtFWanS
1pcKEwaqjrGUBa/lWUd3xfzGrnHsL6TPpgmLHk7E62uPS05/2VCKvVDzNhxq+y0sXaTW3mSf7l71
0jjnSXU0tdu+EddcFoY4JmIwNrHiNjM2GeDYN4CM+CS7IHRUVqm1uXxZfBbp9/dMcDTVfCJc6arT
SxSyN4wLXztvYSF0fAFFpPV6tBizz8fRUbGYjVL0MGW6DLL3QIfUaYmqwXSxbaNzesxVJOT4K1Kq
BNKRsBylcG3G6fUOXzVxxi3Gxlkj+TL1J8a8tgZs32ZQhReKo5ul6uahc/qLAmzzVqCGpDx+MXeu
Y4teq0Yd76zk7uJma1cf4LAZ7ymRYIeHkND20H4UceI1akRzGDfddU9GF8YhpAcA5n8WCU07sIEr
gJx/+EKm9FxeMMH3PxxMhVfj9zqR5Zd46tD/9KKaS444C3HyLDqBxWLRs5CbqWpeyfB0ESq10oVN
4pAYHnagXUksoEq6mK9Q0ApRKBjpGuFjhWJndsN53RrCUfNZ2+6fMTgC1GWsxTKWHdkofvIzDz3D
006cnHdsdHokyffYZ7jglNqDWHOqWOpVkk/K/N9IuMCQGBgaFc2zxxtC7Xhk5kxZfsS52qdQ3oGe
WEuSmrR+yTu5CU4o3pHq+Pa+yYYitC8aC5gIT7K1G5B58He2UhLyG7C97rwO4XDNhzQiMyCGN6lU
ktP8nleZeVyZd3t6Yzkx13TfdQYwYmi0s3C0c6yWobgat50+7IKxo2objVGcPa6/1dufBN+xExmG
S0hBhVE8jI8/leRgkhSB7UoRUjtsvQJB5l3GIlGXYGHaFR7jqG45bYE5KPH20lHsBd4PF0vM0eCQ
W68PW7Kz6TK+NZmvzCu6RElQ2l6p08u19HGxVRwFgcP5JyZLAe9ZlKjgfQ8lESRoL4VcmL5XByGm
krniUi8GyrKukLQQx4HZVTMRsBlaZkbszMYoI6Vnz4lXWJ0/0ck7Hk43afaY3tqcxI8NO7asSJ4L
VcTalEhCOjVrh/9o82KEHfARmDo5vwyBSqMZMscOjer18go/143WoRqU6CZCLZkYWVNjBR7Zs25b
+Pzr0jDaUjymFodJ3M8yfHhziui8NBS7GoYeqewR/wTi8kBrvUL0EV+tvnVDXvpKdeESw8/8Bwqe
fgkKnNps9UMzJFh1mKR8/UaEJHNenVsLp3qsa13H0xX6+3gToJi5TWCy5//yNuBnAhZJMsjzeoF1
fMTQYbGaAj4ujQVcH9NaP1Zzl51+kY8PRnu0fEEUHlfiS2Vadbvqm2XGiiSWMx+/TKg433nR6Eje
aKL+XdZmOjF0N8J1JRve5+4AcWRJGKD/Fq3x5bJgtk9uPyD5Bx3/xbEkJ3JD4p0QvbUT6DbqE7p0
q1KPzjHBFtsqLjEX46sDAZQxEZ5hMX+zWANmPMm7RroliKhLHouk5Pb2Uh7GgeihGwXVmeYQbl7F
/WjDBtP63lgGSBAb/sMN3aIFgJOM+eAJF7no2U/wPT4Wa4S9Yz7JuWTcUCl8expMz2mVSDYJhWHv
LEJ/ZRXbpx2qBDwO8gU07mM5R60C/2ABd6JR6ZXo/CDGZbNe1+rfO3CxefN7kwnwKGBzg+jLupjH
zbUrVIdiZbCYxd9yLMKp3ujBLnhHGf/HvaCYxqlZQqT+T5d5udw/Bs8OrZkup53kW9uK99AnO08M
eWg9WR/ojAEnBRDzfK65G37A+03RWArameRlXk64I//8Zp/pcS+AwZoYPxTBWdPxfbgYMHTo3TI4
mXPv9f8EXqWeZag1Did3YgwPrVLPHBG0F7J5Bw8A7dPULtx/oR28mvPuJ/7kOHNJtVE2ZCAMLLJd
QFn87ptMnWQBCSQg80Bxr3qVNsxwARF+v7TWiFSaSz3SY4m2Vza8Ve4p/TFPjmddNsUQsxpu+Li+
xPnA5L5vt52xt6EWy3SaWshikAtqMnePURnLDYs+h5BN0zt9Nly+Mggrf8oxl/o+9oKitiDrI4zC
wmAOIYau1alNNswHcVr9xzpA4UVprGLl9g/YKwHG+PrtBt6IF1iRXJyvM75gwAteb5Q+iH5D4N9L
gr4VLQ5ivCWyqY7oby4ACjHmRADcqI1wzxoGDdFkDlVy+dDxPQX1T2GCCc5tKqVbsUjpqWgqudXQ
ET6rOoKfSxPg7TerHsIzyYCJMXh8zdhGdHKvj0ddt3ysYejJxbqrly56q4L9+T34XBc2RWP8y/ZL
aJ9SRvbg+oEZazbc2Bz3Bt6GorriG07j7Uh4f32wy7uyq1LurpxiZtOotJPO7x47a2TAkXM0pZDc
tUzz3tCvYJCJRZ+WcIattRENcd7gICplHJk5Q+kWJqNiR2V6d/i7lsGTiL6X9sbuC7nNb/hc4GLs
l6yc1e0n99rMF3abn5aO16KXnSs4a5jnsYqEGLuo7UkE4AYObVMJg1+4TFVk9qmdXJy5R/YnAcda
x4hMW23raZ/R5iL+QAqTZ/MBjMyZUt+MDBQGhMgy/2GWmfTS2fJycNQTt4vr950lFkyN4MA6Yo5/
muVge0pZhbhp/WNgmSgUA4XSV+2OlBVE15bBa94OC/HZKQ2kcdFckHgXgXssL8lPBWtCn7ZYmBiO
LjK03o/05Ktk2mdqfpQ7gamraGFLHovEMLwoNFWUS7iNNP7bHidyyb4SLzOrouoVra/23pVEHaj4
7/7QXUVlyzlMieJSOHP5nhmAxLdYeg5UNa2PsqPO96vH6TLkGXmUtRW2rLnJqGcPvBnC/Ct9oON5
MoLypxwrdD//D+US4WfMTtWLJUROnXwDasgEyMunT+wgTTyjs3XHgcP5KJSeHRJ5G4/xtCpGSmI4
KljLdtSbaxEGUfMqrW0+DU75XFgyVMsHKxfK/FR7i5KWL9IaYO7O+wOj/7QltWeDbCVjxFHvrdy2
mSm8XU932SqEtNf6ziWsuGenyDT56GLWNNzyu7Pon6kw3A1LoiiE+QJ0inwQWSZb/hezEbrSY9Yo
H6I4wcZVTPNwODpfce20yrO6EAp1RUQ77W5F9TAdrtG1wNoAns8O+BwAASkt4WjLNWNbNMu+x68X
vCHI01DchmjWxhymK3CSlz/RZTcUiDy4xB2v5OfAk94slgm06DNr8tEPp1RI1wKndOXY+vg2KJCX
QIohkVbShxrVSzv2IyEfYiYfptF19WCS2bpAMIrDZzBFE7cBXzH/kKtn4qqQ3AdKGNFp4jlDph+I
Po9oRHGGuk2UTKynGtAy3OTjSssCbe2YHD29sGOENL3B9SzoXbBAReKILAoNKLab6znXNswDOzGw
TyJEYckvsHLd4FjEPyfVPWz8k16BJa/2sHwkVU8Y98lvVBC0jo1RdYgaCIain+YlOVH/PKGw4eYF
O+7uBF5s2CfMZDHQQNncZO9ofOGUzd49FASU1kZQoKTQBBAPJtc+QXrnHWrjETTeQJDp/u0xqMj4
iXmwzzXsjsEc7WVwtWABLl3gNKRxhUb+lq+i9AD7QIgGPk+hCeYrKxl2PijtLXOEBmDUYMOeH3Tp
8ddVIFACu5sktGidlppBOcIUw4/zgLeJ010+KEdcalM4a57741vNfnbADBUpkmiMMIGdt6Q9xUuh
YDxpJ5e9TeooceJFGimYgM51XfDjOkqbEdUSJ4FZmdaasgMXffNHtm79uNqjnWiazDCc44UxsJUW
cOEGom2+H8a5rQQ8pmrADAzwlFOduRV0/FBnCdGgrxD5MkPFbB2FuuGfCkiyadS6Zg0fQxFkmqOO
vot591Agwk40wukk7BWJoTgegwuGEGOgwsYI0mBOD1xuF+yCYPFFuNAOUvgIeSA6fQNt/XtfeNPc
eLGCgggoxEMzi4D9f7TkYhRMwPDALR4/3gHzkuPlPU8fkW7eOuoKshzenV3xxDCahaz3b4qtU2ec
uo1H3iMaKE0dT4MEO73ogiy3vUZhf6ejt/2bpmzzeqU0aOz3UZ17L4U3s1MlE/BgZylJXGshfaAS
XyNsrIun7iAqHMAU8HJkw0hy74wGnGed05n3IV8oLfrMo+tDRSdbzP/pgggvexw8UKl0yDu0Zkw/
NSXFydndHLf+yy6/afC16D1Yek9Y1ySJHyhEk3ehmEEDd3DdAuB5J4IZMjXJgiRZ95TAzCMChDXZ
kqWoGxUMaMK5PE69wzroKdEA9a/z2L+ITdFkwRVaHHrevH7imMrWYVhNNre16lzHtC5yrd41+zhC
R+dXXQNGKh4xGQaPks2kZf7fF7J3Js3ElEwlGW0z5NKo3f2YlcvKh7s0129lhttYOYH6E7EL+4/E
x3UsZom8QPl/Sa3gfkCeK1euPMdUwQS8R8ZrCeZ+BD+iRn5rAo+Z1+jbpHz4xoksVt/qlS2cTaOd
Gv1NOChIsyH8kI9FRDgSYwA+M3JP5W3Dk33CUkh7S4titTCUzaNdGXf1HQETbjwTS0YOSFu9nVa4
1gKGkf0PUQsVFgPotHIOk733o1z78ml/1Lnjnk2l7UL8MBK1EJO7r+b/AAupIpm2lyva73hqUt7l
Ohup8mIPoYB9Caqvl5CO/8cVGT533eoxLJ8SLsQYIjZY+XDLTN7S6iqBYekMnQGabudO6Du26alL
ah1QDBZswXQkHSkdzvcNbZcnFB9E68AgdvleGa5LMQcirG+5rIVsU00+gpPHdjNXCoIJufJPxLhQ
nyEhVPl1ABm6VnsItH7h3bdhYvilLuDbMCIile3o8tIoj1UdKB7b0sUD3+D6S+DmbEyRxYHm9XGA
sRXJ+YTyyRtZnuFHAgbwCsW86+Y713z5mLV/hFH+wU3hwfcWAKnLof6ncaeX+wFja0KJIqmGo3dq
1kCkaUNtBU9qqcWri6Jmh5x6zIgvSF1DIE9iTXHTaD3wLHqF8PFU4n6Vs551MK780YDAdTES0EBj
JQEHtpY4ktqySdnAnXDNyzkCR3dKc8DZVssckYt1iaKaTRmE6wjklTikbR2WQlVqg1y4pQp71a0j
MPCPAUm03ZILi9OwFjW69zE8MAI6WLUHn4XJ+OfXxcOTm/yoHKhfd7jUqW7F9jph+8EY2t//UunA
FTgd/0qwb9lhKgO75wgvTEMPHwZYm9XC6A0MPmJmd2FxT8g1bqvOIN/TJNf0J0PDBZ2Sn1Ze/5XY
hjUwufhgffpoSuDJPn5VYsWUOJX2LKEsSm10v2OnjFkdGP6b/1NySoNPkTCWSYlEIZjD5a3qgnzV
T/lMDusDO6lq1bXR5bSkkuo8xZ906wpKaKrOZMz3UIGaPJPrwc/QH+Hnt6+3giU2VpWMsAyWOJig
yR1p25YDITib5xBEIyGtfua2TejwvhthcrdWfcdQhzGBQzftVf6PFqsapXwk1Le4LXVEdKeVnTES
qu19BsgQWNeLGKqao1J3xb4+eE7/4NHv+gjcWRTsW0Zk8QznOp9KtGQaSofwvRWqpDutoDSPDVE0
YF5f8l65wEr6IRF+hC+78S232pEsoz3aND2w8tnzQEmKfB991c/M/T/v9Nk+Ic/hlhu+ZUYU7Ilk
yUfqfNKhHuf+c5mLLLUXQNsq8VkkTNILJD/gk6Ek1WYsiB6VL/uYR0rS+isjg4uCEA66KM11kAF7
cuINZTroSMUbMF6Svvt4syU560hX9X7iNbIQizOSydKl4HpzuDYVNm5eRe9Q+HTo513OyctlEVhX
bPmHzkm/tExnrTzzkYcD3e1LWdDAMVG3JStR1YCQcm3oMlIvmgxzfmXdfCNPBiFEBaazCaEJaBVu
Gyo3GjVaxH8703zSHDck3ee9v0fQ6dkmo2W5H7DRT9m1dJECIvS2Sa/PUZSLl6oIgDSNj/kE2QUE
jNbxnsKKw0dF4eMfURDffgm6p8XD5ExtugG0UIOuWrL+J96j4wkUZY+Ipwme5Va0asHw1meyTCWK
EHVy+619hBKdbEY9eHWDaJ55ZZpEwRWQvao1mew6Y3rh510kWjS+oUOdF2LCKdVsCCZW4fETsEf3
kDF8f9PdK+oJkkR7JZwcVDyVIU5upigF8QLbyeLVDlcuX7D9KVPQOMYIcadKeoV5jfnnJFhXr9kH
2ZbIxeloZVulQYQ2FkVVb9VwlFlIuKyo3ALMl8n2Avecm6VlnK+z0kKRXYZ3PJ1p8zBlf50POhHs
UQFiuCU5XKI8G0MeTtuHOZ6mxB/pbxFHjKUqa/+lAXpCU1GrXcCLd5rO+sRJ9PRWKA8BirJmHjWG
mOKv5BAsRvSzfAKsaL83jP8h7fnR/Gab//VZuBta2QWEuWGfwCZuCndMxiEY2FJDJT5bcIRc9VmX
K4bHdM7/I14MKLXbW9aO5XKucS27KnlxESkYr8LAmHySC61QVjKIiFfiGreeuk5ZiBkEmgIEhXBx
xxlFzh8hq3awpbQwPWm/ScQohwwP/XMCLw0DFZf6Fqv3VvblWB7e250PgoQuH6uKN3mY0ngT29cr
P6AA0GjiVEMHlHJ/ftPvZQunBhzhscPG5V+/Zck+RreVO7SnRq0L2u4ZL94zzNJGBsd1AHKW8sZg
nEZo6m6XYneumakca8rFgZMjWa6/OTIVBVcdfDwHZXHBPDa4yjrtwax9MZaXF8so83JDulUNyNzx
yRRN1mt+e+dJbv7hpi+vI3r1TP8HUzLmuKipqBsPCXeWPfkA7M0YKFon/cpkZei3oJwxsKlY3KhH
VCS4PlpNu5BEfWdDnE1huLuXYCZLmbh6VXnIvs2IAJflX0ydOsEK667jhQNOLXJdOZltYXILFpZK
0In4y7ZQXfD0CYRrYkk3MN2U9GyF137Z6cGsC5DrembvYDifS9p6byuyLghKuZB1R2zFKRmFJ76W
dkplbfWTz9t2aHUMvSLWrM5gQUtwU4BgkAG4zbUqRebiv6Tst/Fntjy/PWUdRANilaXnQn6C+RR5
AD5MNbl3n0CGlY0vjD6DvK1uqErAzNXN6g8teuJFCWNPJjA98N9WaBXhxiDO4K7tC7ql6j7rJKGh
ZCY4yNm3iUrn0HVVkKID1guhTGARKTgbS3HEyO90FjchAo4XypSpAzI4pji8Y+OYBZOuUHiegTy5
yG/3zZ0S+EHyptI+ZkMLSIC1dsOKwrpdn85keWo61NQFDaZhWW5xRBYUnAp2ZJZQGLQv7ajJojM9
Z6VPQY3sc2QLfkRSJ96ncTt+ZKbwgTQAPmA+FQh3H1ptn+i+YlPIbzhhs7HOb72UKVUhIlBH8b+X
A4Xi4VSiqAk+4Sjft+bsUaHaiab3RGO4jgn8jbKuFAhLyWiQqKCLN+K89vghP+1hSPvZUr3pOnwp
y9rFLvQz8DFMaZug5mIqW+E+GHLwdMUehsu2fWzYF5SqvhWoSuwtIdm+GrZT089hxrSqLNxrpB/X
WndfZr0P5rBW9640DZv8XJrgfZ0+4t0LOOoKgYN1C2FVn16bEW7oscfbGul0ARN6Rsz8bqyCmvw7
Ys7YRkRLLNQsrxyu1drcJR2YnGL5E0oXiLj2skfm8balUjeILTyjDM765bfo/pESzKYcBwX3Tdkt
pMHR3hTAzv/LLV3mVHZuv937exvWjHaMRj19vdjZ1SBh5lLuwdRL9LnhP0S5Bs3to2qWqsjmRjU3
e+XFIxM4CMw+fdgTwSLDiBcH+zyObUdF54LrAzqZvC4zBj+uMibDwFsvaCCbkI53HrezS+xiGiFd
b6EbaIh/ne4HcvVDkYidwougnOYnh/lJ4ouepYT6o39sCBbPZWLtG1a3HIvw4/zpjP4tuOg/5sqV
v84CtpbCswqNa+eErefG+p8FGFpYNequfUUBXSI426BmWXQJMgKK9v8mT4DnqK4NQ1QA5B2PUSo3
mRcjKvNddmjaIwVxvSPHMTSrSsWs6jPqnzbY67koRp65e+Kyi3m4YUGAKvplbpzoROk0broXewZV
rl8XbGKUQxaQzMC77xdEwMJmhA5wiNhfuSjF09e+mu2sDYnj3mnKN+5QUcHZG9B/du4SF7+hvk/f
AmmCI6aL7EwfpuxeYJgDlgXWHEGVvP56Rw0lotie7qK5Yr/ADFsQrgDduSPUO+i2YfJswGe8NLOz
oKcLiYyNgpNxUy4omaFfuO+ysVHrt8fY9Ny3wq2GnMq58SDytZoqiIfRzRY1o6nND2YI5gFz2XAY
KNCtNtSDuiBSBFBCXVBfNlJ6ij1/znQFjlk437e4lw1tKC45AhE++ySQu+4rb+Y1en1Vmr1vPiwL
8A9KOR67KBe8JTzMtVPA1RiTg6gfe9FWv7QdJnlYQMR32GNrYHQd/WzRKPKOhWB/oZ5l0bsKGMbE
nWKTeyDbTnLUD+swbchPfPnkElapC/8Qgs5X5JWzX921NLMYzbmBXPQqyuUvA/QzekAhJYLS6LQ/
7XAgcjQBo87jLt8/QuuCpOhcGvuAEouj+0UtKxuBWrr8LSC1JScgBxjtObrQ6gAT/8hR8xRuRjLS
4eCow0IDRRvYjNGhCJyNGnDJ9CEsDEXB3PLGCOkauigV/hK5qs82S/a8UgiU3QaANyJGLDa+kasG
/MvK2AeRS4WwV4uUzu0VezycQQOb5/aErCf399ZceSCcvCXM8BQ7jrjSfxrulLdOVK0XIK4p0eWe
4dOyQ2yO4ThbLu3rmmUdxX8qyZSTfMKMse4ksHqIvHE+HThUM7wRYQiExF73zEtn6zOyWdeV3gr3
0klmEhdTdFj/H8Ss+dzr9rfoFtFHyN5jtzhsUMxbE/WpfnVYCjycQ7pODorTrVO23osobiet6TLd
zZoI7SpuPTnoyI5em1/H49F7AUS2wW6sLjU228IurpNONdk2HWpOcC0Z1aqNLFuaTn7OQ9bS/S1o
qL+QjODMqWWOHONFjTTCdipjQppX30G9M77F0NUKr6Oox73dYerZ1Im2BmiZ49MzA40gNS4OOebe
MT8myajyCsXo93rkTlmM8RBP5Let21u1vFS+R0D2I+f7ipSGpcSZaw/9S3mhC9xtJN8VcC6IwFNp
iGPdZMleLqqUoj7XHI+flrflp5c+70PbqEJQS54OiLh1CyK27GhlgOC6+/2O5VwAi9W6LBx1Yz8N
WK57vcXLOhczPh/FAmkfZfA7G9cG16qED9RfJeFBMtBBtwWUKpVm49yLqqvHMW0Zu/bs946oMK2c
2FupOgDSLuC6Zw/ZBA3jaBVN3by5EUXT3PyftIwkEKwGRc/KLhzO5teweYhllCgBez+hKlroAYVu
Frq7Q7MClZDaoFKNpvPj4qoMcjAjSyt/WSLaMk+4UtNXuR0tpdqry4Dbn1r/56ioPrwFS5ZZtOAD
a/phCYg4tPAg420cU602XpgbBiG24ZjPr7za3XrYHaDC78jebuskH0rtAVCv0pgMyJnBnQNCjgMz
V0Er0B1su6Zm37RM4JeGh3+ntXhgbNDTHbT5AvnFcmeQzztLcvKoCR6DT+i0LBXGTPA5MbHjcyah
EMClRrP30EBCyQnMObMCSrXVDBto+3zeQU05HC/1bWFy/dGVXq1q46BZit8mbx+x5iJENvVcpiot
Xp3pYD8lurcvHsXawfv1Oy8hrEbegE37WwsYzIGXa/+PiKFglhYNng95UGKV6ErMbUPfuTb6VWXR
1wLmzQkBLhDElNHIWUL8oRMxIWKzvGxZ10k1PNpxy8rE50xTflVjV//ROSF1EBySERzQ/fk2ZSJf
nXUuhsSoY9GxVEHgsK/9TCmdxpEwNM0AkhonjNvtVpj7IlOel5rQcv2bKRMuLo9L8/2a1a/4jrKS
SqiXD1CMqsCkWXy/p7pqqcXqivND4FI7pybpDQ2/N1Ru0/k6Rxuy+XFbkJspMxEd20QtyckNfhOn
gw7Fp/b6P3QT1MXiP75qUcNViOnZxGpYsWNFm68wVTRn3OMBGaYKNTZZA/v3fekdgK54kjjxt7oi
oXKql8UjmFRpQ0bZWLmd7qDkfFgRcGLyxkfp8S7zQ8bd4bnRL6K6MW79jS/h0dA5WeDuZR6FQH2R
Zcj2B9YhAMaPTaefyJZK0ZYiY+j64vIqL6ZM1QsvoxqGmMW3K73ngBuFqaDWbQ7bzs/KXzx5SIWJ
4o7UoeNjm0t6dBNL7oQYHolbt7ndv9S2G4fKLipsFTE/R8WJh3ZT/qI3HtnUHuqFKCi8Q4zZyrMv
bQbsz3FE2RF2QQ/3aaa76fGoaIWXRBXOO0KEqyCRFr6HOowpccktsqmqcjNzqnMIraBsop7xKSGw
MLfdux72IoqNTGTxgnkHTZEaIgvKqo8GhY17A4Ji2JrFYAkUOJMbtCxLmUqRayVMKwkm8GPBlpQT
YcVp2LEIV5ctwqLDsAscSOU37/eRQUvEnNsZoC2L5EavrnETQLqpDDAxcr4lXg9Dz/CFVNuEmEFA
Fwc9IztCtc1ezC2C/3XUDLUEZ2+q37UMk5/y88iyW3avUoxNmcQwsYv+M81EuQEk0TWGnDjRHXEb
Fm/4EKhHbXBfmOQyhsryN4esrfHS5vrwpYnpJrr1/I4m8lZcfonJA9QSz7711ndMODFHps2APK53
eH1dDu9JmTthZJvLwitf/BaOKPSOWwvZ2x0Vl4H3yYq/82VGkI/zMhG9nZvjdODxGksKEwQ0V+hL
MGF7ZfeboV+Nfse5V7JDk2E5XlZcMaI8NEG03KXKh0wlIhDuwvK0O8Yo4P++UD2djpIvoSPOwNvb
4m8Vowos0Tw0SLk58GQ2XjlbOr/V7Eev5MZ5Y9wjgCXqvjxtQfw1eGmK7MfzJXzLZbARLNqg5c1i
iE+iOWF9CUQ2Z25K+zLsmN6P4IY4zolFN6HKuOs3ZGl9uF38SgNVmusEgK2JXJ393A1x/q2f9W/0
4EigeXT9lbcomcm1zo2Jsf9wzYpQJ5BABEGLE3HrZkFuoMSOUfBTFh6EGBSrW4npylD6d2Sz9pFN
sLNK8vCv5AtGHSefZw538rkNZcFvQqNlfmvgovMLeaI90JO+s27yjXcL47Ov9fBHWpvdR9joH8fX
O89LNEHnEVIa3e0RYRIMt8wV0q5Rx2HSRDO+UfNKJX9AkkKAspkta8sZOsY6unODsh+Zr1N2RgR0
z6tqSvdaKfPw21X990I/VD+G6fn0xz8QP8EZHyufy0iEX0DXs4NcIpyNZtai5a4nD3T2mDwjMb7y
Cgh3wkr25arsB71kJvhhHEAeOqnr3ROaHU852MlmKaxf1YF01SeXEBYZOcC1NCaICcpuiaQWdndF
GQ3LYnxwNPt6KKPX/bME8NX+ashRL/J3zK8Vr8t1flKwcm+QI7UVsKNhXYDK6S+bXbv0iOI6mx/3
F7uVL572GvJoJm56IPWxsFSKpT5appRzXNUlpDtAIMLuc6wfUbsFimah0cNSj2z3U/NiKWg5t1Fh
2PUQoWAwE5oPrpTdBjAdqhmKZwtVmwBlTa32xyevRCMYaPZ73wZATcW23ZlzOM3wazBqJ2Bfm1pK
72AR3klpMoF2uCHNhB5vltd/Npqy4vWkeuuwmH5CbRdE5CrCSnscSsi5641U8/XJ8N/gSSoVSJjt
A5+o+KuSyV4AYK8kuJ47U1k3VfWSdJpcgx51G1MF9dZohZWzc9PHxt6tVOkvXV+TGTFQ+tX3XBBk
RBiy2rOYrrJ7PMnO1/y/mRbuRkT/G4mlf5SOt+dtG4WP8KoCFR8hsKd21VNdF9FptpCADFS3szxc
u0fDgZOd1WAI08jdqVQZkZAUiVcbez4IA7GY758gFOJsXCQzNNauArMS0iLVPCyUvgxkxPuerZpx
eFB0/ltzmSEadpqcgJMHccwuELas6n1l5O3n3cbNa/tAxjXWtg4vdcNxB9Sk1WQFpjVcXtNPfRLr
z3C2z2RIkNTJcwCy8XRi5Wwr94Tjt9jLiC36RpneCgfO3GM3f/OfmCDFiZ/T8esSdEE2W1/p5rhx
NfEeM1pM5BhVuELRWIJtB9AbstjPe3d2lrPWAs3CbFGxF4BMCBs3mWdQlpA34d/RV+DZ68M0ZXzq
/2W7We9/RnpK98yZUQ+f7YnW2nXQTusbvb8/bGCGYfewrxLEoQ4y3cnxnHUI3g0A8nG7mx2wB28X
IXLoa5Oxau2RySrEfKvl6bpQ6DZbXBg2a6TsGU6pbuOd0ZtviBvx6mIM1TkRXA7y3KoLhh2gE8HE
xUOXHotk6Nm5WdgwI6Wlai4IAKsLBo0k8ROfQf2JnV83bEF3fla5t5PFtJTf5xvE5dJroX1YsDzH
vPruKT+lN+cTmYFDsd8kpzMWMACC/pEYutXczxSTfqsYIaLkd4uUOnQUT6FIvrYry6edYL0jmwvv
5h/AHG4lXKLhDVFcpYgvD7VG/4HdO28bobOtlq5PypIJIiKvpjZgucQO6uWVEVwF+X+Twk1hYJ+u
qf1pB77tnQNE5kaBW4iLvcikUOSCwBf3NtdHzNcAdR/nwQXeLM+DxaypX1UlJQx7hCTExumNZD4j
f+mi2dgsbxPU8HVRkwdNm5K4qjscqNL6cYl+PDvkMnRJbNFBOeVU97MxVtukn2CXzNfjoBias5+W
zLfhR78bSjka6vBxD4viY7FlU5vu5874dMtJp1Z/sw1szdUHNvCjk+CMhj/laXgaDBj2J62cAaDF
2jxqhnr9jO7KZVVGDCZQ7kuXgXVs1W1pRC7IFWY6S/ayC4p3bYwoTn03mRnvo+olTUrpctJvp1t6
BhjSvut+lMWVys7m06xZjUw7Ad9Blhy9R0hFL7dsJv6IXNX2/PWK8js1tK1sMqLnFXx1zhMeEkx4
1v9qIcrl7a6O9+H2iLWSQNwiHKczNzPN91aav0Z1vCHtH4IH2Bn3FmpynEX2KYI6mDp3ZudUWSnQ
q0txZ/WcSUrsKMbon27NQ0+mNK0xcegCLBIMyq7nZealM82MFUpTBR0+DzSXHVtGOe/jmoLUwCv8
UOx/BUTSJZprnaB4UIrBwgmAaQM/hdphfv7mq50A8z2axInRbNYLieMNBkCrvUVnJjy+tEcx4UXd
Ds3Cgdgjfc1gMUyyJHM0P6UV2GJPxha8/bM34BdvA53a5HFuCb753rbbFn2igFDJGncq2Ty8XDNb
qVaIrmQkwCWiL1wDEFnZVqpsa605yMi2mGVXaa9wQxpIi4jVeRMUPPDK9aCBi5wXneZmhA5fvWpo
7rdlseO6rtZYyQUP9+RwJDANaRBisz76ctIviuSml/m97xjMAY32RN1V194WXC1JDAG6tQIbAXOS
Bd43SE++eWJfu/K4s7j+aQ2QSx8qiFnavsKz7y5pso0uzt/ZL658Cr8+hY6yY3GhB9vW2Jf1qzEB
YLXaMHPdiVouwZctTDrtG8rG4mwjx1SsmILYPfAqkG+fVO9QIMucwrZvzKEZ19TuOY8cENdDIzSq
g4fqbW7q4yfxgfzlkkB7fddOYQSypuG1Ri/45vMwTCxQuX0Er4cSAhXCJLYyEtYp20jr3RfwlM3x
fx9fFodsaoRU+aQZiSF6OaDzGCjgZxWuC/vyGvBQP4PDGOAwTiJrx2WefVO7GoUQVECdTPhNhsYt
BpXTngO1MCWK+2ena4taZeu9xCpxs2/PyvUtrhNJaHxpq2RSody0llNCb2kcyJstiVINHZ6eo+7a
vWeG7xDCrEwXAoySAsn85GpFBIe1R/a9zROj7VGMfJZRVprT0Uqs3AejtnD8VhdKySoBVgbZENIR
TVpuKUzXS9NpTJRCd0QTdHZF48vRx03yE69oV9Q+oktObwoD/W7OPZEcujYfHk1kpLeMnt1hDJFG
sEW/oKLH/yz2Y7D7jnvz+29W0FRlmUuqlkgq3n+g39OPj+E/M0yxLCiDKp2bi/QOdgdjz8ppybWb
nTEyA+0A9gaKXpDUvxFWp1pYxPFKkRoK0zdz2N55UvoRxjH05tPe6wnMYJBkYQF1NL6Q1CE4Ujtm
/xsSzQqM0usS7xgNfdIF7yAKTbiIL5OjZpiJ3ywDVyLKY1TUKZvjgSkAXB60QwLPsn5Cl2x3JBV8
U31vGCPzYS6aBA2rXmsH9Hdybq08hEsA7sT+vo+Z2xkXf0Y+ZPqDaCbD8iVinq5WbH2Mqht7DOfB
H4iUiN87Mo/XRNMDbWzB+Fpx+sV815++1B6+K3xtVc7o6EbK5PuVy0OKPyWMrMjBf+f1clEw1pfa
Evx073CmXTyM2rfDMwUT7MKPa5+iVsF5tuFZd9G+IWZRjMb+37WTcLGPpkh4w0whkoFWlXJKF3zx
mRtmkTKdK9LfdlDtLlST/7i+N+Vip0apilYWkINFl9zQyNi3NhzBo63kf77d07EIo88bEQf0Ipsn
H6KOX5hjRKOjgPmKZ6ls2WttkzomhYlR7GhFVqjlF3vzaYAy64+stVoA9Fb+1ETr+/ZlWMWBUQSS
LQSvCnEQlwLQI6x/NOvCjBG1U/Umfp+v9AEqRnxfA+QwkBhGyryqPGAULUWWbLQwH/oH+tAeFQWm
JqCTPbu/dBw/wmJgIbLPgCFn4xeUwWlgx3DbUFmqenZtkSO8h9wf2jPgcLPmbprtwwVZpbJZgLu5
tsb3HF9k2SAH1+tAjVjXDg7VNT38gSK/qzO5D6iBZFhY9sAPF9kqgwGB9iaxqQmNdpE4fxxHYC51
WRg1TKLrMbwHTk2D1J8fyPWl+NpmqGor/eL2x857OctnxIAtjvzSgw4jFht2qip6qBLRJwd7L6S4
xB3U7O/LE6eUU8yxB0r+Ls5acAi3igHi6I2hcRhH1HLLPFw19N7wFPTGZTAMRSHXWi9u9GSEXisU
0zwsk486SCAF7Zma071afFV2t8AGZnvYZxQtiBJVYA6lXo6W5YDy9EVu27lF7Nv506N8Jjg9m22D
CN6/1HNg4S0i55jDgSY+InNLktmfmVq9M1oujHYyFCEdgYvAe9kAnLEBnz8HhYR2b283Nu0VG+pW
PfqgKhw09D1N9sriHCvY4gXOkCGuiicg+mNDd83igHZXe1MY1AFTKuH9fX6TFlKalvaZoHo6Zgal
5NkKz7b+IhVA9O+lbqGI1WSymvzYRUV4jnu+qI3TFZ0xxsOjiry8wO7TZeQwfIPsJulb0NbMzyN/
46Y7H8MrIbWoSQWnFdpiCONoJoRb9mRhHIKZ4J4buyqprLPoVBgkWp3qDnYTwTHqKZRDYflQWNC1
L3fpAw5Ctb5bty6evitJI3GxcQPZh4xDALsW61FwkZ0hHVKfxmNcou1cohgRhenq/sZ4P0ZwIwhL
Q5baxO+a5lPgIY6izC4vZ+vpTgzhInxWmsUtfBuEhnzP+3OT3h4mIuegsaeB418CxNX9Wy3zqF+v
Xb0mulu/17G5fzlxJR1rqM1X66A5uwBRSmHbkMfz3MjLrO8Tq5UFp/ssHot+1VBEafS+ry8K/rVU
ekFQtOk75r2cfx1Nokc3DkjpIVSvs+eOptrocWo5+0ZgdQy6KJvH7o085+GgED7p0Sem0uakXBe+
5n69xAn3IJLi82zSWGDEwbzegFitFWJvoQcL+YLVeTK/15mH81eGSeH5oVStpNxc6HO0dRnkTZCG
Yp9m+PgrI8dadcEQwKbdjF1FcbeqUeY6gq/xdv4xgbBNKiWfBINkApXGouo4Lc2+RqDCXcxe1uII
SDzcPBTl9UsNgSkcS+sIdqWB775k8zrner7hpodew7+lrpbCpauObNFRhOzBwO634JushU1JRsmy
c0sejbXTvv5bI9nFdakjLMdZ7meWpTOz85B6kpsNdwd/S8x2uNXQaOE1cHuLuYv9dKlKe7nXayAM
EK42epd5fTEk+SrnFXjA2E3at9TEBabb3DsnBucXO2k+Euazki5y/yTfEqnsXfzH+lbqV3H6RD4b
Et20StDYkCathdggOoGTWKDgywwVT5itmnYv1wbkecZMgY+Xjn3ptZP3EO0ID/DPVCaKn+rMa4DB
o1gAO1Ij7MiF8LwHPfRJJ/2IrTwvwmLt4jTOKp/SLW6c56Qge/RpKR9sckdrNJ3sZxJnLQLPTUuF
rXDQonSkliFN+NnDONnIkAPwOghFpVbDvXBB8e9SK30W4eZ0KOYv71dH99ZkHJqY5BtfvnkkQivq
oBwny2w9zGevnJL/C3kQcvfgKZ9JVc3ILEmc567IXfzC5pfReF366UVbxNt8vV8huE41xqBxz+9L
rinbJy+cxWwLXxEJcuHx7QRhjbqzCwBaBf9h6FSYxQF+u4I6NiCHtc/4J4X9xmqD+46XSE/DJfmZ
+VGxil7TdaUVk4Gq8IGp396DDW9XbH9AeFl+s+hDVbzgNNq3J+xzhNR5FrYdJE54I8McMRDNKGyG
feB+Fx+h0ic12SDpS/9yNP6pRoNycDwz23ziocoQ/4fBgMO7rcKrj2McvVQYVMLI9sLY6pG6tauZ
rAeCa3ah2Ok/mlNOXp2Itmcnd4cD8HCxdcxdlUe90FBoz17Z1nbOwSFeuoiAVHKPsjes+ihbYp+Y
NLwWKN3hChLuvHXbJ4l778YGQrTEHc3fFzLOVqf3c2J1ugfDwz5b7OzLFjpgqPNi+ULYn6A2eL6e
y5vhfulyMVn2HtyvkOIC77LXEXYiYTN7300XFzVdl9AumkVmRKGPQqqzcFyNlryXL1nFhvvU8+2F
mTXoqeEgXRpsoZPN/TEUG28Rada/GYB1Xft+oq8Vw6EDgdUGXm4Rd/YuHL5cR/Kl21FsYQizb/8W
QISw4SYgXG20J8ftyTtQIbDaHZRVrK/X5AcnWjuoOjzwrTzWbteR9X3Mo/+TcLxFjdRkOONrMRkg
2Xk32GySQsdNPkb6gVJ/+TrSlwVUaUMdgq2zjAtC6Rtwv5D/eTxrTBKrK3I0C4VXmS3UovtH6z/m
Y/MqjuiYxPCXmiJhhZaHMJVmpBPgAPDKu9aVjbh07kWIbX5ZPHiwPi3BrKZS/PUW+LUK6Hl4Zo9T
TbtfGopkE35jRqwTVrbH/c6BXlwKpq00zmWkqAeMdyW8oWLQM9GQsIx/ssh0ab5oTCKCFS3L7pqP
R3LIxYpGQR3CBWGNcLHwZk7qJDQjhdZ3S9WmaXeRAy75wQ/N7xDLOdUrK6UfQinb6CE77BY1Cy7h
lf5JBx8IYHdbxX3NGm2r3s+7OhYEZ9NzqVImLw4RYsX8StxA2+MBvGYvEhJix/KImqxvk7wnTsks
bXGnVuv6T5BU5Kc0ewPFtvkhyUbbP8YRNWIUiF7aHtOdNdMfG0Pn4yUqU4AsDzVgkXeY4loJwKEE
D7flLJr8FiOwC6IwQdbX2PpqJb3BhmCJ81d9T29aLJo73TofkQxnxBesbFSXF90mciujTQC7ghet
pKpKvrQvcPExG8qEuebFl66kZMr/XWPMaS/xAADVmCD7vr4erJWtjx7pvWcgLm+GeVfRx087Az9T
Gq1zUeWq1usVwQCqaYORSUF5eXmiuCvJIQ0x4GYAjLzmSxA/QKrqWUeWVSDmevU4RjXKEupE6jrm
mSd/dG12rEv1u27vMvG48UzElmiSKWrwaJpyoti0d3PuQJLgwpDbMIgJaFbW5cRhzpRd6hQ0R8um
GlAwZUJBHbVOzoXVT4cEqLTCCR2JVy499HWHh/TJ/NLzUKUun6a6AGzch03UpUsgpQs/jEOoq/Qg
iIPtl6GX7eXMpTHZIVB1aFr5dUQY1MExoge1nsZ0tHUQ/Y2bGCiiWCotmMo40Ep3kJWu6khl+4jZ
/iQ1CprjnSSS+WbVlRcTVY1OygRncELTpNMXbDfTXtPw+wc+2eGy1ZP1g4fXAcxBf7CxrBE99Ygo
kUxI8yok8DIcIiTmQqUtKx0ly38YWZj+vhukmkL1vs7SwhYDPGd38b0m5TJKP7KAQ3o4cb6wslCs
nvgoJi1Ams2SJIRjqkbwebhoipgeH/DGbk3kRhgoljk2BMv2VGUdviVGleg5sBEj3lTp9MfIC3Fv
kNelfhxMY9hQPp6dHAYPUgbPnFhBA+7tcTtmkmN/HRjCNdV/lbt/796T+RQ2kNnTqECz9Fk+5yjl
vNQgVsxewrDUYSi0ptLiueIwXSWPWfdEbUfbRj8mG8alCcrNhoBj6iurEz8FmLxkoV28m6LQPejE
G27vHSJiVEwuhZVsbcLnw3We8FWELSA7V21g+0koSy4YSPBUCNLmBhHWORTG1S3ibeAPPJm1oU6w
z+A8Vp7wZHsf/58cfOyoze2EZIotqTStN4p1+GPLYNrfqvGwUWLwreVpS1nhrrSqjUyaWLvMsYT7
YKtv02EQvgB72b1FYRNI47lGXY1yoO+70Ds0q4BRbhp8/CZ6+pNT7HZh2z8GBXQU9EN24LLLOzeu
5S5xO+AbeDsfvE06+yt2A0Xu8LQbYRqknolhX0TU5BogFNW3FaPiUX13lqoFCqRJefPyQ2teteit
RheMYNXcfKQudlgEEtTF42ifb6ghiPFs59hT6/mAwBZRilb09JLH0kpQgL0F9J0h0WeVMsK4Lxf/
R5gnLfW4hA0n1Wev/bLkEeK2QCmVjsYSR9RZCkt63X/rWaz9UyU07FgHcufPHO5gvxHIcZw4qKPk
U/n7eBcvncIOcHMyaFQ0WX6yjA1QsAew6mtFnthA7ycUnjoRYkWeyFk3p+6m1csUN3LU4pLvUb4x
p+oinAEd+Z8Ae3J+VvCYtlXdyZZ4Ndz/ao9S0BnXzEu4W5SVkc4EAfMi2k9QzrfFVKf7oj1cjkF0
gnyivnElScg0OEHLUvJ9gHrQYEaRPRiS8ygp+CT5H2uYIKlv9E9R8KHL/ofDKhOqB6FiQU+c6nzP
1Z9oy5b1n8trisnbr4cjZ55wPGi0AzM99xnIppUUpONLPNtBzEmqikjyXxnz/mCotgAiHXKmvcta
bYY42ASKeS6alVMOGkzb0xRZV2vtvQDh53m0I2+4ZvR/uXd41eA9DHDx0YqH+n1tq+B8TC9y2xtY
OK7e1/8+9BYaQKHGOAWvMojjttSjcX+9s+jP519x1ucYDSEw4v/JcdRvf1vAqVPeofam5ancqzVo
VTs96b7Bo7hPxVd3dbqJbVIks20pMpgfTIAq2fhjcaIcKG0sFTS0IDW9b9u/w0FBWaiBI9oPIm1h
LbY1xm4Dq3TW9fOSki/FLK3RYB6X3P+plULq3qIa3AEanRaN1HHo/vJMNBqRFL9B4F2RotqbxRmN
BPqM65p0xlAKMGwsYZgAdWKU3Q+q9qsInDuiwM82PzEFdsaMI3WvTw1aF5/lRD9QYJEHszLWE5Ju
XL8exeYOaxjCIwkKafMwmXC32w3ht+zsRxVC/wkCoRhhufgbWD2tAk0YOy5P3lqZ7uwRNWzHUrTt
vcm9vY58GzdAtSMjzjMsD3MGD2ufJZGoriJv383HfyZS5qvZS2beqM6GUU2ODrJ/8F1BjAQUR21c
gAtYpXbIkZr4Ye2g3Kz4IC7tmhEV2wQrdWsFO8bUV495IfqEk049IyvfQbYkq1z6oEFN5TyiZgu/
0gK4nLJs284S4UoNNSo7d1iJsVfRrsDWaFAJzLxU156ngMsa6KvuwIfzOX3sHVHzKYH/StqqnyZn
TeniE7DjRNtMndk+/APxMZVdN6W+DjlVXAecXNYUmok/GWiySycxHjp+NDClG5GH0UYCG/K6RbfI
k9cEvn8BTUOX5VdnVtP2vToBY8Idbyo+HGA8TgGZAMa3ElodeGSLcbF5mPXjMKbb7yeN4hsizqNs
oAsg1yUSLGfceXGAKNCeLVkiE0hTNvlkhb5s/U/MzEiZpAyDpp8RHWsqXwRAdQ3582OUmaWaiPnZ
6+a8AJJEqnC7SnskRwY72OuRvfIVYfZnHQp0x4x3HEvk0Ec8Gir7LnEsNOSd3cbvPBGLuP0wQ035
fEc7tcJ01s8a+WiRGPhCvvD/riGUjtv1JLTvccI0UwmDrLwEMmG51mDIE3Rw/M58OUTrT+HramKB
fLi3mlpZBIidmSHuVdVhaIWD6qXg9XErBpfu55Wr5dE5b5A97DU40mnYwXol47uf6QoleOCyrb79
fTYvMwczBC9hAbC/gfuqUfBwsE6iKR78aM1Mjqax5hE88vO/KwQrhX4h2x9dHzNE80bJSmnVtZnP
Jt2HPT6gytsiG7e5Eg1OmDFbO94swYSfOLdGwX+P6tRr+LKnENWyhnnNf5ed50XlNwf84sCdCMNA
2PCH3NsqzVA8uqNPwzMuFW2AdA0zl/bij4pP7YT+tbLYoe/nemIM/YpAZ6LyWVxTIAElhaAWiUZ6
4oOoWcGiFJZJY9IquxivJXBQtcWWsrZoLHHRvWkKnbKVLWLa8l07Qw9zzKs7u5cY+DRE4xnWPeac
1EYXJ0RspKHvA+O5wlu1geD1LJ2aL6CRov93xTZsNfsoKmYmRADXLyBn/cCDxHuFjNPvgLZMHkgX
VAMdiMJwmFODFvlwqUrpWu+K23V/47cw9YaqMtOknnwkiw5oOz1wcPP+K2lwDvD4yhwh7H7rh/j8
JgEtA06rCt2/EMS/z/jF6shEnoQ1bGCPbmUUxe42hhS7AN0LJ/0KfOjmjU3+pOOEuaWrP4+2qIea
BVH91OM3Rez7Rht08ZmNNlafPmNy7wUI3Mx39vJiZNxzjBVyZRc5Q8df+0eg0t27g4LdKQ2TF6Li
jbslF/7txG4DzUSuQ3eO8eNjXSuKPUj8WpKpJM8Zku7TqKNqLSiz2vchegXU7SFMxp0/7PxLvMCa
5O3lUiSi8bTsDMEL2dC2U0uQgw4dAThcy03yqxtqcognY2FgmOvN7tMCu/jCdnpqQ3yG5slLZAC+
1Tn/LEVX/A/ieMqYRh7GLb0CoQ47hw3HNA50b+XBHp2kWErxpTecJ7Sfyrle8Tub3byFde8vnZge
HRc8qC7FkLAm014K9y2ugqAOvGYa8Ixp8wgDg4rTQXO71F8NG740Nnge4MbtBDszKJgQqux2FnRD
bmZnSNzNVexhcceo1FvxSn6uF16Qx5R31eyJHysGAAsFc+qmvSiuUkEXAHnnwKAeOYcW1vX/zpTT
hEt/IQg6xO3f0GsPF6HF10kd7xDEGa8Mrne8nGWNaLXijqEe2pWHQ0WPhnzqUcgJ5pb4h4/e+QM7
Op+jXj6/xCrVFKPAMYAoF4GYCLQ6V+96PO4rgiVel7vQP7PaBih31FPaqv/nQy+qJ/szwSm4fZXZ
OTNvcuEuDGhgp7Cgbaa9GjU0VVawJXxYx2f1S2hCSb9M6sbzHwC1k4E3N7rlrLkS0B4a+gex/OJP
eZPDZ/cWsOVEvizkG+Lg0FubiVd+YYoxwt3KvIxkt0tV3EOx4Lh3Dk44RLirH/vBsqwH3OUgGc0B
FUIcb4XwZfcz+PqEFavHUkDExuwd7ruDSFU0wC02OyDE8RxFwVR6ar1qYT3oHXr5KSv7gRju/Bo6
fwwje3mbwzTLW1jcK2bza8DpzkyiP5Oj2WRa6+qTaN3g5OxessA1fcT2i5IBuCXLqYoafISW3cne
dQGR7D2lMAojjFEL/FUT0Um2Qc9YeZSjTeOXv1WSRqraB3Rh9h01E/EI6FX3L4xi45jQCnW0C540
HfM2aZChN3szGlsCY0E6m56S+86jOUSjoFTYY9dnLInSj0a57KUiXUeIsQKSPrRThaQgrWxDdBrC
mOpQ7qvQKQ326XQ4wJPuUfJnSEFcAlovD24+PGxCYzRVUG4X9SQJhXkP4qTA8FYy7rUZpXIzP7Se
OUQ1FmSl/YxvM+1A+0n1lcCCTT85FFHp8//F0xg5/70rL32ts0utX7ixseMdMFQx8mXHFNquVzTZ
Lz9cqagjcRNfb2ARogLjDcBEgmzW2V7nmlU3EGu5pX9t1vq1vyU4WaC6Jy9QriSEGIjqZudH7qZH
SMr+2bAOzHm5OzR6hvjvmUetq6vdqOaQXZcwrN7h2jn8wgSStkntodnSWGh8i7jfwG5ipAuvQ4Fo
iJAo1cEjcm1QUUvT7kejK2wyAXG0iucYrWcGp6QK4WZvPYdSVlQNCY8nixQ/h/mhREqdzg0eo7X4
b+6lR4+9mqu48l8Z3Lj9aUxE4XXDBRVxHOLlWwlqyOsfy+olTS8yfMu9mDoFohSeqHWwWzeOPMRt
XxlUXys5z3g8BivpZPLs3yMylytMKGdMOrrZQcKej6mMpukPJCgDSDjxLbltgjebIJhACv/FYdex
gC4nr3gUZbZAmyJ9M4ITRrj8tdaglI/bdgsfIKy2Y48X3h0/7BgEnAgIFIrt/nscCgCblRKjjUjW
j8/Zvegj8MUU+eKAjYlolbMvVXwXs97HCFQPFnS1g802DjXSA8tmzufkG+6AA9fEZZvRGacUFu3s
E6539bYYTES60DOnWmB6Mu24LeQxId9H9vVYpN+vgv1A7QIGb4qeKPKDZMgV55qLYGAxihem23DP
xUStQxFmQ2rHEwP88EHv8eS4ZwSB8g6+VAWOYtdXtqzCIcYg8vlPBLZqeyy8Bxtk8g9BEG3Nllmi
CSWvJZ5O3VIeyl7V19heq0Q47NgiDK5lk5FPBErDIWAfJ44hgi+1I+mSSChngpjGjELGO3tLEH8b
ojTBa8CjHZNyHWZvlWZm0qL+FTi/s6fka3Ug5PBQGS3o1cuXTPGMMghq/EIBiQTeBdQbaxQylMoS
VmkGbxftXMHHpfovZMdF01AsMjJTAEhIDmFe7WSv63Yu/CWapTzNEbdYkHJV2Z+Oaa7SZzDoDctb
yfzNfizbtMKjXF6xR2o8g2ki9c/FOAeZpg5XHqhhSkQKkp+ERF5R7eCfoWvaaApJvWsOQoopI5B6
VHxA/i+ZkezIvZW9aizwbGqtnUmXfoCWQOe8A2x8bJ3SZ67e1KOIesBXHU03gzqGvZpcQNfkVSj/
7CszlX94qF5URFBgByeiiYqI5LoHDU4UTQBSlxs3tDBKiK64nKKw4+37W/q19oT4z0+imnZ5jSgs
3/MRDSibcPcL+m4z9ZyUGCbe9H7qpfnwN1c9eCdtf9o6PDakSHLYA70qDOCi/ASdunaNccx1iMtn
A1nC/UF5j2BMtO1lw131rOek3uOX61P1p+kQek/8KzoJgfQ1Yd6HT4PzrgPFUdotrOrWgS5fY7tm
zXAybPAHgZZQ5cQdDET7+2Qcba4b1Ul+CoTss1QRU2KR2c2WVnixVisNMDoue8ydhYaU4ZMMjCrb
9EXMv5DW2fx2x3cf0nGPvWRJBqFHF8cq6X6hGY6dbnKPcHpNNO/eSdPiQ5PPgt4vp+/Y7VmTzBpI
KVh/aCoGsucEw3pAf9HPWCC+lHB1Np0lkEP74z09YKSirSl0GZck9lJMpvkrLRKYDRBdq8nrPUcL
R1+2Pf9akV4dTq4jwuoKP4onc1IWsdJv2XtVIPTuhxN2Q5zVaoNkrXIuO/0+IMJjvYU7Xd7rUYiY
q75vOgquI0mKp+u8sFa9j4+/2tstLEyTpgxiU4mKbTdkYnBtxqXxyt4OkkbS8IrXOAjyxxnDr0hp
SHSCWG9tEmXcP/ADsE3KOd4rpul8zosSHmWjFrqfvKj4YiB44KvKP6n4NmGfbna10RcxZWUDRKok
3n6cr+2NLlBbmtQJL0lGZ2qC7u8UPjgi5Uf6a0eyVkF3pFOISrsnka/5VEGeMpuPNFm4tIT5gQ48
NOIPfi/Sdqg4CykbATC1rfTi202vv7bECYWkme/46MdOar/Ub243xnRpZzfGgZTN9QzCYnFTP0XK
90jqIIN5c/zNu4EaKeRI7rCoNguBT2grLLEJ7OyJT26r7nqAiEW4qfffif+nHquC/7oMoLjsutCS
OQsJplQknXRPbZtg6XJc1UJ0pYTJU9PvrVieU4N5x0Gwl8Mhpm4UTa7CYUUNrmlDkVYfxdl2OdzF
qFCO8/ihSL8Vsw29tDz6//AoEUkaLHIIjFvIFWgFYzgJPBnTse93m6EQ3u5xRSI9FLpFeVq8rEUn
g9qSosgWqs/C4p9YD21NVW5PZL/c7vGH228TCdH60l4eTfPS547oJZ/NzfdWtgJHXECc84NwQmSR
/KOy56mWj0JDtWb8U1P4fI0UQl2HfDjmSGQC6Ad2ysNH088m3xnQPSaDoNqpFFI7rYR4npnCMQcM
79E6iTZo2rHo4iLhAWMWa+tqb1ZyznO5zbd9TkkagvlkWWqVk04KShaQjfsOaZyKffzWQtDiMKMY
66eJL2dwHcCLrnBrJPGUVcjykFTCRrQPqrJEEnHLxC5uiG9kNFu2rYwUBdvZM+UNYDupGtgjqsq/
wjUKvfWtzUvRK0+O/HsZaWytN9Akn1YGPAaLDLXEkQ1jrbIfiknoQNTQaWeTeOW3aZwvTDabPMdO
r+/hsBcRCNATSR3mbczX+T3j5UTvnpiCDCwckC1dDaWU34TWKMGkBdPz2ENC5eDPcXB/eg6tDTqa
c/w4cdfxgEKcpHk/BEoL8bXzdzoKL8VBlLtwR68h1e0lSOEcF+PFcjk1DFq8kFUl0JfrE/GA6Gqt
hhSPlWu/XbusAuXgUMBoNc0lDr+ZOVJjFD0hkjHbO+MKq3a9bvfqrAaXuGUUfPKemaxCRRZvjb90
N9IPHsmwd4jIy7SHKdV9vOETd5I1+eYwDeioSaOLJqjs6oHgSSpIBSr/qlXWPY0jOAd/5INlh4jo
noyK4vzQDpJ2txsBGhZDeut+z6IkW7QlvMpCukdZh+lYYH2TQmmqEbqBvWaYeu+CSgYrtjfKecIb
QR1LtBBGWlbgfdMF8eMw58yL72vRvgRm6O0ovPemFHQpkZt4v3CShXXi+ZEZDcCIBd9cRotV4kb3
2uLVluL0LwGm4Nni/l6tpyniGZ8II0BqQys1E2ynQyCSTEsTKUyZULSauvs94G6Pha6cNV/Y60gf
2ulyR1KTPM1VM/caRKlLYatSBgI4thkjyq26t7D8+HyNJW6mechyQu9C9mzCjixW09R9b+aH4ghS
OaMm6ayED4xM7VQ5p1BOvttAGYhfxx2gnjgPbIh6mjYh4D8eY692jxJV8GkprYx2vEewDsFUOfw0
HVkFMC5CmYnfs5g2uDSOi2f6KdlsGRL/jouePN0AM+Ks0axr1hqmxYRn21xFsqXlRpkMiADRxCLg
YKnH5VFOEAUIxhMU7INKALu+vZmoQV7ifNOa3qszjiOILdu3xlUyFchG/lV/ucwR9ZB1hZrJD3IN
8QHYWzK07ZtSuLpvqmDfZsUUd/ks/zEfkAcB4arvtsUNHkfd+0eYPI3MytmR+TilQWEXOFqgBq21
K2iVlkSVGjB8m06479gl5iG2z359Rw2lB1Nn8WLWiIHeE0zoHSlIyimsMu5jwnE6EKeVo5cE3tA2
uKePBXAi7Fdh5iN8k+AeqLJY8h6RojdzJH5CfKaSmWm3f/xv22aILhbs1n+pDyRQsjsn2v0qPJJa
3ZUG06IQHgMkIbXpCTyq7WmnpquR2R/aCEZ2BU50zezWemXADWbrgR0ZCITxZtI2YNZ8hQpy2hcx
L3PIaxAQSFKwvRxIhKZ6umii0MQFl/TuxNdJB3iE/HmPR/cuqTtUQLNOvuZQSSZ0ifnY/q+vPB14
wx5QGJK+Ryw9Gy+q6+s3m04/2Nnm56RWF23cbS07kLPOgUX4Iq+p2Rtm0uWE+Hy5qc63hI/IgnE6
go7h3/A3hxaAlirkKwBrkgtZcAB68onh7vcYe7b+hHcs7hI/Mf+kzfw4vcXVOiPI3z8LVFZ91IcB
VCBknMzjQ+4nIWZWQyGL219hgl6y0267pB39WsSkqqXcujT8feJn0n+bcl5qegF5dE+N22Mjki4Y
4MJcY5r5M/SiwrJw6hKmhM3In5G924noprXPrlDJKBlzvqIP0txdQVYO8RGX4SicAe/ZDiccXNeI
xIc9xDGm2CxaRxTjF8iaSF231bqBEBn6v5cqMpmiiDtAA0wIR1BN2sFPrrYx4MRjIeExOKZlyLK8
r+ikeP0CQqJKB+qhi/kugVADLlz+hy2LD1wNLWmzPtVGkeKfnUWK7pxvDa2+jMG6eoWbZXayu93D
iV32IsQszMTMHKsIuku2HId0j3Q53qE97ThM/S5VhThmEFgTV8E6T0zKOVeN8H2QIwWxu1tHd+fa
Thsjbe/0EMmHrv8QkNlXLjcbfQ090cZgvQqwlEHO1GolrC+zVdng86sejRjws3TKfeJcKqKrgoeH
I3Kd11QDj/HwyR5T0ix684p6+HLjv93ZhKc6fBLKai8XdWeCmc++kH7viL6RMBZU1B//dCXi1o8J
3qlmU+0BGn/HI/6NMAdXalEv6zH/+354JJ4x72nlwb1ZzqWm4dETNr8QRvg/YqFiPX2oMqKRLcUZ
5xBxw03hitCjNPn7yjeDj6AXjToKCVWko4vMVM5lmWbac71mJgPIzazY421dNPPg0ZekpuVVWsk9
8+mri7/F7bet9jhFrnnZp4QteYs9gwVy7T6189zRXprz5yQXIXVK7W18G+/reYCYJ6F/dhCtskY8
mP1ZUde68dYyrYxL7CVVp32Mof/uzVDDvN9E9eUOxQjjRF7aMqPs1toCjHwmLAoBMF9bWsWxgtMv
BLZK+f2SsCL4tVefH1Zg+OCMd9cMMSXk9B8O6ZCgn/PQBi+pUrGTF9YpDiGkBA65Wqbd5nmxrlpr
zsLV2FyIuGJo51tXnK+3VC0XdgrZrenxck15pn83NjHA2YipBdFrz1bqca89X3LlkhlQN+eJD/GT
vnNyw80UhEcpyEApKIjBVC2jUETDeMTM0CmPkwCHGb/wAzFEjskowV7a/YSYNpYLSzjK+Zt3+V+z
3zYdk42zoeuf5J8LsbDIPjtCB878juuJMPQV5KoJuOVavJdEYH0f0Ge5zSDMyn4J0ZbiIX/+jpA/
YJxV/vq1cknVcks7JNOuc/KSQ6jQ0wDD+/7bFLky1EWGFYNr7AUJSTBMH0GtnZ7O/MC/OdYbLmBj
j81/zxlrKDS3GT00rNa4VroNL2Jf50mwQ4Xl2ZXtX9khSFJQgl39YqX/kSsm4TW0nBUnldLdnCoK
gj8JPsOAceGGWA+lmpEz1tO5/OQd6D6PT0YENgT0XokICmFP8ynBzJQN4sbG3jpeq90ouCDC8XIs
cF8OY62bCWlA0pi2nzCWtZOsEDs2qknMj6Qrkwg1zrxH4v/7pBVNYmjBWY4d44Tvz01R9qmnKp5Z
O8Gbqq3vhHR0DbWGGh7tGKo9WVeyJrcQt6yHPcqbKCLf0oDgDEb1n9Nd4CtEF1HKJSHAZewRHQpR
c6O8xfHPyc+Oo8YHpUBOb/i8Bbf/9nQ3gL4ayR2xUDXdgjxL5S/G769kcb4aPmNf4kKTs6ROqXmq
zI64ah+y4CGieX7jsNoTuyVeeOGb03tm0El8nF7omXlRnKntuu5qocjvsF7gE82WFrg/zlTTuXfi
4NIiZhO9mGctU+xIBa822F+MqwDZkztb2HiQVnj4jTy5twKHEzAVSX8cnIgYVDHeEFSwt7EZOv8X
CqQl/4RpsHeNd0ZjBwUE+qwlg7hJYPgjwkCwSjgRIZSD8Ay4jyTQ7mFAT8CnejPf1oSw2+Am+JXt
2USDOphMsxiNW1lDjzYCvunp+UmkIfuHmDRJkn9RPkkj7quxi/0ub5GnhFkCP+tQRx1EBLlAnnZC
B0YnTDhbYCzhUqDE6ef81QYYGwEvNz8BhU+zSphxWHIuEhfUW6pIGytbkxnFlqj0Kib1MQrOdCYw
uz+2B+IXmw9nrihZIC1rRUpCd5dkZZj40WMMAibmwj4S0VOtlHE9CZiIXpFov6kTvQQgSH0Nldve
kRPHIWKBquru3+wOM1BDmzOGPoSUfCl68oqy5ulTjmakBBFQ+W8ILlyj3/kJLeDVr+sD5mR65A1S
gNzT31SU6uLmhfreVNM7bgEFaei0i1wViv8hEyGNCEm/5HxB2f7/DtzWuXcc8NdEN5o7iGcQr1la
P0zUbztR7ijVBJkuxTmMXs3LYfNr0BwkDR8leI0oIRctWuFU+u6nTvYLrHg+9lxHo5tnDyA1T4+v
QHZ/HLgsomTkU9ZbaMQUaKp5C3p/FZPOhe28CA/O4PcarWJD/hDNiuH0tvtKCRihubhOxfJNS44t
paBlAR5ZFAe5tQzm02/V53vYSo0dD32t25s4ja0UNItCB6e75mbP/GQ5W99BkTQD8VD28FalN1K4
RGdcQc2h4dzR8aSYBXCFX1u3NhwcD9qLhPgjsru5tW3kalTLckt3ob4G/qBK5B0W4iApG9ARkqpv
LwmLl/OR0iXpY03I7rT7TewkrR3REH6UD3ZclNJdfv4d2IYB4MKpx9ObEBb9iAmGeL9pv1uPil73
BaPBT3tiReYC/SuaeyZ1uEPqxxRxa+QhhoM1KOAzyu6Fzt8AU33MP5Acp6G7Gzrj3IXC8S6g7NIw
f/KUtgjX1fhM9Xp+u3ujnN6ms+dsCKTOAnJPHAwAYr/19tt2rsmr9yHcB18JkpeF7C6p9xfmXyhB
PFQxvHhuk09BC8hYl6ZrcpYHQauid48LrX05/bZn9wac927jVCMjfFtVVOezkBjIzWf4vAbr4xnX
Ji596itBf1iOQRqEE4hj4AhPHpfQLdwQBPimG8zsIPf1C0gK8gT2RDVOOMbuHjviqrkw42/eLDcJ
gIkP+DW5HGS2aE4c+393iSHt/f/tdtA455fH6LCtRBeWYmuCJ7xt9N6JiWDEu2YYgc5UddTL+VeV
0R8xnAThahxYuYOZJps8wOrlfooEyymJ6QLPwcPra5yHYFwTe4PlW4DdPGscUlEAIw/qnFxwq5+I
GkS6Pu7QcR2RxuHgsjx2qe7znpkcP5S6kWfhNj8fuXQrTqQL+0ehH0+xaq1mKXlXA8NlXwHa/iHZ
ZHJcbNsOLsBXHYbuH0sOM23wPdAYlMp+/MR40nCHtjFDtutKgfNgLVPzOjusf4vqm6yb8cOS5VFk
RJinZn3C7Cd1QhvM92bUv5d1uvybQVMXJMX5l65oTBijctA0t6N2wytkqmdzJrNlw/TXVoeACX4t
53Sq+PjTwhrRkD2bS5B0wvVNFqPSuuKIBktIaZgwVP3qAv+4oAAZOhp5MyXXZZOlwwyok5TFNkiP
wrXWeAMbuhFn+V1pm8oYnj//Ewz4/zaKOKbE9UoZSWgmnHnMbUEd7/gKwAoF3fRwy3Mh30qKdQWe
r9lVoee30uoHodEr/v2AuwOygGi1XU2lhmRZXHSV/P9p9h8KyYGVSBno9Py2t9ICWYD+PFtlv9v0
FHo+vOx8hxBkFrweNJxBr+9ST2VPNXiOmSmV6fZEruOiY37Y7A3y5lSO0kt+OAREZUraGKFq/LvS
8K+Lb6J2OtIOCLwPRjLt3E2hKi1q2dcarNJR5/e5d4nDu9gDzZ2Qc3es/AJK4C9NM93Tz3F9pR3C
TPL8n4+xWRmT4uE+gKH8E1muoUqWsAzY+MVE7G2zIRTBploxFo8lfZZxG49Ngykg+4kSligqtv46
B4VnOV/pASk5hkdww0ZOQIlzN/hM0AeDkDG685IiYuWY/HCMikA50bOFKSXXc0A6PYWuDIGek8rU
yRrmK6hPaSQ+gfxeI9BV7mneZEVqrBbmrRkulvQ4E9Jcp1wskXnjdBB9IuT4h58dJz5CH9ri+mpA
oPHCQVpMmw5dcZOzNBRxnPjVMgsblHoS9JabnlxhWrxDOQV4YFYGjc05Q6w0eH6khjuaEPlzYFCg
+035OkSHx3xyOoS2aofvylrV7U+s9SHRfQeqjwUfo2cLemTBh6vrdPe/zuJLVBZJX3Woy1xuVlA+
lSBs40Lq+2dz7/ivkYGLAEHJqZ4AuTEepgDQn37KTtfQSlFOcsmg+VCiGSyzmuBkT+hqsY7tnIuO
k13Sravb59YhqXm931HaevvGphWgoD0GOvTUoquzUt5z8KgUQj/PAAjkrk37ukAem1n/NT3oVmV4
WqV/8gPcClF/IPgRt/mVYLutBOdm2o+8C/KlbGZeHVco0iIAHKuJy45X2k6ib2u82nd7B7w9rpoK
2beOWzsdHwXllZxH8Jxv9B1XGnj+8EIuCBryL8cU/bQOxsooHwhcNKXYSQBp4s6ZWmYy1VtGMVeq
KmI70vHR9Ls1Rxah+sn5MGM+h7i2trs0d5JwGdTspXtxFUxf50n1bySi8yyU8+qk/LB5+k4/tD0C
2iVI9c94byyX0Otw4o1W2Ron6DwMx97E4XDaZsYyI4AnVL87YZ3yV6IkBtRx9YfB0doDSRHllpDx
BohbFmR92yVs797X4/i2a+P++vWdXtvgu5pZSMuyfFKen8n/dBOpv+DVQRm4gvHfGQky79/Er9nM
8xic7rNVp4cZ7d4Kos1QqYtuKox+9f/gDAJRZ23TTdwnQfM5CZHMmbH6DggPlgpiW9FKjRcxNXmH
banPwixSxmhgwKV2iCqlA9IxGA2JWj0o73ozKU3G1lm1BlLHVs+o1ddMDMPhF0i6OWyr/LRVtJNq
cg5VVTzWVR+BLDowMtsQtz+mZbyj0srXYBVrx8s4hA6CbWIAYpIHICdhGgqhpD6ApcUL6pKcta5d
10XFtViwoAdPL8hQ6i74ypjKLhkgdbKlfzUF3vHg7+9XlN94nmQPRNhgM31Y7CRvcrrrxM3XA/+i
f3NAdAdS21pze5N3w8fma5sbQuZSGYGoQKZEcT/W4polrA0rovmC+1nZkwvBMNGZezdGvjKRVGvt
tzNWW4aqeA9e3YpYPoF4tOxyCbV5K2FsDZmOXHKHrX8PA+hqdZODm6zAB+xt/YnvxwVKJK1pMJXj
CRRXbCWU8nCccwdIjjw/+pzSm7gZdiE9DDRRxqg/rCrxK4WM+vRkzx97bjR79CL4lTCc+zeiFfxp
1Ehv5KJwg6zOWczEaXUBwtmFKnk9FA9jkXkKuPtEX+Qe8xlJ/5ZubHtRAOBQnAvbvJ1MdV5TK4cb
lbmx0k69HHoFDtkCvSRvlaEnTm3I3+YNFF4uhH8z1SSgvKDvcP9ziG7FkRJ++s0tYxBv9BKoCNhS
O8SN3g2GH63u4Iz7ICKWnk9aoSPUdvx3iAKx6o5ObmU84C5PTIKGc1wfQmbS2o1e3faCxL7xV4dW
Shf19wv/hp13k2vh6OyjXXjQyjk6og1UhJihCIOCCNy+ZnRESYiPHqlXUQ0Wz+Ki8ZpF25pQXIgc
gTFiGonmXFdZ52qD9iI/tb6CyPrOUA4iQotwrgqzX/EebDniSk6ADVi5w8zz2NHlCZlTMCPQx5S8
mMM5GOHapv6iLJOdQMhOSCCjwVkMnsG7gg5tnOFq5in4Zr++gMZ3oZdvXxpRhxwWYYnExk86Bpsv
zi0tzSkahT/rVh6wXNJNYq8edUWU1ACGbXnI/ogS3OphIk8mixm/3DJwUysFOPP4YPb6Q8EHGLZt
r2rISlR9qrJwlSo3I0Y2b2C8ErlgQHUopVkaCyBYdUiFPjBtDPchAwWBIhePuOWVj/YGfp9gv6Xz
HIDjuXV29kw51PIjUvpfCiXgvgQTRQv+vnT5U2edJxOAjpti/kZOo7f5fMLUMi0WzObUKENQFBTt
tk0IvtXxmUSkLV0BjhaniU4Ahle9HPLiQogPbPYrMNVg7wD+NFpQQtZHgYF2Igv4HkVqCl6lmGF6
Zr96BQMcJQTeMDxx8W412jOEulpxS6xdlcTtGAnFmxWE/RDJJRNzp9O/ypcHWrjJ48HXEQPtZ1b2
RT2ky9CjJot4n9qIimP0hiZJ/bC9W3onjvS2e1N7Xt9//OVgvyo4Y4/gd5DnpizPU6VKUHHjwGPg
2zgXCJcfpN1cLN0qdxcNmP+opWnp1sgJI9Ve5YcQnkW3zQ74D2GwftD9ZnIMvCHw6VJylDZ0TxRc
YnUju/0+g/jSjy4LdkM5cMzdy9jKnCEj+JvWdYyAmfteHgRkvYhRnSXtx771kkWhcmiwzw72AFo8
VEF0/0ICXh0mdD166BxjZe8/ijeaMnr+zL6cdskE3aLOv4TWXMXEeTsrlXIl0NByTCES25MSSy+y
sd12+6znoaKcbOYg+c4NGahucNNGkr2BbEKQWFkP42DqdWMsBW27EFb1fD5ZgaEcyFN43e0jyZo0
PFcytUqdEnqtMMoChEh7WC28WFwfB/PVwpr6+IgA3NJu4JV9gwOdK/m3SffFgq9JYuVTkRR8JOsX
GiFCxFogiXoHjml7AUYww+oFnrQwSUYWJvWhtkzjsupyuy6vbHzFi2x4HfDPgRvC0qcSkGLn5eG1
WDgV5g3ktH45x46iqxixe5T3W7LqhK+ji/ki4Y0Xm00266FZLn8IDjZzC4Jb6c5iFo67DxVdGlfu
exOAyngmynVlhmWGAUZEEskeAyc7qH/MU8ccoqjNMWa5OUFBSNHfjRWDOsEiB6vNv32sxgwrMDf7
e4BhV5gP9o2bO1jSt/KBTafgZaAYs0pvIt5OsTldEjowuSn7nCBnAMHSGf9S2Qzv5yqcnhBRtG7W
d0dLJpyKQM3Ll3c3BXr82o9oM2/q4Of/u/XcKx5bPLU8qrw3gJP2NPgVhQmn7Jl6TjlBDrFwO4xZ
GwqIsf9S1lgpgd5ODvR4guct/VQ8pTO58V0vpPzq4K0cl6QyAh0zWGRs2JnntzQlrmCpJzUZIyHy
uzdJbliY4Rm610gh0ZUOcjbjaTYB8wMfLHHRnKgfF3ynS3CCi3iZ66C8mxBWNrJ6dhiTA7KBs5gc
4TuyN5XW+sylgwek3Q8AI2gzGHZJlp4oouBOSOHL2DfIV8RvldzpPps5EkQ42cQ/alXSefcy2p52
LwUXbT7DANAua8N39shM03BG27Ot4QnwyNGjn5Pn87227UoFh1ZpXUyuldiQCgXp2nAl+0I9g96g
j4t5s0xKqI7x73eyksfuk5/Tu+sDYWvl+I0haGGU1KBI90ZCwTuAtOIrFzuB3dat+q7nLvSYom62
Ck9XjCOxn5tJ3jMxvIVhdZvLMwNGmnhfBVOEf4ftRnCVhLDopfTeANit7jVFw/ayKl40RQ3Ch2gQ
UD6qfFTJ8F7Q2EuMmWZBWxfopclJHX1D8u4an8H07FDQkQoFPzRb9pVCaq3VZtn0HRWRs9K91LTf
SS1W92nT3T4smx+aUuhCwFnKlgHmV8nOLteZdNdrTC7hMuCrH9p5/U9WuhPJGENdpK5GC4An1cAs
Gj1em6oQ7FtEvaMKVuRW6VN2fbAtBc+Xzsis8pryqHOl5nl7DBZDvpjByiwMq46qr/CvXOjV24F0
h9PiTfwNCSPVrZf83Nu3uPd8GGpPdQBr/iG/fZMi8SHmMI2oyKlxHiBjaoddrtX2q/mukopRNc1I
RETXSEfyQRdpN3vY+QyOfRp8gOqLccsbopnXpkYa24fjUFZOAogqSICGVN9rt9vbyk1J0ulpGrhZ
Q24r3qKonXYDIe68DFN3gqyiuk+HbsIkiMs7gNbPfikz5/xAN8onf3tjDEMrR66WQ7e+9oUNrfgH
TbdNE82q/foGZFmBymnFmWHtZMpInhBfp4ci0C2xc71NyBQMBBSErLjECrjHstGksD0me82IMhCH
VNuy06P/6cyp6ebwiP9/cF7zi49J5+zvbwdyWnYVqapLVPwh0E6RJI441mf0e93K4sZbXfpnRvYI
+vqW2tefWUWu2oBTZVUPS/9fGhBukjE+ahRe5cHouJtqLWA3PmW07pVwLD6FRf8tXvVzvesDmye0
Oy/+S7WXw91PAGh+OVoSajwvAVePkiaRP5OB8mEBOxV3VqFI24H2+ARfeCBrJ63eVQRkyKyDJ+LQ
tWeTeWj342pxcUlfgwKvV5WmKkXkmZ3Wxqdq9h1eUUDuXAImEDhdzYPKqSem0+D56EqRyvwSG9Ps
Iez4JzYtyTofdaQio3qAxkbue/B9FUrYnw/F393YvlVun7mU2bKb4NAyQ2DfD/A1I+haPx9gt3QG
XPbbEsHpvBcPPd+GWAHNHG/2cWoSUZD9CchvagTB58My5D/6N1hCU7vIDewbbULG7kucG7xFsRA6
JSMC3AvQi7vScO0Wwc8VHEFtPIZPUk8Vv1n6XWAVsmdtq1vVSoF3l7oqEXD5PwKVDjQ/1AlHJMbJ
UO1+van934ZVMNX8FxX3Gg/YHOvKG2S48K/QXr/s20PkIVOMwZt80Gf0KrUxvTtkfLNqiVlWNtR5
IwJVuoTM2/K54FeOf+GXMjWgzv8RY5aLkt5ApMOOJky6ebBGndop2X9EJfkkrQmELkkC3wZ7ntjQ
qfHNscvtGj5ReRRQRHzXbJkighup7sf8S5SAJGVAgSxathdzTogoIGhqYDx1LH7J6acefsDMl/cK
BrDmRMZxVCNTmIGbGXEuLXi8/K5VaS7HM+M4ghfBP9rQGJEIGnNBdrUS6F2wdf9Ytq2ZnSBrEHFE
aBQOIEE0QdFK6kkKVlpXZUCQxdYdvfoa49jcEn5/peH4OxvtOaoxy5Twt6O9OtlfiIBCiCVghv8g
kfYh/Vt3tjMawnr2OmDWEeS53X/Olb/lQjVqASOjmi2zlIrAPuzSxHf5jmv5NEbv0dClrOO7CLcZ
3LANBq+LhaYeEtLa8MdfgY3u7bf38riKaO+Xk/IP/eVco71Mrc0fLC8qmMvnmNE8bDWwnMaTUwJh
5GNWla6jAnZv/r3WIA9/SFAw9+Qxrr1a+3lAxmh1OSpqwRqy8a5VZXha3GVi1hcLzuL5PmvSL4/H
ltKy3Omb/3HiAc2Zv9Hx7s5RQL1KYkbz3/KEQdq6UblGoTOrFF6Y5JCZqF8OF9vde+Gdw8/byYhf
d8pzxov0sLmusmsRY7rWLis6LpboNAf2MB6n2Ch4Yf2Z9W/fDYIvEmqVVOn55x/3zKECBreu9cnt
EDAdaxZ1C57w+47p+eyGFVqjBS2cmNdScEdFo5epUagOCKbwBf5QcZRWsqk2nM9pa1vW+YUF8QBB
lL55sjAyMfQbbNbUllWeHxwGtzvGY0ttG4Wk8D328DKbLcWr+HxG5TB3ghQFVfazkyHgdSqZ0x2W
qdSRL3r9OgYLewOn3IQsKk964D8Ex3KwflMBheKuq6OB4sUkyKolWevNJdas5gvFMWo2ESXfcYKY
ZRkSyqCXQYQOhok97IWbTKP9sxb5yewLjR/q2Fk1kAPDKTmTixaE0N5Qn9PFbC7IOL6BqRz3Uex3
Y7prRC1ITGWD3MfJeKAevYsNWJUr7H7ozmlUXFzw2ucZVJa4F4L49A9mvi+h01M+6QG1CqzyU2C2
GecGF+3M8EcRk/CPbMZ/94ivuWsr++httxdKdcxDCLZ1Evw9yO0UHcV/NmxkvGVNGEpZzhVSMKE1
seMc6dKU1L/WSoMqTJjQFlKjAUJTKsEh2sbvYl/SuhU3pum4G9dzEH9Z9cdp4xteuvvq9k/0g4H4
cCpvoF9mh0YKPVZLU5R4Gl+iV897wPVoezQ/qyJTDldpZsCZP64bZjcqDbeH6oy4LGtVgjV/VcQC
XRLJQvg4txoC1Wd2N4GQbVSY7fVYzgIql+W7JbLOXrsK+sfmcTepij5TTiuqH7FcpiQ65xtSHFed
UbzLN7LNFSh4idT5e7WrKOj6RExKuq49cGkH1tPMlnb5a8402bpeeafLc7Q8Z1bciIyi3nN0SR2q
ODeKXcdYslgnOWmCouszu2M5T17Lvv+QeMY29sZgwFSvofs0BVJebew16OP5KO9YbnUSjljvK1cB
SfWsE8EoWVhPhh2EgFa0jVYkz32Ab3eKEdIUrLoYOX8UjgfjHazj/QrvAFTJz0A8W950dqnBWWf7
K0tZcU23SNK1SqT87l2LQoqKYhbnMMQEJeijrd+lLsvyxwTwHo3r4N+R+BmxPjeXoGqpWmi5V9OJ
hCxBqwc3EQGbhrGAOz/ddg/0SesSsu/gkIFlU60smE6IOeFrlghmID+XfZaQG9SJEFx6veYTxQ2H
O2NdDmoHdubfs5BHNVUaS3pXDaDqcuOH57PlzoeTomDZcriDelDXPdN+GgDx4RNF3I63uCkUrsXp
qqzQIDKeAiRC1O1M5ENV2CmLm5FKWOO7xbmSgrjVWIeOzA1qouGyT/XH9iAF97Wob+DjNLXSuB7w
5IBppSUFnmZWYXx6d5FWLDSIWIOELsKr9tIPC1PzsTrTtxwiTQ8aqCR/fJjpDf4Od2slh/pUFg9i
alsDoRmtJhaPTF7XXke7dIcd94XYcAoY9cpIvEsrih0kY1lyyTeO2noAYpt7IuJg1G0oi+drBpO/
CDs3XKt/ZOG1iFY4P93zdDKyJmooQnairBQGVd7vT5pYSLbgmgSPzQSezDUoTKzNWNf+wr8PZI4N
Ji/WI6UfUJ5MZktTjbUGN4ETaUGuW7sV/GrG/i4BpsHeSy5MpsDS3FKgRkRktOgX3DFPYqqnZYd/
X/n+DF6R3yVrtDSjPAmoG3TY/YPqSRhIkYpo1Sg4anKEu09NZMqh9rVTJQKnxFW4hZANBKnNofMy
9xH6TL8bARP0ypZeZfFswi7rxyRQIpKisXJlLI/P1r5qedzvuSNGvhtmicAiZnZpr2rsiMnofjsp
TvtfI9joWEv9IwYZJTUkuicEUvonWZHJb6WuzmcEaRPNH5rrFP1ED/av3HGjFAy0dTOH+5hJVrsd
wwD/nSYRcQx/J+97xwSTRkL80Kmst9tyVM8P0zqhNeHjBvEal4eEJTD6pWMcPLfhJd4aSuKm+of1
q+jyYRqDkTC38rWqKWZ+ORGYF0hTBIGEAKmxA6byIO7z28e1VOVVa+YWTw53lVOZyp5XxZb5Q6UB
TY5IjT68je/pfFvCCZ3v4AAlohczSX5sttLhvrHrrOWOigWJSEa0JXS5FuyveoJ+BPtF+PzKcAuB
BU/o31esPQcNDT7SuAqMvGFvnlYaugynTWLaUPZe7mZkQ9pRlUS3HQ1Wdzkj9pv30BgQScNsSP9C
mnfD7xkRW0/XIbTeVOef6GpfxIkVf4GlrB+1jhSEIBYWFrBSXSeIg5rhMa248mkrAvNhYdlrceM+
rSnI08rmU2v0OkOsqNXENgbXXFA+cMo6GFnvUm5eX1gY7BbN+P30K91YGK5rVYYOxyAmmA5SMkaW
+40iiz9H9+vbA3/0gioyzh0zLiy2PhnrLmUQ6d0OPqYQi+4jEHdhSa6TlUO9t68IscxDWvETyhCF
mGBcxPliUUv4itnra2kLLA++I2FAO3BuIJlGa0vp0oiRaro8DptPdDB6Z2wWSJlJiRzqhx3QCUzq
++36MBV+u0ABn0henTjYgSuvVsi3b9W0uo3DNNAm8GY4uie0SgMMqcKRjfU4M4xrD8oh9hDMh+oe
PqT/CSPUolnuYsqfwgHFOwOgcBx/8Mn8Gk7nhN49GV54bdnSYPyowwN5Y7+AHTWqZuaMSWauMds8
HKPsCBUkcSBGlbBtntqtjpqtXKFWslYnDrf4B8p3o9WDByPAbLCWjU/r2zLBd26nCxH/H1rWDxsO
FGzypKODha+SoJ0T7+qtLEFfqSUw1OMRFSrpwdQ1gsb7IRmHEenfCDTEFOShKIwfImgqrxPb8OBs
4cWUuWf2K9wtEQRcZJ8zWeYFRIjH2G6mc3ATKRa2XtMH1x5Ij3zLcFVmGWi5ENdiOtLETESvaeSe
OYZmVrKhXWIIF8bOP/6IrYIArN9A5t+J6IL7UQU4Y6xTKdifVxwvZj6WnwTupFJLrB07cNuxexA4
Arxl1jGFmR4cb6YCPvspW29AO/t2bVcLbsa7Djn1Fqx9JAHppJuhQBbyRNPzc92QRhgzbmbCC+j7
SzH32GFeGPgJMKh5sHnsNQoVTERcn8yKDlRnLvdoBvpRX2iqPFYCJQBLKLspocgm/tCVAhoZ4I8M
OCtVgK2ss3UDdTtIzR9jBKpV6uMwk8o4p9e1aiFvs1RMhSFpEwN3tQbPRfi7QDWYO7jYA7i9rf2Z
Ei6fN8eGG2W6z++X8k2wnRp3AiBahi9sUmeUuUeIn0j3pPvG+3B+1srGUrXOhU7lb4Leyup9HO+p
ZDrO43ZiE0B7v6YN/LUcbNmkQ9f6VC4O6S0AdQY5DVazjGcW6ikaULWetI/kdaYAmVosgkvw1mD0
7H20FfeRkOGSWDO1D8PbcCHqVidzC1jFvNSyq4THmlwhYN8BHOF07miS6Wy4U+OLFfovLuDx7M/w
t9FV25MpJYVxKtTxcrTWFxLMVFk4wGDUwIuoEPvmJqKZzlv3IbRFptc+Ry/0iltV0coKViom0nnY
M+z7VsNrv9ynf3Njwt6h4yvK5oAI6EXyI8RAnEsC+/voq/akAXUv7iQNhPa/2DNoz/0Zm2ue0BWM
dpRilM8PfodEDXKipFDQRSjOv+Jklzz7/InGT/kcOkyHEQa+Y/n8KKWZUPPkL3ibtixy25sa+gZg
hsSc5oIzOWB8RKCRVJVK3IYqNLP5vbxQ5s4RE08YVxyisAPeXi43aVnPnjO0H1f5xEWQ65vlgfiv
VS1rQeo90LzvPX8yF4tvE0voQvFchOnPoaORopJl3APBNUnXycuRa/Zg4wi5McVY9NYxyhazFx2/
9NMkZUdJe46Ufq+ie+1pJZLUKFcTig7J87JxDVOu4Bd3z17n4A8Du27Di/WDaqUhkBSsTXqyocBy
2GjnhLzv9EolX/b+6S5x1Sbp+sKgXRkkjdsJsOU88jHuIFyApEKohboTDNk8ZN0wHCp3CDrozkCr
ZN0zJoVe1u/rZmLBnaGRrR9qVvzD+q+SCUy0vxRe3GgRohXZS5dPr4oq1lBg+9O7mqubu0QttvTM
80Jb2wGYIWT6O+QT70x5naYFJypmUSgWNl9qp62OLx8pEjN421I2VHefcUuwaAmMA4nPeL2NQ7fo
xKcIMCc59cs2OSt3oIw2fAEiJfaET/Rye/TuyNL8cehwTgwCpn8aIA/KQsJ/5pP0SKeo7pU1PoTF
Ycv1CinORYkr65T1ZkSyvl+mcl24Gxc7Y22iyEqIS8uLfdKo/Ace22JMN7pf/7gRAeGHCAqxHd5i
FoTGCZLr8Gp0B9wIVosiYSZHnYPsauneQCMFvpiQH/sCnD8NzBuuWAZlV6JnXNivTFVpGFJsBlfZ
TdGDpyF/2/WlNKES3KJoZkO7xmgtWvWLWxVellAFrDdpL9zNd4Qxpb2UUkUDZHcH6JJtoJtPxGlC
W6GRLoFIAU6COsvheNxinOWVfWatsKNx4BLpWlnSuH0Wh4M2juuy0BJCXF2t7UukVpq3DzEQ7hAk
FNsF4Bl5DOvUYo2qkERo6oG3Ah1joMoSNcgwRkQuEa+IVCr6pn7gQ1HkeFiUr7cIFcNd/2P2zQ9Y
MVg/j8ke8JV5zS/cBIVfE5K2tFY1sq4+WCHPjSWe+DgN4wwCDN8jPObJRbIyXKWcjjAdmIMdf45Q
6BPbLY2hcVEEUdxLDs1fBuQb/tUievo3sGZu/neq3rcM/v5S37Vup6St120aP116FCx4PXre8oHD
Z8RnyLJhSpC8uM1I99NNDwmW14PfCiMp5dn68Z2fghvY0YN5QwUvOS+rDFPPxIOgoyaheMD6SsW6
7OXBSU4Qs+yoIpOs0icGVIJDz5gF4JqSkOkJHJmyAOguzedLWe0S2aJPhTxHL76CnhwLKiLrU3Fa
zA2ReG0aTLwL5zZ0VDN0sPE1tvJkY/V+1ReqZWaXVQy/DyAXMojjiBWNbu42NYDlisvbz40sU+kU
XfxRZdsy/hhM9EwUpOq9E4NseuOUqcOMWsNfhbY9i7imBwI+af9eWvITcoL0bt6ljfhTZPb/nOco
6AoAa6ZAaoVdOaw6Kf2ORDXAmE7UP6Db9RnfdNeebQ7MlC8YuODMHB3pfKOpQG5uL88BvzLfvf+Y
snkkQWKbJbHNU9znl53QvJi+okRPODksJ8QRxgVz/KuiPSy/UyFvQJitH5QxEKDphOb1g25C/558
toz+x+dZADoqtmFaxjnK5OGpwTikr/iqdaGGM6l0L8qxapm6jy+EXEXHwzFN8CqJrSWnLqrUnkZl
+4Bcm9cPqJlfwHvv8Zjz6/DuSvV2vaunCwDzE/j3TwqF0i2ejif6VE6SrZVv9dZUFAUm4N6QlqfD
M+YqTaM9qKpKbAvkAU+lmkmv5J/0uwdQnEqzpL2X8q77/CjvUU5DZflMwo5jj92XX0usiXuH1hb5
2zOJk5MTlaG7enqm51tyoo9CNCusRaxP6oHosSGMrHhlT0sotv4RcEg1itUqaYDiJQTwCvOCXf+s
cpboAe5yPnXs1l+PR0XMoWBzrRVwLI9m4WS5PJIzcqJmCRFJR04r3pD68vnbOkZBYb5Xla1ulxVO
fwB9PI4Y4RmmDiL96zreY5mBqYBsk0QZ21OYMWmI8YFywfSu/6svGxPTfn5HZvaIglTGDxqCoTCU
TQr4up4qEMooYCKEBcLwfuEKQrV98Av/s8CKrAQyC+X1KeO9gADJ5tmsSjGeTHFnCONaTqQlH5h7
A0/GoBgWE9G5nas6oy8WJt7+k6BtPAaiYh7AVecytczdMzi483X/7ljkPHhxLTX2H6giVqqEfHl/
+MwdvbciHs7motTu0ar1Ig0STU7FMv1UVIugii9+/Dq7ySyEsj/Q4Lx8i3WQfSfd68PK2nLDG6AP
vQq1xOOj5xg3+6rBwe2rmEFPHK/zeHauslz9VTeU/9liulhfHIHnYHrzd5ADLyv46pdwLGXtGmxj
OsCHkTIJfjUZ1fq5G7/myAfsDNIeIxJ8+iKnuVFyFqjbElMWbH1hfeqZrpCQUn/T/xotLVYsIubI
Gc019EXcs2hxNwLv3kJog7Amku7XGy27A5LVwLvj6Vl0BORIvxRzmuBiyvFTmGM6z8c2UmMbV6Rg
nJzh3W/8bvPMMxyTQgWsliWa9zCl2nL1eLONrwZY0YYBxzYZhgYhn/M9lxl9rRHcZ0QBrKnEHjIL
QmD6e5c0n4f+hJZ1qI+rym1ryvi/Lq8azi5zW7SUDo6Ie/Ol3SaPlzPMfHz/lcZOVCqtd6CTylBQ
XpZ7K6/3emjusBiXPD+kOWAdXHk5S3N3fqcBYkvNcCnCdzmUabkLanLXfix6cv7tORBiD75yOxTA
7slhpGsApRT8ozH41k0P5RNkXDgX9OxHDgBSo/KJd3hSMemNQ2qLR4X7fnXWbSSyGmuQk9ibKav2
cJ/djHhilmb3tXqykNuvadazMNUfCuGdiqMxg0XJ1gCnoZPA/YrRB2MlAmx8M116IdnMboFRcHFR
RDDkum6BKekRd+o/6rW/WT3GzDkZHTGwu11OjxHQmeXZdLVBLUu0VbqWnOO4lpkZtkFk6bLxUNu1
QLD4SbsVqGPdOKZ+TsHg8QURxJpAckiFbZN7x+jpvyZ6syzn9wUUEBV9eIdihQOcCseq8BZYUlhU
HnGBAEZ1SfpSzyLquKb+M4I35K33iDzV4IzZTipQK9sbdVN9kdbCFD8Bqz9zvo12HB6rRYCr+MDV
a9HBwRKkMTvuGi2qJNQ52xe0Q6nCMoFJAV/licVOQTpZF36R0rtUHWLEL7DrBOFDDRflioYVEKu0
TBoBU5KDqUUGQrczKVPJzERNtNIwRRdX18Ogw3Ur90gjHMkJ4+Yr45GZt6vhKH0hHLHGbkfBla6D
XNsRfrnhZXgfhcOhYzUsNNt17szLrb3VvoWNdbs6T/VnCn3YaTPGgUMi0VuegXKS0Gfr43zNDZg+
u4CWsVjjGqOtZi247Gxr1tZA3OmFRm+1ZfO4BTkJgxiMKRdBDFDrH2/e5N7FVFb2LJ6IVllPZinx
zuAtUWipX7XxIfwTe0CLjJFkjgw0hAc9hPdg2ke/ytqZjDoWdjSLD0N5U/o/b6A36YAgxE2D7U6O
oGyYjhhW3yJzREy+X3C7df1y+Y8bx4kYe2iiKELddRiyo3QscNtJ78Fm5uuPJcKPthrnAB27Oi2r
rj3+SWQSkM/3RgZmT+3FqRH2IU72g7q7pK0zbsB8LafW/tjOG22SBGh8i34lOTTDgc8IL4/GPNfg
0QY1J8QuWwslIHY6Jv0OJtKm7dcUx/Kk8bsVs1wSgvXXz3V+ftXkMzDxX32krNzJ2LKoAGteEp6n
B0AYw0aIPmLvKDKZBcM9yO1cnfhLCWcSEz+OGA6Y9bWEovBWSoCxkaaON4RDzRDOxQab+4uNJSiv
kvnXrRjxoyspgY7vKAoaLqPOkmKUa/kK/4h7KtZfzPUeGZoTnq+17gHVBZeC//rVsb8GegFEsnS5
qercPzPUF1kg7NUKnhm2+ePpsEW3Ar7yFIGWwuSpPio0BMwlcyiYh4qg7CFAGuQ31V1rFSJ2nVQj
Hfgm/TWMUFd1i4vSyu7FK02Wqa2/X3V0vXTbZPwl1W0JeSh/F4Fqr9TZUgWJAPHocq5gNmFYug8b
qsW2ZXxrLH+QVIXrEy2WssM1MAOSzGMdi05M6O8c5Q/YXal9onB5zLXzlda3pWdy2E+3mdXreLiI
vduudCTM4DZwOV9qGnWu//9V9YIpPBr2USq8vKCrPW25nsKjlsrKCtoWf47jKGsA22c+Lgr7lYsr
TtUb1oxdLODSst5kvQRr9r7KzoLaf3FTXoiakEucvLcvH/w6hubOHoPp2LgKLbMFtglcq+zgXIk+
dQ7fiS2ODxhse4i/EHQo9voynLcUDIN8KtD2TiF3ZWi0NBCBPNXOeQVFEHeNX5/sArB0syJAK1zx
FYfppLHwfakDamq21rUcHyn4amPTnAoycMVyRbND/w++BiZ2uInC76lPQL/vZrdWg4wu0214Tj+Z
ISonBJZnK+1MBem4iBCOB7+uNpuAn5am0eU2A5S9cVwMpKWin5O9C36WpA1bA3oQ6upNDqBwkEYP
PbEKS9ry158i2PLKTAkjJBg0tGUO1xg0EG9Ns6645+2a6Koq6snw56fn/Ymu+Wia8Rj4v0UTkf2f
ExzRjuHc/wY0ntG/Iae1zCuEpckuH/iNF0AmiQxJelh2XmwUfzm/+dl5lh8TH/cOI9QIBPnvSqIT
Y2PFxPQIroA9uGP7ejtwkiLFbViq+ZtDDbvxzVBYD6d3R8Jzp94dXOhM7cG2Icx5fF5juzGifxTQ
VAN1JZKX929QgIRFGDLIdZCyeKizV/u1hRW9qz2ijcCEuX9lY5/bhaos66zIGZCCrjpSzEt0CUpN
1dEdILszK9g129mjHrGnEtVI6Ijh8WHCPtdew8SVQYHi1130PwJLRMLljJL09MCJQ2Eeiat1dsEL
vPUC081LYk/UaPgV0RQzvwV+SgkKXWgiu624K3li/ljOBPxUI3r7khjMI4xEkgrc5xAlXMiMFqbr
4CTdgy5hwHt6vj7GKLSucG+J/Qn+9A2DGZ8a96e8pRCbKcXI/b7hEzbk9iFQKSsXBqF1nH/2uJuL
b1wsYKD8pzSm+zXKXjcP6nQeCyYy7Jz8VLypzDNPjrJwvMpTPwZgEz7vK49/rd3qfNDQ1h/u0IRY
sfz9tQZ4yMNs0zEBKCYDohCQQO7nBVnY+DldGns1XQ40DObNtSrtk9URhaJTW6TdqYgJdAyavfrZ
wxIES8oveJA/+ZylmEMftXJ6xKsFr1iStEjrJH+JtG/n5m6bDfGaZM6xS2HRtp1uZ7kn/dmZLZV3
OVmrQ5+nG9UBkfGikB1J+mbX5meKx+Fo6wCTYeYrzo460scYSglGozxXP/1om+77Qq1wT7CScHZz
ZMxsl27Q3ksZsG+03JUM9cph3cOxHCIp1/5JgH1HOrZbscfkmmVv7DSzm0shSagZ3LUdfK1j+q/s
5STKxw8lV9yMiGZReYE1ARr082H5bGQKGXmOulMum5bJFTzFgqRfixno3qmSxU07pKZGonrqFbR+
LwoLsjHG05r0U64vWasWjvAZRAt8o4EqCmnDCGPzAsEqByysqacoea8fyYAHx6v7uWK0/P3WuHPG
ROtNW7S4V5nv6ODTk3U+4Laq4Z6ERlsLfOWcRDiYh4HYNEirnM0OIL5St3FApuEBnk7eJq/Bks1Q
4UHev48XCBuchkhHPuSB4XsiIvTbuovOORmedymoE6Rd6E+aA8lRoDqEukVPSkVHjQweVlsZk5QN
qJDr40NL5uD8hOSmCMSILf9fXPhR26H1eMoQ5VqfSm9xFlzCwPn0dJDNZ2A1/Sv42mmsoUmfCfgM
UpdaiYMpu0Y53/1Z7SenHZpidMF20GCxDicZTD4VDViDUywhZ0osU+gQ9QaXkOSHxbjy7PvD6Pml
JUpIwv5tzrPG3I3/zijotHl6wYJCuzshUj9ZvKWfHRBPutlkp6xK5HtPM5oh71GswygZGA2VSJs4
Ab2qyTBe7DKo9DbsCrpZyz4mMLryhOu0PnRCxozuN4tAambdZCE0CtPHWtvH8P9cvpVi68dl6YcI
vAiQy88hffld9pbpFSfSfYlX+9t0OFlZblULPuHYoyV/GZXuHgaUJlZ+Fs8LYn5Z5tYVtX6GSMlI
sYD8RQsr6rvukHcMXMsBl1LKfLgndk/V3zxvnWrfHC+bIuBCdgryrdYaLkdzaBz2UyDW3LQYU9Y+
g8PBxHWn/ZPV+6zYC465zr9tYpk4buJkForMFGXJUfzQ570Li7n7uUp5F2ZlooxcxEetHtKgFBPG
0vjH7y6s5aUzmaBA6/ksWdnhpGk1zcLimCMDoYRB2nttWdjoSoNMadrMmbnPpTk71KYSdFeKLVUD
QtVobZC9XBg2PNXAFCHGS/OwLZgiivHYNLt2IYAy7JbNLZQ0MTFdfh74BHTvDBHhc4EwcVM5eojP
dYehmFnAOvMpkhGvrKYPlVljV3mHyrxZ8XlzMcWDoZyVjXx1P68LHw4wy3WZ0bzfxaRgAKECGwHR
pGIKD6gbRdty8tkGg7MoR0/odYX0HmdQ9LktBVoIzdS95CptU2M/JqWWqLPWbqieaIPLaQdrmp+f
ySLXW17rgmMekISVljURNBpToY0MaDzLy7BkI3ZeOw1kXk3QqZSofvJLrAcEZWO7k/kbxTgCosCB
2xJlmfJOoSWvenMkmGSjJndC6gKqbc6WLaRD2J9ZkFvryD0NH7mougbYQPeD44w/N1gvS+xs4ZwT
/ewE+0C2xaaJxGcwc1K5GeW8a+9xFrrTEJu191cEiuQrNkEe1cFEVMC1WjwkYRHV/MyLF9kd2SeG
wlupXKfE88/zi+PTFZu/Mrki7HEg83q9ivxwIkO/L+rqw/T/8hk08VbaEe3ApcRJSrDHKkJo0gDy
DBuLldCCwM3J1fdHkVnr/NJvkoIkAw0Vjt/YcIT7XeDY2SmUq/kq4SrDmS8kuNz6QlaqRyoBePJc
cSXfQon+eQ6P7E1+FA+/RwOpmirG3QTNKf0NkjbzD/Vn6tqRQhTavOIWrphGfRVb5OZsRCsxgK17
EeS6hkj9+lGkGObqRda+vNaS7HCZryVshVV3i53IIR+ctVAdurAWKnZbmfuZ/yFYeQVhy1RSmVbv
9Ql4EjlHerxJOupSwSCvfbvMc6tuZ++XxGnnnLMRGPXeWCi4nlYCJivRbpSeElMytqIQYNWZEGLI
dAGJrzFLGNKW4F+6guDecJKKTigzfMhdxwGesNIniIBgPGmrUVz9jeozeNwlHP/1wO7SsXZVzsUU
Cj4e/Nv0jOcrUW8pVNdOHn2yIcvL9XPEjdkaUYPqbc7/lWxAdbVr1CfXYi6Lmw1GTqKWNC0I8Ut7
oA+rKXtffv9e5a3jmJM2wYIMHQk8lhJewo30R2MdNHQ/0WU3W3BXNcGcS+ufpGjuy1svT8IY61A/
FjRK74sP1VrSTVo775EV7m5rziNCsu3uOoOTKiwMZ+2xCoItwCIrm9936zUipWcGIAPcunlmfZK6
nTS2+NYmxam2A11dy6NSGWkKKEJ8PiGiTL/ep2QJp508S9MnFpff2a2dOuHsl8K6S6KUFxbtGnem
zlEtdGB8KDXsZjtFOQ6k6dJR1p0QQlTQbiSlyKFaukmywJDgTroulb3cs8tXsVMBCWRumAG3uzr3
xltNkx39WsJhRz7AdTjecpK0eMxBCGNSjO7vLFo5XeJQZj7G0NO9VNbwckwRngWwamaXvM9QgBxX
mPfl1w1tb+kGgYA93aAbcyh6t3+jX3h/zcim2CRoLKWtiI8W25HqpDxuySPAn/7tR9YK9vfchoXx
5vtbNIAOsV2VFlNgpFHzcCfdazXVmmVDOGPQ50GoPx3/o9qNxp89w46Q8v6NRezH50tOh+RVQgZq
rnGSNuFYBbgnObKzzF6GTw9QDOVuFVTE7TgOaHQ294eXpVNx5Z8k4b9cPSrn0DNzYWQHov+xUaaJ
LHBayQkgg8+rF2T2vIIViYwoj1QB/9S/0YqePpOeNO41BUtsTWJY6wuMUVTm2jIf1ZvwETHaNRV+
sFe4lQvxc7CYPpKDUXH3ZrrYA4NORm+Q61/NIMOutJe3EeJxy4PfjLjkGE7CB1WIuzQ/Pi68nNNM
UXXkZraNNCGWj7YqdBz76v0rhMxbpejUxqpSv2kyMTg7iy9yL3e86cTgNEHZKvlIo+CSum0Isxcb
d/upA91xf9t3PKBwtZMBLz05rsQc2mikh/lmTaI0ecDuOX38afJTQ/T4QpoBiN5mdxzuk6HNvOUI
F7LP4DRcEU6xxKwU/SZ8D47bGQtDvkx8xW87JPUhydnrPbXFFi2d0JUsqcbr9T+Ts56LM7ojrfMb
XVylFhQCx5EvlcXDP9uydt7aziL5I5R5qcUSrRxqtsMD/KdXqtRwJ8ubrUvs6J6g2QRgFgLOLsfd
r+F96IuGgpMKBk9lOl7RJAKR+UUKHDaNYAz+RuAeIF7IvRdhshrWOCffFjqNQAQ25dosYe0g0NDF
wpTkEI2q012/mgYO6px4ps2nZ5nfuO7syjL3HyTu3MNYzrpYVNF30V40lDE3NnDUrxHjuwvKrnno
4h474y2MX3uXvqi4R3JxRHSAaPLZWea1z543QVllJIP9o58RBzsmq8N0X+lzvNs/1TfXuHJCJ7tR
ikIZRbyZJJBJ93enopiIA+4Zzsxo7HVAlyON1TICRXJK7MGzhtRYTNBI/KpzAba1mo17CpQ666GS
uGm/OP4LwxL4XYIJu72tZ39Uw86GYP3aGFMmYZVGutm2d4gvoIymyFz8Zg8IExn7auuAJjVtTY4f
QsbJvntDlrwFyH4uK3ZCJlP0jnneCMXT+FwVfqngFTE0or1ALF86bay7daIxOOE53FsQryAFRjZK
XxSbZrDQVjO7l6OEXOPabPrNM7nwukpTFpbUSdQ+4mHfsTd5c69EAOrk6jiLFzbWgu5zwSIh0rym
Yh3uuWZ16QGNEPEdxviQhGeTJQIbEnVUkrNBCtymx1rHQgnEF+ytLenOD/p7FyY3SEjga2K2OwTz
fQtHupGchc7he+rgfYbKU7ONrSYO8ouMP1C61Ifwmn11YRJFgzjD2oJ++7h3atHZLPczSFK15txS
C0Ds+9wFDEPzKK/jwK7gD/0Kv29XjdJ/G4EU9MtTlsaeX4SX6y/IIMFE61bNBroMVtoFaQ+NRvjg
0wXG04V038M4SW47HI0jQGEtg7a74MwK80iV38dcAso4YGlBpVoZ9bWSZcv+RbJxW2QV4vt3GFXl
QaEPFnq0IZ4FEVxa12fmolwvhYlmlsqODV47LfQ27t3MwYjT5DWNtBOR3ne0SMAHALMMaaIntoQU
IhXtEMZzA2Sp9BQs2BJJnzSRGHn/AJ1MAWhH1Z5YkCM2+VuaFUU4YoMlrcabxQ3Xn71Sh0+f8DJH
tQYG4ui6gRfM4oAPmwbH9xdXH1BJ4C5JQjOyxE6P+vCc/DahUCbVy5oLWvhVuN/9zO20y6aAH8X3
V9Q6uL2UH7Pm3ZibCCG9jHYj4MTg5OPPUhAe/2ivJLCpRr7fqJMqrcYkj+KgiGVdDxC0cmi+aP7N
8KkAAUSDSoTaKuIkSy7a5tMmfTiyvTiBdKhrtYm6CIt1Xe1/dU9aWmZtz5t2vmi+R9hoBd0P1Hdg
bqJhTSnUIIVueUZdvF/a6Nyai78SlXcKkjiURtqVIjW2IAqTEbpxI2b/vm63i/JNgbOrnDU8/6P4
KnC5BrpPDnx7Iigzr4lW6NcwRYDlwGK82iCqkQHdacwtMmTToWAWOPvb4apN07QY/PAtyKkrTcuo
rVzcTbLUhvoMnj0e5zNctSyrWPLWEY+K4UkOqKJTzbi7Z+NBSiAGhSdzEa9z6tzqh8QS78s2VXTV
jJB9Cz1pb85m4A5zh0XLFQvXzQxhvbjs8C9rpa54q5MBrEts8PaofovFc95FELxK2oJhJjAiV0uk
XPX207zEo0pWqY+SCqiRpjTs7q1XqCrS6ICnf3H3MOQsIxCBjx6j/vpnZ4GxtrNek48ku0LhrswM
qgNvNg2pJHWLYSa3kLIpF4HHKLYcaOsylRnG7XipOJHdghKSU05kOSwtCsGiEP/qulwqllOTHd1k
EToxlZIxFBfgFAuKrZLgljxG4+unNPmu6W9LCLCA5y9hJ+aikCu79F/s3otfEx9xRYDNx9uJo5yG
ODPGYCAQE/JQ6zmlJPrPB3oVWKwjQRla9NBO7VwjbbmEIqkk4G9ahlhXp531GNzPo864uT8QFhGG
G+FY+a3QTNKHQqDCWGgndVnWWHbzWthJa8gBE+IKo8TptzoSdvHVvDOYcKcyDcjDValk7riW97+V
IAlXrDpg8mKAx1Mxz8c6r2nQ9R2+WxWYT8NLvaWAl0ApsfW6AqDVzLtzshp51o9ysB6Ik7Zu1KJp
WsF2oZ8CN/iLniWqnhlFh8kcKeEnRM1fLGVkjvWdIFxyV4u0Ut0nWGazOsS7BkuRbogIqN8Q9IzH
Tg1Yp7q5R67CzptPYV1fClH344G9YLwrQ53tsSt1bLsrs4q16wqq+5RXhdsh3w5D4hMj3Zm678GN
cvz3gaK+rcHfHWHtx/B9UD3urxN+s9H1J0yrabtfVNk/CwrZOrVuAPMY3OnwPcbpMq/itYwgAUAv
cLiFNfFaS+craYK1OxXr90EF18IL3VLWu1VvUbP3VZ61zrJdyT71nbuVF2Q3/PEmJQK3qs7/hfFB
zMhlTwTu/aVRBjjiZdPDAG/5PI+1pEHKONnELZcQwyNJMKyFIXb3Oi34/q8IwHJAVSCNeYvv+8bq
Xj37U1M0Q91+oU1yheNi8QfhyUr+HSDAS+YxgVprrRzwd6ON3h5Rw65nNAcsFWfLm7TFtOAmPVtk
7Opcwl/g2pNbQ3xO/X0KLApnaael1qpV+NX5m3/pXXPNhkNfeVfDW10NR1bNRJ9ITjxLefanw/Q5
+29GLkJtPK8ZrLarn4x3w+4480Ag7koROxLUHAfPEihgM/cjGogrC4zicgCfzJjlZa7N7Vp4pCPG
CzXlZDbMxbtVTR4/Y6eA9f0y5Xyj75kbyUNxC6yCJa+BrDt5xHlqWvodg3oukykM7FPP36u3iXHj
RAIb6c1Xdq3wrcCXYy4/SFVHT1Og4sodE2tSWKsAub3d3oG8pID1jN2BKXM78tcAQKh5WWUJZTVD
MpzT2SwWkIA3ZKMtSpSJBuvBoMmA3jr6xLUaudJVjmf/hsmUazRA2leBtYUxc/ComNBI/NF7SJW5
B0PH0A18DJh0Vox/fGCwghr5ZhF0slO3HACq0YHYLu+uwWg2Lhp/aIv7MqpF/3UmqL75MIybIOXP
A7+KHtMA3Z4QLqO4I0jLnSzUtfOmysn39QDf/ww3fghu3jalU8LX2+CeMojTXjUL9Xe4Gygkgj/u
1Ybj/1w6gUcmvC1VDaxbiFVsP1cyShRg6VxP4pi2Pfzpg42lK5D/nDotfN/6mmXwN8tY4MhHcOWV
CimZfp6OwGV/NOc7qsdVK57wZVfwJdVMvwfDtECS3QfDZq1+l3i7KMiCfPqGsYMr0EVtnQPoJKuY
TvG97lGChGKXImiKuEy/yawM+y3CImCZP0Nvp+uEQt6Wzzx4lD82+3vZJcMj/fVJ3TB+oeQLlo4K
u2cEldPAPtmVBrjWm6jYxgBM/g6kkg0looEiph83W5+Yp9q2NxvFH59akbG/FsBUaW72oPx1ZuSr
lIpmiC3r+nJdlk6cX4+R6f2btnUiMFaok6C5zJFETOKfLPfyYrF2kNTWbrPyO/sz5o9Yk3UhcXqv
cRte0b0VPZHWxUa7qE9cu9Rxw+7FKZd7mhvvto8Z4yie8AOMpkNE0sZyIXZXTacajuVAuHNBPT8k
UGpb9jwA91j+aPqiJc52PM8xHyNgqsFFQO5J+bmxHu4UgmCsp/6kSe//p3JH0KATDhqTtw7eV368
HwRZns7icL7bf6BP583ZqIC1ga2cUxSmDvgu30P8KpOE2hrA90JleiWt1C5vZQ/uoyCVreAUyLdl
99Ph1KlLu0m0CRS6aH3LCytazGHZoycAbzh1XCVaVTn4VuaiepajlM2IbJwvdjrWddI90r7KQ9Bp
Qcyh6IcTKcRHf60nMvGWF5H+oo0THeq5DSOMXWmSUT+QaUJNg6UIharTMOc0HLDNnplFcMEDQImx
jyx5NUrmNAfTK+oerzyRAETIvhmt0UhwBctO9YwQud7kyt35MFhX74giqDW/qi2TZA4gfk7seOOU
Qa0/SsVSLtsabRZRePuurtdoZoaftIlImAyAg1kTb937ElarFt016qBPMB6Hqh5a2QhjkUE+R8bk
O2US9tL/AFlMHJP8X2bnVu6LJz06wvMFSuNCqts20BumM+aSzs6eqKm6HKJPi1R99gewxAJDVIxE
fSUnylyNQPYGVOXtY6ztR7ebovQd9kE4uzI23oLlC1XPQWIcNdkEYsjfSUZ1kvgdAPmAwuKwTp7r
xdWJVL/cLPHaTPT88A5wGbQXQ+HciMOEQ24dNhAFIEs6JApW+//rJQiLgCMB8jKuyeOiU8yUjSLX
ds2tuwt9Q9vtrKLlr3kzQPiKghjU9bcpo6w5xVH8JaswO7gg93tCOBB13KZ9Rr/1Ewq3OIfStes9
wGyBYJP5Bq+C2MtlYAY+up21BQqJhwXBF4a3yPyZAUyzORPRRbN2anFvpmH3nk7d/e1NOzEXDpPj
J5QAVrhUQz8RFwi5Ta2On/yP31jhZOcbJmwa9Tk2XB1XqhhOdJN0Do8r+fh3cjwoIdehPy1ce8z4
I4nGiInQb3PL2tHa5y8jzz9fwewnkHKIk6XZ67JfE6Qk7/lxx9o5Eyi+QzZgdHLGZtqZRea2Viiy
EvR6Js+eImw6hmkLox3TXu/RzYPHa7V/4VuNa92+EaKsR4+Q5pqDPqOP/x8Of3v8QYos02hwiMft
DdpHdsclssCM/DINTF6ADQ0MdLIvU5WXbB0Nrgd5PHjDJP0NIP+8+BAIx3dTWm/SkA/4IJ3NJKG8
ZMyKBSZa52RRG8Gm/tRqaITmZFyNVM/HrnW5BjQY8zlInbgrdqGceKQgI5QflffYqyHzkPA5MLJi
Kn8CNSGlk4+M0WPvFzc+4SmsFxsDCJqsnLUpP8nA/1PBuc2t+sFaEbH6jbBzC8ISNNXQhEFIO/Md
cS6c/N8613PR6PA5AvjJhCWZqozB+zUiHfkLQZmFU2m4h1ag1ix5YcTIaTNOiLTLqMQbcGHzvnIZ
FI4bpf0vDeRd3EgRNPN3qybrcuTZk2YDo2p3GqeOKriFk4rrBcyBNpNN2762gLiP9bKBHVJBRVoc
RGQ6tKukufggRTc8+DGzAXYmBZWb5aERprjq6BxnJija/EbyLzPNU4D/8hZCyrPWwmvsgsScqk/9
Ogohp8r6Z5aZTnCOjGUplBcq7152piD7QuRTpeoLSaXEDUp6Ldu8q7yu+4oRd+ArZ9nx/gmbwAjC
XL7X0Z2+JhdqC7dmlX48phJQrqiz1iVcMD+u0RU0zh1/uAnRThZhLv1U66mXyGrIpNuGpILtj1xw
6ZZx1O86E/2U8AZGEbqStaDVXUDsskSPGQO5idVaSJGqYlLt9+LBdz7701TaJkyW3e4sLWZAl8Wp
sBrt0c7bSXO98m/eTkYK3PZOgxXzo2DyFugvVeX3sEFauX/iRU8vKQp+NabUhiktJBsihV1hR0xP
ORK2rbBIRjfX4GU+2WNjwvU10shSU1FOwGUz2wQi7D3L8tPX0FWg518gqTJbjMqQolg9FhUtpgjt
Q83r1EQP/qv9AHhzuaSz3KWML+RdYFpDTVOk0lrP6MJhIj6gdCjPGNNb2RTdsIJIHMU7hX9Mt7fd
ZiSrNUHHNkJBHCBYyb7K3vBki4G+eWypGP3QJP5lh0RlYyxSl16mL8MFlYUdIA+VMrrDLe7IV1Gg
9M0gKbI0ZJoY1wIZj2zh3IY0LAykxoJtEQT7HxygJZw+muL2oxng1ZhWdLZkZRKX9liO6Rgg3KzP
aCRVF5xb17uajFgs+wXDR9sPSq0lRGv5FlddF6OL+LRROl7rGDB0FxjuAczM9sdT43YnUXDYsonp
/OO8EKdVTy8tCqfMMbIa6FbRa3t5q7ixobjKMOXEGmoZM0n7nACZ5zab0xUmjLPbtIhq+yokmVjG
vSAJyaQmJmq9mwoJBrO5XI6dD7As803PDBcOlzU0u0m87wcivlXiWkGPcvRxZthfh00YRXHUyLEg
QcxuRP7qY40yv10SI4kMnt8OuXJJOxlhu5tzdpfZIDMgNJvsLyz4qpQCJjhPPgQvvA2INwndJtPr
sZ9Kp/E50Rjwl3I0RU/Ku8X8KSYpW2ztVdbgmdslT6FzvGXWa9cgMgCUYWv+irwU7DsYUIU1df48
98UaYhiR/SAcO7+J2gzwbB92Bs5c5wc+Pmf00gvXrnVwnt529Gqok8ISw050WD0mN/ISrBqRL/GE
hqrTJmjgz7dG9qRnJctqq85CEhZhMoWLw82yPENA1zUqCMpPyDEpqni5yAH9j1KVQyWLJ69P01u6
JfuCQw43c9w0DTnMA/IyRoTr58iDiWhIlRJ+Jz0Ow7XpbqMOmxDrBMnhHP912BKyUet0HOphibKl
JOiNeQP8F4wVI7k2Doq0jR3Y1IzqZy3hpdtyu2xPQu72+36nH6xASqQex4JrIsWHTesNh5bIx0qL
nHVJprM5LdLrQnopx0JrgZDK8zHHqZ2WjfaKUxKNwUZ1Xpnhmaw2xzDDcpq2xD0ExCILH5JCVib8
0qIoQru5nsiudZoxZPtx/Q9W0CKpDVukrlDSmoH75lW0tRDniVWSmN94lj0kgKBJ6rc3Rhc+X5ib
lRcm7UrUlVoXRS3Nnviea1iAMFSvijGGs0FQKBoU7aBPMi1FKOTB6gGDCv32of4q3ALWvXycY2gi
Z7kdFe4btUSD4pYRZ+6disEMCCVYKFO+piiYYE3xpoPcDdFzPM9PUtIHnuVaa2/FAGG4FZ9I4Vlp
qOXQ1UMwIj/rH6guBGk1K8QwzYrob30M//EML3dq9YLev25mAHchQfBKTuUf3GyCl8mtU+v0L/4Y
z2KHCMMSrdgaAD8DkVSw43Sw2AoAc0VQTvPAqyHDLpK/Ku2ef3EO/COcgpL1SeP9UATpbE75rzvu
xtgxki08MeFjkv42jTB9eN/P/rA7V7lmPSNStI3OOTL3h7q4ZcTUZGtBnXE+uTywUlSMh69QNrAt
tNCh1AqV2l50+gvPUzjuW6O5Q9Mt4groHLw2NetVHm+ESFg4dQn2niPnr+gGVWaAmUYMvhdJ262e
/ekVuwzngTKAWfhtvUYm8TPst6NHIm5c9+eR1/t2pO/9RAgMqMlUWtHvZJxOSJQdQdNdgkSTiL21
w6cz5O/m/EHFq3EWjMgDkWHN7n55UjXDwm9SMv/fBT5F0c686+zsVo5mv13kKeqAf9oPw3glVICm
zl4KggHFmD3HBSTYhgNUzayFbPSX31+eAwTJFgXKUhevA2V4oMidqL/dJ36FKvI4CeFxOsB7IhMl
pOPDuLT/5tOwUYSPR7obqsCSLuyVI8qYewPb7FTFGtU1W4Wq6AeqEijBy7HMVw4ubi2LGMkBcN3f
OAZgi+GpxEbUvrurrjPzJ4+VEG8xFdmuycB1I/Idjahz9+fWfhHAIq3xDCIOsptIYG29U6eo6ERu
TXzwofqEu7V3doSGY6hzJu5qlrC7wXgXw4qQ2ciqtXuWo5LvqNxaquNYwZcrg0kaNHXzjJ9xICty
3Osy6BvBOiSK+wpxk8q74nJQiLWlUM9Mxnca534HlZwr+SeUrP6Y0hCW9tKxgegXSbPnGd7cg6By
yCv0L9c9JNwQotbh+dSZ2cjxSi4/dcfWcOlXZpgt8MUKQWFiEo5k175chXpvb5lfl2dtGOcvpqKa
hVttM8pAIzz76EzSiQA/2+43vmXlo2Z6nqmEo6LbBNB4H7gYJRr37+Wry9Mtrk0E3cCakdCIGwFe
279w012Q2d93LHEGtf/325D+7ylv1cInm/C6q/+7vif+9jVBHfEMHSUt36+aIaPMKI04kYareA1n
v4W709f7k7LTmHwlYv9FszS10fP+0xRIQa91XyxmLK2JKO2RDcPBURFIC9xg4DBOA3oIaAbGjmYo
GYpNQrIUFEJMconVFfgNL3VGkqbqghopb1ziCo8/bfY3KL/J2tJRocX0dN0JRMBmIdtdKftacyBP
qWA4R8M1+TP0yb714mfX01rOuVWCLtmHJVDGgrOpRI2Nv8AeDTVlnsCnaA39N17FTsw/U5Uk7SCc
SdEEiyX0KWS1thoq9IcfN9rJvlqYzv4eb8U9smfHzBtjudsGXFlK9iTu/tlZ8/STTH28a1gn7QpL
0TFUtC1G1/okuIchVmukXVXC/ZxSEbG9oWx4a7+GKPAVXBnZHk5KSZ5pHi6xsiVv3LbJeGnAvftY
NjEVOrFXFsNmlVH76z/qGGZuUY4PjmGN9u7AQUCt4iPsc+/UJkYP5jKKFcF+B5X+m1refBUAmKRn
dwDTw0Uv12Prqf78HwPEKruDpkNaJ9b1WKAEAk+q7wHF77ogvjgGlyVLZ/tANNYh+tYNdP8Oue0h
CzI9lyHWLD7xj+qNc4a9y0nv9qfl7rx2EwLO7HOMRpOeENBC3nLCwDRfafKcp4sqGKeWoghhSz2g
O2uGm+otFDkFe04gCmFuEHbwB10BVE1Doy9GTMi1DCa3P05EARNHBuDd45VQFaAirYuZrwZ1W6vF
RK/ORzI+WAm5JRhQ0I1MIsiwvGyfhywzgAdDVtW+ziJxJnSGrtrS325K8MPjad/0ztv5iqRP+Uri
OS/2Cu738iHGMKLC/XcI7Q+rwOnltoBOBGGRKKn44ln3aQza3XcZLe4Q/EcLQTTumPZpD6viMBiU
8A0DprkmKVA7MlLL7232TyKY1tFbhQVMIEObYysnJh+AXx6GAZUok5xg/2zyOcZV/1lF8ai/TXzd
z54ZRfh8z5Q76lMcGDpanqL8csPjIzXMXCc52B7CtQzzgw5nof9jenZbmVpvrVgXW+RGmGGalQah
XdHZiXXy6C730EpDq6ocE4WRmUrcxtNMECQrNFNWLHRmjynO/wGxZ5wKxg2iOaaCy7++8Fb54tBI
nkju5C+wenVw5hnnbCVAtYJn7yJLVGcoI2TyRJTO+03akPveJHt7t2OM4I82YaDG/SH6k0wGs/p6
fQ2TYHzu02oFa5pUq4EmTA4s+r9nwm7m7/BWEyTYxe6iKLMDYKhQZzB9wJRSZmuCU362eE5Z3A8E
NMVEVR/a/69TzFyoRdDjBIGp5gQxl38y2FlDTTQto+Ch8ai5QRUpHE6EhIpeYKe1QIMqZtbTjN0e
0Y6v9NUkBXtumSWB11X7lfs1Q1Lx+IqdjPN5uC5ocqFCFLFRda+0fi6RkbX9rrvPjmn0BA82Qal8
bnR7rTUqSUZGZZFXoosGnLPgN9j3p5eWfL+P9bvxuhh3jIeu4wwhprhqcSTe67RQz/LYOwnZr70u
OFTalFJtJ/0YHPertLYs9PjQzcMenMcYGZq4wrRdNTSb4nYYkyZDl2OpFgMXF2RQOyWGw++CZ8nG
xlyFLliMqS+Zhr78F7WRBvOyaXFJAdc0JVJMqYp4NSYX19Su6lzbko9aetl0jplkiPQuR+TYkRoU
l9hFwAFQ2q9Z0EORaEDrqtSs6iqyUxHpkYzmMLfZqQTk/1A65cYpHnEevu9aoqDGSJkL6+/2sOWT
BIQ+I6NIB1qNN3ZD0sYr9nCn0SQ/cd4WT5bKzfVTv6VhCE/qx782Oa5zvWd3eC7yMcxwQMgOZqQv
rOH8S8OXcNjVKv0EXsb9gJKTuS7i36Jagy3HMd5GQV1CX92GHX4rUVMvTgH3L0wYIuK+ZZQc99h9
j2a2LcHrkNn8a2GawmNcx5+MYt8C/YiacRB11w/SUefAisjrLILGh1woybwp9TQEFZ4ZZdKkjYZR
wu/ZWnkEatcKqr/L3fH+ku/IJxzjRSQZvKh8ffKez/DFYRYUI/YZzf7zBBVLz4jhPnrBZcZNKVu2
3ZRhKgZWuQCYArKN8O3xpyyvL05b36vSGh5P7IXXXI74HwuETgCDVHT0KSZcHkE4o6QZcgsvfYYT
Prv0h+xydvbHfnRTdZWyxUINj1pEIvgXhkWlHn7B314CzE96m2VBQVSklZPSEsQenkBgJ+WXUfTn
yZRyn6B30WloE+7SkIonoOAFLZzK+lbXUmHOqj3sL4UWKAkTVVuKLrFDttwuov7Ah+LIrnsrQ9Qs
RQ7L59F1zFrJXmU2e11S667G/+nkKNIdz/bpMn8UtVx5r+bJJ1I6wm4p2lKvsgetPfQ/EfzbOFLr
UX/N/009qrnen3ZYv5XAgB48YjRaGx2jcf2T2oqdCbbSB5n5JRXWOuUWy2N3JYGY5aLC+5lmB1sv
rfujqm2AGiMN1Ad0/177qtXsv8Ccw4wpdLsACzpDLRkat7yvLzGAsrxTIr8zatGy3rmOOgd0d8ai
rZFmB3sXfi8bC/tQQgRILMDH4O+Kavz6th7T2xd/ZpthvcblVVRxpnqpG8eYlD14p9HjDBl7McNq
v+W2duX+vE9F/WQRErf3tYu8RSHYHFQQazSXyngMf/OITpb0XnrY6zdBdt4bogTelqazNNqCh0aX
RwGTikuKXDV6N1f33jT4R3HYqx+3+c1EKrc4qzP8esGXrv4BYtY19ebuPzk/MRxnprlFW7fAUXVX
ucDKWtmhXs2na9irf8M/S/3FcV8ETJORxyr9bxXoqncHfgTW1+N0OBe3JhnwJW0t8KC2pfAHWytH
DKAxa7hDCVM7TG2TSRJ70fYBf14oqk7w5Df1fcigqfVs798IvA3Fs+udUBjQahs+eQ1cjAtUSp9X
tTn0l29gjCLwRaI8i65nfhbHO/k7etu8zzbH2xUjY40ev93dx+C0WIETW8S2gPXHpZ/gB4pCyZtX
FbgcD0kDJSXW6qJpAIT9TAEQeM3IIe1HBDm64CBitN/9fbi5cFJ8N26Ogend8zEzcYa6VylPRlpQ
kOMzCGcFR/3aAE5qLLCxGmoFIrvnWgN3P8mzYuUUcp8dEVLXWSC/hdFK3up031dKX842qpAbU4g0
Pwfae0/oWvTb7BLfAV9z5vGNj2qJAvxjf9gPtOeM2ohWXb6LyhejGF9bUpX4bYKhZNHij4c2ZX3+
fAwRLKWsSvYnDh7J7nciP/e6vS+kVvMioMyNQBJG5dss4PPyyH2/AGk1iVCPeUmIeFzuI+xTHDXw
HHyaIQiLDK5HLRtgzYwTLEdW5D5puyXBenYsMTPrxW7tglC6k8XY0Y0oOImzxf5PO1S6fYWRg5z8
raewaVutaunkUqnKBV8p+X3T/xQTKPBbZRuoisOZGiHpiFlUOFLYELLPCSACgqAnllnPnzu3apaW
6KpopRWgvUIq3MUxlEOsrkxvqHgyj7E+L1A1HefTKal8r8GKUfu1XxWfEu2N6H+iWBM1y561OwD9
RpJJYfFGtoNql1DmVVTzLyuMRaiu7JSVEaxYMmxsnu9hgmZZRUmn9HWmGU0IywCLsy7WsTvvLD6I
F3agbGVsSJa3/P0DF8yyiZF7wl6kbcJU4mAJhbfeyVbkOzw35CkV28FS2YGrNxYjc+WyJk3iOtCG
wAZk+QUF31X0qZ+ZioTy4x0nJwkOghoDes0ueVhPbDBMDAa5d42RF/MPMzv+EAeZX+/MU9LJFES3
7Dlz+OVQrCetwklGfjcpw+ME2WlWJVPWbG85298n52XdmWvK2fl3GLbVblHZhIdiHQXtnTTI965J
scDkBmblZvjfxoPMxawN7mhMrIbIjm7GjtJm59khTgNax6aQqG5wE1GDPkISr6x9iEOD1vbnsPWm
xoyqK506BCMY9+fxWG+D0/6a9u2uox6LZByqmWV3RFB+6xpf68l+x8KMCb+iY+1mkibMLEUFDVf/
jRsTk4hsO5T6QEmXl3U0QYebvhLjb4iP2hPWxajl10Hw3iPQxKB6T2VU7J2vEko61AQu3UFWqmlf
3A5+jeLE+PTZMMJMFmB1snOiSLcf0v+2I8DQalU3VwFD/CJSEy8yHNWExszvr8zTSXn/TGAFdT2J
JvgCgOEBBvyOHS1V62j5t1Wg/v8NVz2diGNbFaHlrIblxDZxkGRbvq+lMAeDMzi4ciFIRg3QNuZU
1i1wGVpVe0eEqIZpYk/x9BEZWpuQ3SGIFgmS97i3VpBHz2juyJlwyeVNcWMHbOCDmYdR0ZfRtg5a
Rx2pyYpM6hDGS6EAW2nPUY1lQtzahr1eR24uG0WLrZ/+w30LNk+HIdJSIgBWD+FbWogC7+BdSWE4
Ikq3nwLOOgRYXqNNXxTR+mX0YR08OrBKx4CD+zkOhgm5hz2d0MlNkGt0axeQ+87Geuh+LBcFp8P1
2HoR8+QWeyT4Yx4aLQuYxVjgq2VOZzS+hg/vqKRu7vtit95TulriEhvnpv0dYcj8NpHlk2f0SIRx
RK4mqEpraJdUa5jPwWFQHjsdYgSxpwAY6lJiaILifjTW2pnDWMPdrpLHs47f+Zt6Q3kFimSALmdl
z59xjy7UT0Vhs1aJYGRG/CNPMp23mxqi04KeLSV6aN+tIIv2Yhao6repE6DfchCLxViEY4XNOS4b
gnAeAwJbSMjcwH8yhj8hw8aCoKWIrZLAoqnnTT8gFLHkMyRxkGFl9MKEnuWgi7/Q5NaXJGvZZZq6
hyK5hQtFJtx0J6tiIUMVjI1Q6F3+E25CYD7nMtr8623V3iIBxWRZToByPYBR9ml99/79N81l3QBk
g1Xho6KW4P44WbToa78zIMng3/xqTJ4qtlrJTlOoBmJUJrle0fHhGbx/vgW+OeDcGsSuKO4H4/RC
67yvdEgBmNwNcW4D8ZAR2/opwcB6txXzhEmS7Anfh2F5HstHzfthUF9GlFWS3M7440prx9iX/fMQ
9dNpQFpgZzO7tfpdZBYayYiZH4UgJkEvlGWHciZn2lXU8HWy9IO7b/SSK3M12SUVaVn49QP0racm
/o3aoPHxOMd6lSAUJGgfs5eiHO1S27nqI9izL8ZbPHa1lHqo/ToPmX+smTWqG18tOdb85fE0H0EH
cyDHCoH8g+FmvrY/OAaCpaoFOp8hEK2cwrA0U9K8mRJmdjdc+GlfqGLOi4lTo6PPOWSl6pdvZ9zD
ROCeFibG/LbMKU5p7/Y4sAVt+11EUpC30Kln57JZ0fzZ40fUzX0U/Ov9SnsOeuksB4jLoIbVVFhm
N74vN6sHp6v+3jJRVEeARUnw8w9hqM5KPjPdAN9nHBbyPxemGl6M7YDPIjKln2GWSkVJhHoPVdqH
sLE4i5ii91gpkModkQXmeqFnSEYjH8DEllhLQTFK1OOCfYwtCOzDPq+spRksUJGP1YuBv4D8n9yC
5XA6Vl8n/evSWv4dy7HxAQ1pPmdwt+M9jGn2z7nE1CRRK5kF9gWSmZhTnCuZhq+40uG1/mT4OPIc
8NfAE8I6ZlYtELwX5NIy+bS09UTDvb5TsZ3wgAK+XIWghTh7cqj5DeZmqhJxm6fCFCGNPCDlOapm
p0MdvM43jcPMI7ztCJfabGKaw6D6WMcczZqutCu0c2yPfkIildYG08EyCxikU2rI6yx3noIp47D0
5VsIDiFVNBDeu4uWfMaOwhqq7rZ4cmjJjFT95g/m6HvXpw9C9dbTviLZfW3687LKxAt3CxlH0kbJ
02aP5TKYlRrxEkZUijtCvqj6plav9FoNLxwWVG6QTowAAcnSyXO5/whJsFfnaNw+S7bFRHjuDngG
PH0qI8uch7HZ3BTdPa0M5Dqu98UggV5jOSSflV/opoHftTvyB2AShj249qJcXboZ6ttB0aMFwxWF
TiSWggYlwwyM+2ZY0d0BdLVLj++T0j/Kb0Nh79rdMnG2fzXfNM44phXzE5Pv8sPctj0i5rnvA7zK
TkF9hSjfUmcfuG+7mLiUPo+HC1NeZ36akz1p4oAEqZA94u7fR4j/ts1W6dCKIueDANTb1x2/jL1e
cunsYjO7l6LzBljZoKSRv2kL6fgBO0IxZNhu68FWXLbGsIgThLkAsIw2tSZnPn65bj/LU9R/aLuq
hRIQlfrmk/SWepf457MrAo6Lxp7M/kMsnLB5Y4BJ/AvcWry5BCIfgOSbsqEvO4L1255RTrpbvbt8
0ykb9zTDfRxPox6qMeZPRUZ3uE7wwqsoLWkQCfHX756lyzS//N/zLz9pLclB00jIa2dG6jCesz+P
O4ugozMLXlmDg+E9ozrsOXFqu4oTISyCWb1NRJcdFtYFMC7VjlEnVc9XhKnLfUEpU1g00UF007el
yJc32YEkjplqdlgg2SFvvPIcQxRg4RjkwlhUgHATGE5yy+XJGGIO5STcbcS8oF/bwopugT8cD/Ah
ckqzQKjIQW3Vk8yHjOO81CQgRad5K4FDY0fzZqiw3qajcAWwI3RHNyMweFgeojobrVIG4uR8tWcQ
QWYkRcn5azt94YRXrvWRSATIEmXQ3VJS8KlsNwK8wvb4dPqDxrl73kt02INL7ntGVoqzqc258qGE
alYuUh5NnGS4UT0IhIV3IebXCB+a8G2lNHUrBxGDNpb34+kKfbacDqDd39T+vw16igo7SUnEQyRa
/zXuLNAw7oAVih5Zhv6R/ByvFiRm6EMxsYi31n/kVCm2d9T8C+pHQIjcgNu6hSm5vb0tWpZBQ4Nj
CXrW+W+zzGmmyhRYhWQuBP0kKyRkprxb3FNfmyJEja7j1SSNWuPSrHOb/I94KnatpDdn/UH1Soll
wAbeAMknndoeXpJ0oFuqM7Mw9KktnQ44px2p9jiuhHLe4PTGRe41lasT8DxGhlHuCWevyL5isGm7
vLHwgaELhwiCrv1On8UmxD9Ej7z12lK+9rEoZBuHhJSHJQ2uT04lfxTdUmnT3ddArhyHpaWcP8RT
6N2EGP8aNDVhwoBnZr4cKfGxjhzu9DQQYvkgTaA/iBOvxjGUHoX9O5rFDQSmKcNSR6b1kbSP/yZA
CT8jPvnGaHYIsdL9xXP+0jlkdYKbN/yzbB0si4E3Hdy27GujCUGfY3dMWZFeOStlQBzvYwzS6BnT
DCAp8/Z9MWWYv9tPKknl8MwsFIvozgFbhvabYxs8K8Crcko81oAljV6pZ6gSUF2iy/EJhxbbCZPC
HYtl0Fb8eVjiS4aiF6DyE/SLHujV/tKD6TdIA9EnJ9h4hm+WCa4CbLpj2l0ykPXBI9OUd+9t4uXZ
FaIUrSa2mjPFIICOg4OcJoahy5ID/KCwlMtPyvV26KVibI2nh/DjaYrgPb4rpco6OWYRs7Gh3Iww
xl+FErKwR6YCwnoJDS2Ritke2ERnQsCsjKQptdehtwGlUEeb/sKMhcFgZjxxHrKCnyEkUge1HW5j
0J41Bs9PymfiwuwbxU37jHckUZp5/kY7xlXoNUMwJFKnKhjyuX0y9/JllrlCuAk8zkgRYGTE/noG
CEHhviIv+EDLwEoa7FolRJsDAe81YgR3uY/32gmnhFHK+y06kCYsR/WKUOyoswQ4Ritdx2w2ciD9
dmBxP0+4Z/U6RnA9trhFWuLe73wfoRzFSGWXQhLOuDIVbUPYxq9ElSk6YcNMgAZMK1rR0INCCPoO
M+ojGkDblQhb1U5as9M6JuAFyqnASWtc9sJIq8PVc6G+9rj3g2LhnccD1zNab/AlH0cTXVe0vowL
K5Ulysxg7bicf7pIVqxV+vfE3tTmADbkkTEgo+K44AipAxQ6FR2IQO0F/f061ZrdqovvEuiyyqew
Bvn3GiwudKyJLFvdKa725ajsT15S+JSzUcXJp5d/FNTVyx+rrhxLosEuiS0TogonUPRLXEKFxYFg
im+LAGxY5dWlcm078AbxXsQKKC8s4bu0fVJ9wbgjGPfy2CWnxh10vdUelkkoQ1u1wjWpoclsGaXT
41h6yoCuxBVThx/HmXEjWiUUvGt41UP/f3kfuaG4neQcN4Wzn3m6ZUs2LJ5sUIPD7Qwv3QSBguoV
T/KcJss4tVkZkZnN9bfIiVZXYbNvl1LfvaQceY3mvlLx0uHt7/81nKVIubtxgRXSkvZiqo6VPRva
0riXRxjmVd1XEeQ4IkxnQpTIsQFUmv+TXERugEepK35p25QCdZbTXS0Cgc4eAVLUjLu298csyEh1
3d5I/VsYGz79/7piau14w2MOA7QudxhbuRWz29fwUSW3GDpSvtBwGugaJlzpyyRpK0i7Xh7T2kTe
mLCVqnzL90xJpEnKsaRohdlfH4vkZkM6HIQ+5wnl8iUM2ZlkLd129/5G/BGxhuyCujXlXMURaaQn
qPsHI8w9PswMJ6G1zCCSVqMYB1HmzL/kM7cDvf3bMlrhK/83RotQ8dBeN3q+Oa0owI0/V+NJ9x/n
LilBcrsqh7K7EYvv2zQNedmB4tPwvnpWgByJFxnL9orFVgstgFomWqJ9uJHUqZ2Nn8d3KEb9ujdc
RgVqEA81Dm5ROIzbTPui9KyEzeZTHmjXsagrZ3+vQPV0ucGfkNqH9RItIsiXUdQsgEi8zaQ3ox7N
LShWwN9MjwZ4Cm44XIQGMd2W7nl2v4oSgVyPF1o63DL85rEtc3UiW8+Iy3fneHZJ75MGZFCfvWQM
o1spieBJeg1ilP9OtW3JTQDnf6lMr6jf6k6bRcv0eurYRwEh0aWHNuaTnSBaHwImKQz3QKn8IF2V
ya5bGh3oSWM1HYwpkuujeWZOOue8F7WpcmqB48UVOipqdpEkAz+YzZf9duDaB9BuyJ83w05QSU9L
dUhOwuxjbpLKiyrdqI02ClVxrSgMOd0zdbWgWcZcsgRD1l+u3TWfUwCt6rBrpkhaEMOUHCQP03cW
O1T7XnTb6Z6ynjPNDZ0E10wYuqSPxO3OfJqaSO+CaHfagu9W1tp7mt621CWoScV7Mfhnn9iqVS64
a6Oo1yia0a4YMUWVZifLlXRs/ts4UYk8rvkVIYKkR2PRlv53ka7g7XtF5xZGO6ThxLO3xZA4Ikty
h8V6day14YhtndBDpqshYqgyzfIeCSIhotKNwC6Sq1+kPcfoogjVyWt51VvknvWYk14IS4oLKwAF
XpjBQzsshu/Vshq9rmjQJvWOCRBl6qVeL0tKSsmyngGnvfisJ50xEb6bEOtDWb4UNX67PY6M82Zr
DO9COwJdOWlmXKl3hL2J7sh15mUOqXFOdKQUSEwBPpdnczn7BDTkVTwUUdHTn53INdS5tJMEWS95
w3Oa8UbKStbD65ELCJ5+rOdBDLzfjbE7XkJaAXcrH38Q22Lw1tpNkz19GadhcRVg9dz3zhFlJF7T
63PgGNlqMy0cGUinG72IuR0fyscvfdo1wU//Rxlg1Jp5GHUCBE8dfPJilomnSDmIoyac66xWqi/d
OE1JFdzLnXv8oi5aPTQGkzqH6bzd4wuBNFW0WybwrXTyZAy97onDEi2+jHyGQJxZwcB1Jad44HuQ
0wpSJz88lpWlVEiHkg5aRIVsL4YVInSNxvB7RQ98pWld71duQnteplluZgBMuz/WCcplyDf2AvzL
VS0BiW8a+cirPd7V2g/G+op6TvP9JV7BIXtJsyhxuxcu4gZYSeqSuYxI81DJZYIXjKiiPy4NJhGj
Xpo5aH5/BD+agcGEbv37QafB6z33mtJmw3DiOmJsEuFhDuJze+unhbg+QV/ZIu1CYm/NCNS+q6X3
PYKFYfOvwpBbDgZDQDaUFMe7x4oiyQN4PqwA/qQEqWkvi3WQdOfAuDuLK80trHtHe4wa/YAVt7ed
7Va/nkdtRVMZu8Q3FG9U9oDrypA5ROq0fKKkpPxPkhRBW1Vijq+BpsNywIZ/Pj/Q7M/h/xiRCnUj
4ktRmbu+g5zQYUM3lGSpMzIF0Ty23d6KNNAR5DytdF9VCcmiQWG0RMJZKtlIRHVPvHt/nEWU3Ml6
g2mLwOCx71y1WtpODV+4gc5a+IUGtRLjFc6/mHr1LImw/l0PhnyaKuyfEi24m5J/zvSkcetZkQEX
oI0uSLTTP4X1lQR9bbXTyWeqfbQxac1jvxclVYtm+msK+nQUk8aF/gCEO7vAh3DbnFUl6qpNo05u
9RWWpCQzovn4j6snEqk13/ShlcuUBxtiMPRBOqDqsqoX3RzNORXi3h/8xgRtqSG3wDQ7hAD7OWza
vxDGN4SzOqKlCM6qTJ8M+CHdHRH77bJXUh46UCKxHM1BCIku8ytpLPg8LdxOMXmVDkuU/TjRkZox
jcsIStEHEcLfzNzKkPbQteB55qirvENNWo2Qw62RYaP+IEW1LWulJ7lTXjUez8xolAwizjeTTJ1G
s9xTw+I5iuvBU5i66VCyJe1Ut6QrotPCe+cqGd4F1ZNv64SnPv13afBSERu0ToMiwBG1Jy+ACF3s
tbzxPtKP88/zPUM5+oBYQsqdYXsTIQd0kWKtAk90PfH6hxagLflROukmTOsRtD+0MoDYtX5V8rpf
n9CHpwF9SuJyHwbg3ZZNRH0jDm6aHhJDPoPOHUYLi+59zIg+Je/3YVSRhQH0FVvkNxJ3dkGfX2qR
VWhbStIBySg+2wJQRtr1M30yZe4U5mt/IaHze1q08nCNq039gNGVdjwGRVbwB5C+8BWbll8BLrBc
CHGw26z/btj/3hzUVxhi/KsGjmixLfra5v67AQ6Ke8fWbk8J14HfblfA+z9AY3ZXVQzlhxD8S4On
opf9U5u8LmQQaczRjddTzZmYE7URJyD/q5OYvYkRfaA6gThcFTydP7DFJi6c3rdxPmap8HZe+/iA
RucdBwODugDFbxBqT8mski1wBrMorR3/ZHIDeevFU4BKqk4go+62gMkWH9V+b9jxI89HqZxdF35L
ncWF1fmTXEx2FTqCkdmw+ioYem0BgCGZNuUbR5eXfY8s9ydAfEwGWsUC12EUdGT+Z7ExASE9MQym
aWpS20Ljn/RGGKCHhOKWCSQFU0OoXxEIRfxbwlSdk1mdReTrUQAHKH6fyf2l1pfVnLcKFypH/56f
u++4topZKqz1eMcXNZmI5tBZHcMGNMo/NGQ0SY0LJtnRhdnDeCFmnNsZi8kZ6LKoMRrhN22hFRRH
nlFP/UwLhjgpPfLt312+5bs8+aBf+/5NARFm0I9ALtzJy66Lga1bJkENJV9hs/40vUEgz/VRuanj
nAkyMvqK58S7qFAy5U8OauBKBt0uk8za5FchNjTJcV+POo01E113y5k+oPsKFE39Z3g1BD7iRKZb
2uO2onymMi6hxWgqvdXPE3YpBZHq82HtfsmAl8E4q9cdUcCyMTsXwIFU/Pb47wezGw6iunpQnB6o
DLl283sTsfV9j4D6W8iCLjUXZxOQ3LkDRHgh45jBWBpCE6xg3kZza8apQNZrsAYgPHgMXZOLR3O7
Gibeh4ZDUtdmq3RUIB/azklVo29zwmTnIaX1atelvko5HpQiaVFkIilm3JdaFfmQ0V8uAwjcdtqK
BQU9dFUeZyGoQMi32ZxGF2LDULfmXpKZsOT6Z4dDjHaCkmmKp/8XlFTVr+QVYFjjE2ewWZKSrJ2c
66XBwhdX2IA8UZCK/uL031HDqXkzy+wRtiYkbsrWQKpx0/w5Xmxuh3wH5lZ9QNY1yYf4C1OR5GK8
eZosqG29BXyYCcgaaNpf8MDWyDQnyiXeJxBJmRpSdX9cQ324i1Jp6ei1NRmAmT2rf3/H2RKb9tpb
AtI63gtDMq1r5XQS0wchUf3gVvarKIfic7SjZ1D1RKn+wJCnodiH5SdQSN5Y76+Hzn3oXKYZuGdZ
2EPesXvVt9a97nyYhdSe3u80Rgc8RBVv9JRAIB5nC2zCeP2QFFvr3OTNkPqWOK72NhEfSkTRUg/H
zgRnGC58Cs0Pgwx3NGpNJi5BwfQipbI/NZI7UvC6QKCvMl234AHCxWHCpcs6hFoLMvD4NUajIy2K
hzRY8mpdMBwU9fY9Epr3xDdHWg5d0xlV0gusBv59za/OSicGLL1fr19NOW0z+i1c3C2bIWub6ds0
E+q+h8B+cExlw+qqLLBQGFFcYCSOn8RVsXL52Q9pF6ODuO2Ap1z3Wcm8euNniaz5hFm8JceHhEFk
REy0x1MXb7/Eqz66XnYwWV6kppBGdqYFdEsh6sTmaF4jU8+LVUa0ocCiO9Y0RR9B4JEtAhbvs4Vu
3u4MYcYoR0WLlsydt/rusVzRzxxdyDmQF/tIEyrfDQ43lP2lVamb8vrKtjTT1+SQ3JtRvmXwKXcU
nD/o/Suxnujf1+H/gNoqzRiID/WD7yThLnBXdumPw9h89DS9Au5S+NhwPirDFN2EcKhBqbs3Geu5
TkPtfSORCwYylGwKIj4RMZSNi6e2W3yGJauANbCIyf0bCkwGcxqq8c0miUxWYdJh//uGyoSl7QYB
JQpoLdgJJxnKfY8Z92+DXzc5FpmKZ4HMNcWC34MelL8HVek+NPJxemsUVOoYQkbB6tHGcb3WWzcj
LFRxIuSfM/aQxHIwSgvYevmPKEqm8QhU2D89oP8TJDAJnZec3Mn7mjdCfVwZQwBQUTD2B27yFrmP
PPElJLOe/1p7hu4h1YsQltz+lIPX8pOcrrxmW1E2rLjkD1DjpFJpxRU/JFT8MnG4zxYRGHMhEZjI
cQfCO2oRhXMaDcZ0ejvbihxgqq3saE9iM656CgOkbRZWHk/ZAb48Nd8dGhJwrlVPdKhrR0Q4aGKD
zAt7eYcENiYB/DJvJEk/SEO9d7cIrrQPvG04PhfjJOa6FK9m5DJleSCVVrMv/SdjmxW2Q7MRoCbu
zYEIBKzJVDFZrf43vQ3tRhpQ8GLv+hhjQYJ+DaHwaxoITpMCMnZAQ5F+xvJwDKvAKyFhNaHBANPE
og8NsMqbbkIGezpjaSVrmyEctwwTmWnr/ktJpSGGxJRslbMKN9/tlCo+awkeOmv2JnxGFtZDRo8T
VozSNA8Bstp0yGP25KZ0TmmwWF2ircSBrerx1upYgiFbo3dophJqbWm8SS5EuhZSTr+Rxf0kyjR/
+d1HCB9RRMw+KBho1Gv0Lsp110gjhXLivlQf1woz23BlYlWBLCt9AbNDpvTvDV9vBjYIEZq6GdfU
Yv1rxOUyDlj36TFP1aTuPaAmosNt24Fxi/avXFydDdnD0yY08yK0CDz7RPis+kYSrQ9+H62GSqEB
KkXHamxcmdgGtbtRfrPaRuUkl++jtTtekB8sE8hpib3i13acU/eo5a4+NoA0yc1LG1DUg2TjPRlh
3UknQWbOliqOeq2xxaBt3RzHiyG9uHCD/vxAvn2oI4h/oT8t4QNaAdG0dw900U174mShhKZ+Wy3Q
YpSLE1e/3K2Ap/j9L+0UANcQ0k+IVQO1WuR6SIml/6zfBBGT4ECGXt/eoDxMSze5bMSQZUS5ImnW
ORgT+OuTvTzmfrBfNiCZfcU7G2z4PIUzjZQ1TdPOrRxzkT3bf1LLTcjsvdPMeFEYnlXal4/9AbmK
VtG6HcX6E4o3nl2f27YlT7Z6zKUwLhSAE9yYb8PTI/iQtRwLvJfe1bRWAy16wwJU6vq9oi5j5pif
brT3tutABUEfLmOhG6UudOn2yeg9RQJRtBGWVBtMoffsrwA++6Km8ZiBD/LTXdhGZUsB6n0x8hRP
32YgGDOGBF6yj138m+Tn7aixhdbkjJhyEArpPNWCfByjyjqBBC8AJTlgaqZTyZt6/79T3L/vl0/+
CrmSKaPrBRD0+YAHsqDrwpleSvp67i5uf0W/gw48e6dsAgJ8z8DFMRlwydqOTi/dGqbUPze7E6XO
icjDtP42zWo07WbjsLmkYBSIIxvcZq4LYqvgOH8P2RwMB9u6j5C1e1YjnJFkqqVba8na8kvcJSnf
/1QbqnirMhWwR3v6vYgixbAndlqDnPQfT8+Lf6hrQoqkHn7/IXd/b6sVt9vcj2RKeffNv7+m6zFJ
M2EP7VazpU6YmzHeu826NonNiskNs3XUa5ZCL6mwJkYZc6tHhIAT24CE4JQfRV8lixIbJSnaq2FF
+kRX7KLPkp583ib0Lgef1hkGZJ4XOBezz7AO+t8Ve2uRVkcZb0pEOpqAqrDq3imVOnYNg13OsvFv
fGhySsCFllBmusa1dywb4U1nF/mDwcOcZp3sjr0nA40PotPuvW0TekGWUAwPW3SQiXsDv9wqxwNk
qfK+9HrIGqhHdrUpndnajUCVKP7P/RKdRibS0WWh5g/muYBDDkH4oDfcK+oyuRRAWwdmpplRdME7
Mp4F6WvzQpQYeyKO5/ijg6IoxporB9moxvcd2UrSHA5NuenUtBQCBbXIy7/AOTcnaB9z/TaZHrVD
IRiiHBZyWnM1syCa9K+LXbhmuymMuanOGonpaFQsD34jFUmcIkX+qlZWeR2FSd2LW3ZWAgYb/oih
xCU19tGinuR3t90Cd9m7n3sQnMzJIsiQrNjoWaOlNthmZyIMj6QgC89Zk24/Ru7Pqgf+CjwHdrhp
MHvTeRZb31qXgUDVSoDKDI+ccfDFFG44G3Pn1j/0R3ayAR8AH4g+smXzlxreGV/Z4mhwQ03GxAph
Qk/rv6gLawWGlyUWXbX0/YUD311mcwJR2uc0+3/sYZgyLvKJ0tdFGDrXifz7cTZyCpTqw8FpHWRz
IhdS1ZfguQ3ZI+JvR8foaWqEXUIBEcmqNUD0NC4DWy9y6aE+N7LiAzy4mB178kbKqx65Ig3akJmb
TUiNzV1ZfjFWqHuSDB/F6DhJIL9NshiX/mrNLpv7QjMJUxdQJd1HeLBwuwMYAu1Onc2KRTnktL48
JrHSxp7uPNVGiavGytWoNwIgDH31kePyqAqmpUPxSfFWVJxJUrBq5YA4qIvRiZyjL77TDt3oGDLD
fIQrueSK/RfTGE3bFy2aug4jlHkqromEOoyB0tBNOnaVif94Lxz/tEfqbcnPKna16RlBoa/XeU0x
pjQogJ4Waxow8ESOsW/kCCopeyo0S/SbdljV8p8yj32KNKY74uPjsXuJqhChITm+dJhM4xFGVyyS
ofQoYsNqijwEGKq91Emfr2ZUSxjRJe6KCNeuUOo0c+DD6Vx1h6uKQWuEBq2njfC31nsm3EWlil8f
MFUKHeOlfp2lftRZfIk03Pe4JG0d7fFWMIO0SmS1su5MfMyukwvhdQBxX56+C1YtJv+t0BK5Yvas
6CQEPHQ3fqz0OiEzXdC22ii2w9kuDrxMMFNtOxblWbkB5S/aTVCJJA0AH1HRvNpIszNWv2ifJP3p
vIx+Mb66Aq3Kcim8Q7X1+/ybt7t+0ww04R4JYlQsbXvJw9b3DZPlU73bkn+v1T4YzF+VKIpnDzJr
ZUoCWMOrdcAfLFPuu+br31N6478rbioz/JpwkTZ1hyvAW5aDeVtJZYiwQtCIfXkA3fA01e2Lv/Po
B5bCT5d4kLNKXtjtQ7T78kwvPtStRaksxh2QGety+8EyjIIfcJzPrMYOGmUHeBZD0cCu8nLnszdK
9ea7ZtfQP98d+fI75pXh2abG+V7F0gLNKcnRSm0q/EcFGxHIYwhubmHoqgFfROB05pg5DatZre66
VT+ammRd2LDZFW4LdMnEsHp5mKF4lIrjJhQnvj5JRVoxZB5tQ6U77x5uXEz9lc4fW8FEmzJ6oGWS
wcSA6P31y1StfCzNuZioQwk9Y6u8aRxXzxwp2mx0o5ho6SDuflWHdL6SO5ShYYRS/JsHgdtg9tC4
8tU6bAkDPsdUOKpCh0A9CXQyHc8YukOqMJdvrj5KjKZfdbUF+sKUtOIHkUzASCwrN8QB36/jNM4/
/Ctp7s0fI8G+10EkYt5wpyzGfSJ7uHBEzlYtn2KZMkuunrCavtmBx3StureyQ9KVPSS6OHTWrZ+t
slzzv5h4IdYCPBojEE99TWV0qgcsvzXCSM/3kGnl7frTuTNK4melI9B1KTycLwUlar/TlNVkILlS
4ezQNdCTUEe/vVwvgLj/HL4lnrBhonDCQhUZm2o9yeeDVx74SWjIp7fz/irCH+sxYV95O/w8qR0m
ZXTEYOUBZNAV9HMnfR25YSxVkAoT/poj79veEko2xsOnENaP8Rum886cUtUtJgpZCFJGZt9eePBW
VaohfQqeCD8vooiDJGJxVqk1y8+fGZPekvO/Bf6jaWB+3K2ajNsL7Gs4kuCPDyJnUKTWdcIW9f+X
ZoYfbFsMBmZ20lZxL29WH7Akg+SHEnB5Ivc4g0YRkf6n+Onh/kIvqRhmDwkRiE95p+BtUGWJXtYJ
S7E8RU0Sgtjm2+cx/t3RRYp78wyLdWE4i9eDxMeHRRBtMQerNmy8o5/rBae87gDJFgwY5Pk75848
gc2bqxba2io02tVr1LhDBD8ipLm/DPezMBm7q5xIJWmR62A50sX6KOAxUdDyAgdQNMkFxzJBllal
/A25RgYhhERM69S3XhBqJ7bLoV0TNAjf2kcUhuIkJTGW6pTggWfB4nxVkAl5BCSGP9stKBaFZLhv
Pir+56aksAvuXDTu5NQ+VUfYipvUamab9OGB3m01kt0YevPoAPPTg25GWmc9UIIqKY9biLhMxW9M
Sim0b534ppt11ahQ4Ve7CKUUP5QISkf0zIWBaCwQ3B9Ka7Pe1QcA8XHynSx3++wUQigjERdUkqh3
R0+R7aoVZsJgGW0FuAPG2OW0fUVTODr8AEICok7mCkzd9b+5xPTFPJLPiHEhVFTwj9OuLm147DSc
d2MX8KgbiN+PT82p532YZO2BxVqQEDmSkvgO/GeQbflohGwrOY/cKo/pHMEspPMyWOz8yOKnSR5c
prUXPQmKJRBcuVUCSECb8WCEnQMDwhWFSauSmTY+CACwy/KHv0/gvu3UGZ+b+lrAprP1hoxnN2Ym
OCvIlL6M/JlDL2c25pUhnPOH23sX5PlkSnr1Ys7tCG4Bd+CG5UAAucR8tsD3OdR9sE+bvre0J7nW
ExWNZ4b3jw4jo8L3LdUbAdhVf0w41PymkzFKeqtFFUiRTXlHQri1LLYwHV1/MT3a/+bPy5VJ2s5J
dJAII7sXkp2IaoWaO+/UIvQEUpJCpP6vstASJw2rsa6kejP3R6XQ3ht7XGgyWDFhYBIMCGnlJkLi
UiZuloIcYvojwVAulw4fAWrD7hjDbFbXxxyy0BYD8rxX2xG/0c1Vmi750uj0g4J5l7hQj46LpmvW
QUczN82UXGot4ta352nV0mHu60XDZGxwRweVp3mC+mzZpl2SG6afqPBtjzBGD1Q8vB7amO/LOABd
ImhqxdeT5PRixH2oIv3Lq+Gxy6HrzpJRi3AM/uAaiBDlr8uSaqWfyT4hJqVXt9r31ZW34FOPbWb5
thZxumnwWQnP9ru+ugCOjNgI/51/+SBy1fw3BDS2tzW4lP9cP9UGhmazyFiVoKDjLu5dAw/n+x3i
UTeka4NNcGvImSw0YJ8iCc1Hwozicfbh75kJv9J8p7775xDGTUYq4We98vhP6vzpjCJ0MF5YLKVZ
sXjGq3dNKtexAi4CNHSYGBbzq1vUwxU7atfpDAyD+c4jGBEKT/XABsKfqk/8dDT+zLpjhPGbvTTK
XBJCW31ZXnzZuvefygr8K3HUxQCPLz2QhO8NBOfQBNOE1BRO2D3EnpaMMlcDq1ceOWGARvc9+f22
WzPjBZ4n9RzOhybJtKx2Q5aYiH38QtfBC8hff5JGXTJQRp9SmxuvlyrAZ7UdAEMoeFYFWVH7nyxG
V9/oPp8Owcn0ua5YMzVhVF2eOCJnSig/ca17pMqnWguzEgNbiXlD/biwTmVgn49Zx6TPDwgNxE74
yoAUky/YYzm9uA3xZCYBDIs9d4AEu5NZe52i3llwgAoRsooGHuFJapTYqdFq8u8Za4qdHhpcOEy1
1gQbUPnPWLX48PuwcTxp3HL12rJhqF/amuRblb6wfyg8jqfZlUcTVojdmAZnFSd/Uy5MtnDMot/D
SvV4HHL+NO8AfCMS0YYyNbKgpq6PE8XNjeVFh7uZWoEJ+gvtG0EWTgVYDpATtmyvuvPedKGVbwob
+9aS4SZbWd6+n6B2bvzpbuyiNrdd8O5WeogVCcoIa9+uizy/UsDWz+afNzzx/VK6XK70kp9xTdDM
CGGOF2aIOfRGdrXR3u8k9pRi8Cwcxm5bvZgB02BpLnDObagtowWOlK+48Kmi4pvIOdA8K2IE4CAz
7ohfLciu7R+Xj7aakk1AUP7a19MkOxf6Dc6kdBFLW0dG1xDDNkgYE4I1YBLYH6qciA4IyR+DMF89
3u3Lp8VtYJDmx6jqCDpaESaVuGnbrKJFTlYQNR5YvyErGw356mZQnmm14q+nZlWnsxqRiHquirn1
56on0ujykSRIwZQkRCbO8KNK5UNjAJEH9S1leLFpteOjp/Zzb7xHDPyaN2MkZWCSjDmaIYgZHeUh
ObG+QEkUadicX5pVd5HvGLkFhZXqXSdIl/bT2+71JlutE6khvW2QBHGLK/AlHEJ24rANqZEix8oB
r/qxrDpL1OffuqJ0Di/PjGYAoaOGb3i1czzcQwvblwqFfHtbBQzNTuyfay7nmy5olE+8DEYflWJh
dm0gqAzo7yNkFTNY6VOVSDs5oH5oyEHGbUhveMQTJYGK8ef/t1QRfVQ/HSej1iTtsQo18wqLsC1a
sG+0D2mGcEkD2c5dl+1uRzK9Mk4ZC2LqgcETfzWjb9jXRFJ9pDgFc1NA3agft67QL8fHNoDLxBDj
WcfNhlwyTsx4POqK79STGTfEjOiEucrKzwvS+XiYU+Tu+czBBiIPqyi+4gmnr87EcitMVTASsmSQ
mfg+yPvbD0QRoEY3SuLKsf49Ef3Rvr8e2mXEH9UwlDzviTNNkMOqC9W2aGgxA28ky23c7E4BVhYM
259hgYprxMWmSdzewiAIgYvZD1lr7Z4VpLEYkInUVO0fWZ5MENlstxfOZH+TRvAT69lcVsHt+Lux
h0/fiGEIdPqOGlduEJBSlsaQdsgr+HU3Q1owz20VyQ99LpDm+XOGmmxzinm8upvF/BBKhXn4s2pu
X6o87Rjt8L2xQcEzP5gRPUm14ra25dCHQRQN7Nni7YphqLz06BMNsO7tgjo6QW+zbUbJZk9ZOGYl
rodm0MUI/+mpbuEMi7DnC+II5mCaYIJQbbVpiSDdEzpw5b+65OSuscrjksRXohROk76BpsinZdCx
11Qd8Ss6AwzWnjJhHi/EKxCcEbPludv3NdQbnK4YLtuRZkxNOtJAe8Q15ddH+ysK9Hi8tr8SgDLs
nokwpRHeMkrdzYl2CsuZW0s4XidHfoSV9DJ6+Z8pRoet2V1duwWCikJZ1LxAYw1Uq9FhOW1Cl6Ws
aZmwBvGBtaYoGxs/r9rMxSDHC5PEy62Jfimn/j0YlVwOSF4fbqBkYxtfoScO4VQxvj5p9xWXdAvQ
mOyEoXhBXd+pkWp9QP8y9repXt6ZaPiv/CeazuOZIZi4OF1WcaCH9oFm7dY5EglrGzFhnVQxd1Rc
Cyi9R4iH3S1goVfoVCnmaXOH0QBJ5HUxs8PS0/WsReuqOBQaJzgc5zciaO8nFw05Dw6spdcWAvIP
uKAfk0jlHfuFPIfPx/dwHf15V0Pu5ruwuVGRB//y2g8KPhoB33Rf0YEZ5Z6jNYVG6HKHjEJkMFyM
JkuJXcqTbZImkux63LQAaI9YZaYGESLKY9J9HgFEP/5t7fmcKuXcBEuEQXLfdlVsh9wkyywJ7mGz
Qgjms89wfJMsM+OPYRngHYZr/j6GIxyEaCMwHEbgVoEsgf7yshP/av0NEpbuM1bYdwBca9OLpoKe
6fz4HTX0Iuy+oz9vRGWziJ0cYux3Ed3l54bW8qBU8gAaB97LFL4wiZOfMozNGQEOXM7W6MmcHJtJ
0lOlHh4m5GQU2STBsXv7Rl59FToGJ5LSkLehp0NG144mjkEY+TP5GWA6LDosvCjqaGc8V6QxXJcp
YnxCwqb+Ay+oDGZnsMXTinAnKx5kMG/2YhitBTJ83qAcqcObqMCLR0xYBxhNNukvNDbXGHjx2Qa4
fSlFz51Q8ruSg0b7amyeUdCYBCv052KpJcd1eALCUqXOOGQxDiV9zYdYcCQljApC+KHZm6gxaokx
cSPpuCL0NliQjqP9sMTYRPuwcunFxS9H7phEz68ni5AQPbw3/t9h2y3t1YKksFsrEzvLosSgc4L6
SjLk1wIz/bMCcbfo9gt7QcAV1pRqJP3Zv0rodM7JZ4vhmE66Jyyhaz1n63Ty9zEshNnZcQv/3Yqf
3+oOOCoN5jbL6UPdwNLQ+p4BNcXz6uUHMOIGEyY6TLHRydUniZ7rzljJRjWn6i2KnGJlOYT2O+YO
v4QDuJg59iIlZCR+sY0ox0m1KAhKwoArnSxvF6uef8UhaAGe+WD7IBrzZGcndVLrEl6sqlHE0W41
5JVU9L/662KngO2HNifpGfEFTyWBXjiAr4vyKU7q9z4PVevMbch6DgHnANp2G/blOb42cfLqKk+6
25fj6gEWMSJmW5KQuIIITLin5XK2aLPiBhvS1FZV2iR6wLFGmIqo3P78t3aQDlIZ6kNF9D3T8FVt
mrh/fcaVwjIY31KuEz/Me3MbBeaM+B8hDTG6Ev+R3yyODrHBxJu36/FZt1nxRoa57rm55SOZo6wD
ki5FeKBa3PI4SzBPyvAz+ar3P6SwlE1jxijsUo1czk1RKsj5HOhXmA9z58WhT16S0xhdck4kiWE4
AtFTTgc2oZskKdM2StWzBvj98UnWSjsXMSXnaatKdrlEcJiMTDzLkeiUPO4hKQYtRirQ0YOaooHw
25aaEsyAf2vw02IDfVg2qwKj/DTlZxgBDYLgwodAv1jwzPJ6SWFyg3Abd4kyi8O4X3W5gukjIo9d
GbNh+o59CWjbtDwndho6EPgv6GmHMLihiUg8s+OqAAMwlvRHvFbXHzW18ToRx2Tzw28ICrorgMy3
eS7E+BGL/by70kPWNA8S16QQ2BmLUCqj9d8iN8ftQjRZxA21E0hJRCZ6EpRrOZSuQS/jZtyf9Zks
TygZjUZkSwtcgWCqrLaxBbeFERutl8INN/30BR1Hfz6A6IbZEg8Acykuj3NIufv/ZVmJgAaMLbr5
UXTqHBPDBDPN7UFno6Cx5u0uZl+j2F483GoXm0RzCspNSW+rckVRU2nKrB1zQarBjsL8//Mang5n
nnQR/FW6Q+dgcYJVmh3VBO1Wha3S2IGY3DuDi5F6e+/kjICD+J01EMO8j2wZWXrcKO/0fLWbC92q
oXRiH2/fThDSS6V+bJBHJkKxzhS6mu6xCwZDudAIthcoEjY224JoI9vsnEV6e24ZCLJ3AoVWTlT7
F0lbVjudxElNkGIP0kMOYrrl5qC78F+aTRUZPGZVV3Cl4/VY7TQafdZ5VI1C6pFSBOwlAVAVcTCk
7a8GpEMQRczJrVUmlB0JyN31AaOogQM38tUwNFZIy5GzGzmeZGWsqT2vFRgxu+z7bTUt70dAuA1M
pTBhYL40b7ZhgXhxN1aU4/Y33+8KfP/EACnsCMitw0i+c9PR7NOHK9KmLht5uci0jh0mpExHl+Xf
JFjjotsmQWhi4vQCK3ctD/XF6x9mYKJX2eLwLMIRAuJs3PEzqlgajf+mID2U8DuMP55rRx6n5dL3
4a9ZtKF0frtYJ+fHq5gtmXaC0lmSvWKo2X+g8IpafD02qVWYr6dNV/oXKA5qnXmzqZLE+w4A/xkj
JVjHHyc8UhyalPs2Z8Fn0xEw+L87kP6Hq45sTUxBV5rdYGToYmROoQEIOBUZULezs3Lz7BdHbrJc
TrRhX1L1++W+xbQucVEnbken74wY4N+zpoMrWouzfmbdtSnJlFPjDClw1oNeElF+6QxWVfbYqysB
EvsLySwpf6tJGVJjQjD0250tolpOrddSrIzqOgAw3Asaxti9kxYaO76pWpnUlzl2qLv4IZd7vJlg
jkox3atKyiVE2cU3jPIdtQfG3p5zlCoVdEazYAvJgxap9+A6LaKgTIaNBpg1Qp1wnHpW0fsfZo/R
Vw1LowDP2CrhVlFgMwQNhFFuipLEk0obHUvQALgJzpfABC0pMbVhgu0vA04McM5FPMcUsUiCcDa1
ZIKgzH/D5BFzZP0LRdLvF6C6A8Maf1MhHzqEPJkBwNgqr+UvZs4Pi8WtiDnZ3svydBklbGS7MWun
LyAcKbO+GvWEPg0rAErQQ02B1R6M3X4FWxxPtsaRkJiCFSobbfkJXkpPXB5y7aCtnq+WNdBIjkeb
E1tImUegVGdGhP8r21By51PCXIiIF6m2w/70kKdL44MOPbUPakyZ2GzfhS3gpBPmKxYeoo2dedHt
E4QLWeYIxgMo+uSzL0nRCa/UYJlVgmz+HUEF62lJwdDdGikg1EoPcls5Kyo8GSyoW+ItZiUTOYSM
RiZtZX5ah1U4YaVx8ZZkTaj2Ll7vwX6055e/ZzclBuHKpXr+WWSZ56WUM1dmMPzS8lY+zYCvqmH+
X7LgRXPHNTUUK9LCXwTMbPJg8El9zWBXRe9881e7PlzvCOJOE09bIkBnGwJzhI4saLCZ/Qj6uAAp
pXtGP4dF/0yxsVub6Z5VUr28kGjxoNF+6B4pysKrJsrJFHMQmlU3TRCl2GByeUsXabe6z1MyKZ3y
Fdi9m9nVjAEAlhZpyJZmOpDEDQpNO3AVjxHsPrKE0ybt927RfaEx/SU/p8MV7w2HtJtJd/73YMc6
1jmluLg0djRutxFdC0mrhIGNgb0QNRfG5AuNDkPBV0A8+e505qIXiE9GQyPifIxkT+n3B5pWBSxb
on+Kr9xHxiQSwokVWancE3S6pYRrAdHPygniAsb8YI1WKcS1Vu3TMmSxywAgbWl5Fbl+xLJumW+1
o/7w0tI0a2NCAHKy9pU+AqcysU7FUNUMEPy4bnyXbeA1l85KsMPDNUGio5HgTHh2UefAjBWP2TIl
nOp3pXLViRc+MhypBYfcHmiM72Y7HnsMDFxT4swtk0TtM3Hk3ZFJaGwvA4m80xCcQFLV+lGBHSOK
Ooq9XMajGnrqkTC6MylYPpDdUb88rMmYvQxKdutYeLeU9zw007r7agqI31RdTniE4Qdw3SAz5VJW
GA9CR52+pp64AMeSJUbSNl8ttjkvRt3APkZ0C9jSlWNofPTIUnWwuV/lmbbT8tavzKd0WZYNqN7Z
U3aKctD5FSbF9xhwPB/OjZ+r7tWyeH6m+V7j5nF1Zo4XUXEWGc+IbnQRLA6WCo7qKCPLI5trU7FX
n7xhb30hGlZDTnjQmYcug8Ett9SOVF4+nbs+/YsUGVob/6a7Eny973V3eJQTNtlrJk00Nd4qFG/X
o3s0Jz34riieG0W+gXoHSum8aOsXvdgAtVFLdiZ5Trh7RZ6TptIgMO/24HKAZn4Y+FYRMT1tx6lR
q7Yhcb/N7EDUNZIFfn6ix1xC+vAQBMlYYhlWl9GpdaugD+Q0MgVUwqN7N+v1grEAHzsz+nTT1lMC
eGzZsjZMy0glaFylwJbZ82JackfXBBaKdgc/IvdhsDtXh4e4ac5E5BDk6595VYyGTtzwcZx3OoBk
0f5ZN6ihDbJzHbnHCBErExVKlEvuugE4gn1crd61iPZhstwXJ7i0aR50bvgso7RL7N6jpeQdZTFW
2sJTK9N8gvTiNTCYXvkf0+uFelanwt7XuCylOjQtdK448EtvQl2kJROYVHoKaNNt7GKnq4l2D17Q
22jHrgtA7Qikec4TdXJkYnsxQPA3Nlt9s8l6Vqovyt6HvYpD4Lt/xByUCtKXl2OiKx1wVzKOEK4Y
68b0mXHOPaukRigUvFCjLi5+q4L7uKiNOZjyXUDEQjEbRHZ7QAjjlBoGvRjzJ0WFOvYx+QexOaoZ
TNdNCjrsOAo0YSucRgiu1IBHMzmNwVLmQO9jCg06ZJo/EYKd4WCnpkgVpc0MV11SahXi4eRGwfq8
O03sVXX71MYuhIgI2Dm8CK3bJ70L3umAMs3LAfn4ZuTxU3yntWpfnbfDJA/2OZZ3dkBQ4rfaLBu+
10QzOlFJe5YITMToPgiGIj4JSFC7jBOvLO3RuxxX+xXkaZyazLplpMBbgMRmrJcsnWGHmWfX6POk
xC02YBMPtXvPhDkNnPV//QYu7PaqBBu70c3FgKhPD9Cy6vHRyONWq81gIKXLLm3b84tLXE/HSWlE
3ICxq7DOBwcHJjsQbEKIEVFLr3YTVJH0/qLZQbYbFap2uytOiAn6tZQLngitT3BtmXokW15ha1WR
VW+2b9KT+Ycjf5tOw3vEVJvyFc53MipM4qY5Fn/VMjzQvw7hPVstJQYJn4+4RGmyNJe0OgwIFuSu
X3F7zBMJPOixPOP0ZuIznSYk1Rd+daDKGW2BNgVyjCJaNEmw9NWgxOwX1ocv2B+WA9SL/fI+Nkd9
gcwImAoTVu9j4yowI08LQD8Z9VTZzT5cMr5Tg301WT3eJ4S518Y+W56OK1ZV/U0Wr5m7+5pdIuul
7csv+oxFZT3lKlhggXKsKWSpm53e3GWDFp8l/cr7FPPTZmbIBdFofYPdBaN5vNHeGSkfBS4CS4nj
n48wZNb2/fP8tfsqUU1JRr3fSRJNUq2dAzuWr4s0FdhbNuHqQSe3Is2xzH4XOv5EZIeEtlbe6GLH
BTNSXrw+4VlYZt9dkvuWGXx9teYS6UTRfl4N0dsHJRnXJNxx080EbxKTGJteK64CbdQWfsbIvImr
asdxAYKmbsgNh3yijAUY2N1cF0ivZaQ4KUWHF/gu2NPXuXWc7bSoR9Yl7Do04QbrdYtiqPa1skTV
QIq0/VOU6mCqwdL5wsdCqUbRrztwr9yly3cSqQN7/1ECjiqtIIl5jZ00Tx20MWeFwG4TTuLcCO8u
Bgvfq9qmbMWNVD1I30nbUGMM7NT+UCLftFqDBveF5UM3NUCuWNpzqjwTt4vMsYWdazbHwPnKeV1D
T1We71QzzorENBdTqicMzTH+j/MYdl54GX8XpZBPJ4pN7FAv2bQEU/eC74saRlEvXlWs53Z87DXK
Rp+PRSsQ8Bm10CURNsK94maldTnrYqBwBwk9Hk88ivBRC6Ku0C5rBc4crF1qcS0AQzOoH2XQ8KFF
4eKEty6hVfdvbjlGr4GRaPcoHvZJA3NvCTjTwygE2g1s+nlRnj36DWjE7tCPlKNVR36xCxIkd9IA
KUB/6MrpFJFRRpdD94VaxlOablJ2y4Hbg5RC+ntOI47+vFXMGJHTOx5UlOhFKWe8y3cCuSjHttOi
K4tojGTroyTwePP/9JBPusPw7RMs0jN2xmGEhLHiUUQpwDDEpZ6tLmQwP/pUkyGLt8mzOPDsqZsB
e1mDdfyHCQoGKp6kxF5/UDk6ewX2UzKJ5+Jcp7VC9lMojWSI8wz2J9nRusGu2wPQdSuKvvrUhzu5
dVtFv2fNLi4XDwT8gbPMCvsSk/wHAnpW2xPxodYsGy0cylfYKVST19mp1k47cPeiu4U9Zk9vnTle
iPgvbOeDH3HTRfRTUcTfCztiQEketgFRgR0hao+rRWOtp8+MoSJBfw20MDfMn+zlLhDkrxpC9Nel
jEQMJ9i7daEcVWTSNl3wo3UzgPrgTgwDc/rxAXv+7t7WDJlQF8l7jpAtkbiIuENeIwRBI5auxKqp
ustPfv2J6g3KFJAFin4j/y0FbAdbDetonfB3+fLzd40vBd7yXkMUQ6j0kmwnVymJhSg8E4CXyRly
cVMYCYx2IZbRZDoy2eV6d+FJXIGChIAXomuNYuD+smpqBRMnMaqAc9fQfSOtKEg6zfA6F49wRlZK
psp/KTjSKIsOZsZ1//dVSOTvv5/ynGTqJmlx8dq0+CGex4lG8f9nDknk+vBINfIyvUvNy+tyrDaC
kZVCSiVFIt74lCrhvz3ySZntIHGRMgYBVu0WbV/dMHLuPMbva/2sWw2liCpCKfLyTiB80ylrenSL
crCzynGd8xCNwoGQI7YYTTGREdouTwSag0dExkIjRFCtPh6o7Q/6uBhP3YQFzHL6oe1iClXDd5Ko
7LMNyVl8cci21KDC+DXefHR92N9FvTZ054AIq46uZ0dSnmH1RRJLMMisrTIfjOdGXDsFgvzsljdH
5ONiDYnf8yPGZwGEQf5hrttFfzbqN8DuCA16kSti2pC9zkmECBaw/lghjLe+WjI5JicdS6kwXnr3
KZPNegJP9yJ/ZCDolEhyy1z7c5zf9LhHTLeh6zllbTCZmNuJ1btgjxPzWZNamuubBdZNJ/wVUzUM
tSpTsrrki0j/XSOFZt4zRv/z0CVPIqjgYICFDW+rvwTP+IiCdA1v3ryrOwI0nfQAKzsDlkU5xyBm
A8DCiSl8Zk4tnqwfo2lZZI4Bw55DnjQqgFWcgFXY/oUqrD+/HQIEmmAZ8Ia3Uq1XwOyef/4mpc91
bltlzMeZsJ6/xhtR4uaZRa7CpGlQhUBobDG9YrifipjtfLDDx+ucWu5nmLFh35spyqrCfS+EzIql
+DFE575LXzGmkOthIUEa3EUmTWeTRGjjOHJpJLPMfZqutdEgWnZL/0nDQhdCL6BV2wF8olWCb3pY
IB4+CWH0c3JGlvWoW3vF/slZVkv4A84AtXdY8P3Udt/wjhvy56jXs0KrXmL0Tebx4e4C6RWAIsy3
0lPONqqdz/JMI7WY/8bveGrFyb5V/jjNQvO5JfUze+RxlVzm7EA/WrBzdvyJ+CEBXA/tojS7TODg
5lRqqOSsMwSfq1C+F6TP821pXatDn3sjaCyCCXqgqY4cP0lGtVmKp73dN57/VaPpVsuMg3Of10vx
iZt+4bw2w3qriN2ujthvM3H9gMqtODVy6G8+KyuIFJyYmdA+sJxmVp5JEwla+BBpRfcM1Gv6FNnm
6Asc+0dVMlU04YfAb6nryzeMtLsQoRXa7k641wNXZrRMog4GdtKuXcsnmndW3Q/jml3z4ldAivF+
bzu15xYo7LTKbafGqExNEyHzH9VFve4+TRuHAbyFQWDs0ZgCU6HMrcJdFFqTCDl8NTdHNoA0jqHW
VzA3nyu1QSpiE+CW/6kYGS1bgnfoGmqFAwUAC5oqamHN3MO/pQneehr4JhDngBlQuBuzWQhL2TLK
64nRpUAdM1L0Md0t3vJU7j5rc0bnvOL7vNwkTBA9soZXHj2upI4PWCld6ZKofgPx4El48KQ/uGAl
VVOgPj3USgoviYiX/EhmnTQiEVLF0CB9uBR3n00cM6gbbGtTnn1R+PL5ki4Mkm5pgRcX8sDViP+I
mrYgVRAP84AzC6moE2FHxSSO3tLZ0Vn1LKGl4K7iVPhm0lmICfq+9oE/EqdWXBcPqF3f/jo5wpFc
AvEeoVLjj8XnTybNks1m1M2CWNuWT9d8DvI/dDBVL6cmeFOIP/fQQc6vxZQ24BW5NglUan+C3lbj
WuqJNAfVUXmBDfUmg+zQUWYGmfKFhGoLK59jgpkw+cl0Cv3B+DAXcWLy57Ta5wE4xpAyU+iZf0Ru
uxQWJdbDhydUFe7oOvIDkb1rciBT3LHq2Ssr/Hk/2EtjYHbxxSATah9Md+myFpR4TcGE6RhmPdGQ
fpLiwwtHaYlnSdOfq2Tfno7nY8dTKVX+OMqvGOnSHPEw7b7UWl0ER7mGuistK2PGyCRCn4UY1BbL
EnaVh7G8MVSCqMYCTcZWa1RVsU0nnfi3Vwste1etj6INCARqcvGsCTi2Sth9+bdTRx3cwA0tvO2g
ZRtbwJ3YLx+8FgQ/TwwFdnFBLFq3wxFnZYSyWdIJQJaCBHFvaWwxTNcE6+vCzLKidYMENejx7ffW
i/R6nuhAk4rn2CJHE/JGFsvCCSNBQbxegSYhFEmZKo8VbA3GXcYOI4AdDS/ZU1Zfl8n/Bo2wrSS7
XtsUd07XlY96YV/9aJuFd0+ME3wOYknD735kzR/fK8LEOOlRxxC+xIdSfZLXS+8ZxtOVSS4c/Uyh
AwivL0BOqxddJxXyx/UG4bOOtlwkPPz7XEdhwqEpioCtAyzn7u7WdcvppPluiU2dpQvY/WWUrbEh
T/fFKAJKsSDcp7lPHD8dDK8Qw0jPf7XUQWEs4ggxenhJj4yq7kJxRTusi72qsVzVYcZ6Jd9ZhBnq
HUI/3o/+3XYOA8ZMHGdot3Exoe6hO+Nq+3K1xyOvud0PmwyggtmlbREQTErU/eAgPWZ+0v543djY
E8KQ+HbX5j5OqnRW1VuW2VzB+NGaZ1sI+8iWLWnm26ynZbSSaeQd/jKVbgS+EdjB0oSo9hgn+k9l
qCKxtKxcZQR7j6/b+mMrYxk6kDdPQVk+PHIB1j91BpjaFTp5dqp8mmN/Cd/nlIgrD7BPn5vIAjMm
E/OaW7GXqoqmRT5nNb3q7fklX5mxkvKJ+nRsBHfQTlG2zuyrJZnaJfiTpaGPolxNJNK78CV+hFvE
fXvc+05I2+0NanyGmz9QB68D7FRFE3IYxgZ7stayGQaRe5K00fUKpzfnJVQbZ272nD65SOWFh+8m
e0rWlB15g5ccNh/Au5b1rn7evrKvoWaKd2QcjUNgaDuC5mXIpRSZGZ2Q8KDnvTRHzWAwWj0i9Grv
0mw6niIJRN8IUo3zBY6xh3H2nOROMZOgEMBZkB4PAumTQD4rYIRIk8vflBKF3bKFQhO5FQMMuiTz
/rVaqQN5yRTbUqwjLrb/eMjr0RWFJovlV1wjeUVALCtZ/rIH7OshrGA4spL1liycEVfnpLgMJYH5
wflqgt42hi8REi5ZMpid2PxN5KnllSRc+xpFlzQMXtpaymc2R6S+wQ+TZ20aCyhGbjBf/UZL56gX
SnrVZP1X6e+iVMTT2g7BEko3zRYLienDYKJ+D3tIvlZYlaj3CE6RoGulceu8nx3H4EO3cOg/+zfQ
0DWpmnhcgjuQMTn3g5rUpybx+Bbt7YGdfr33lBhkg90s9qzkvCnPQ7n0cpaDDUciLGUWU71QF1TB
/025mteiTufJCcvCGLreJg0PjDwIzmeWd0iWfhs2FMWZiG/0JYxc73CJKnd+F/SFYSY9xIBRRePG
j5wIoSeMsSsMKhGbWoSo6dRGVWzoE2BDYkf5vjSWmvUy1LnaOG6AGWIVude8klf/9z6FEMYrCt2x
zNlkoAWGofE5I/GjoR+KDCF+L3C9llTtf0AaXeBw7bf/31ojFzix1VWeOk7P8sfG/N2Ty6ospoAN
yz0dnrRDxLVqI2CNVXZ4riKakQ5LpNUy7Uwjht1QUvxp3hqjkeOrNKm+XS9GBU17uMB/nMPxH+et
Fd87sH45QE1BH1/Hkp5kCgsMacLrZ7APJ7ehRjq+DmfOWZf+U7sF8YEBsnCTgC3ss2GPf6uesT8I
Bk5ky0+BlYyIpv4UZcpvcjLugf1SmofO21VEk9HiXtUS/HXiAaJyo2FzDblxyxWNAPzQJtESuJqf
IoJSnasGUpZMqVNrSiBOG7hhBN/F7X5UGK4PfjcP1n31ztDeVLdAJiMAoVvca1qaqkbL1GBvOSLk
m4eAxHYIR3a7T7RZDOxO72Uu05Tq9Odgjw9qiE8k0q+bzp2+Q8AuRgqMm6xMIQzAycS4xJDWqtaB
gMn5oPpVmtYSK1mi8ygMSJoQGONGT5VRUTg7h3dQR3XMLgU4kkExKrElE1nvXdIfMr9yHAe8kqDj
oix3fxmF5jdR8sLRFtbrt0PjGQiSO2ZjvmFCAE3CGXWVdwlnEedUoGTXM/yS/kZ9rbg2dRCfvjsW
Rlfm5kEUjcFlTTcJh3eOKLd/37eH0IvgnfZftZLsvJbYcMFsyqW3n+Atnwa/lzUsMCxruJ8edtml
VpqHhlfUGGDE/yn4n+OOHhQ+8syd/hUSWGWeAExO3e9vIOq7X8FrNI44igOCSTXMrJDwsTRKz3Zn
eX+dlbdOYqF4LoS+kgR41cBICDC383XwhlVrboHmM7JEIty/Xsu6FKGWPcwEiT1Oy/vR2m13qP6z
Q8fZQJrKoBkw+3heOl9usIqnE8UNnN4z71JOS1G04RyngM/ZNAHk+fp3xBjYLewH0JTu2eF4iYxU
lY12NtfGRyM0JY837b7m7fmJ2ppDsxZIbrKq3asF+l6KBbEwvQDCHhlz814v4sIY2L96gVEADhRj
/fc0mgeGKe2rNZM+qVqvqEygUEijjthvDRznnUHvSBu6klps4or2WHYVoFeS70DNYG13uRbY6piI
wzbEi76Fu6hRay7NPBpBUVXFGU96QZAjz5nvCoZm5hmcCyUcKimlFI1SvKuIV09egXhef9u6lwjP
GRfFsrHZ7CJbVkpxFKdcJfy89YhuUW8gHR3akGwOK1HX80YXVNlUAL3CQofyY8cTt2rA123BzIvb
Drji5YU6y6WP6zCgB2KjSFF9Yx50PDaIzSlADLJ1fdLVP9f65qr0ZBhlA3/Iza0fqQ3brln4KZng
LhSo5zCtmAqNOiB/QV6Z6brg2r7ZKtWkLkBG5SvRPLyWpXLKVobxkmqMGPzuvihze6bxaLPWqpvC
NoUKDnKZybtUliEIEKPl1Rg5DzlNos9vjM+Dhc5fetBsNnDB496AAQec+njIT7ai/82H0PNH2nEV
qm10a0wYHPplVYw1k27L6HAOtr6RmoLesUR1QOYDa3C0IM0aZDx0yx6cmo3nezvbKBkvc8NvgG5s
6iGodHVYHlettWwaOoS0x++iEGi91Hs/BzUp7waXv5hWYPKqaHEPyqfw/oW7qtQdNTAkCYKUCGBK
fL+D1aErvbkcE64DcT/cXitbLWXKtmIhnmSJ2+bkPHFpGnUI5DSLcE+OjNE3E2CoYQa3IXcWZfcs
LlTsQCWlyIgtJwcU+omODWLOt1IeMsPwlr2m8Sk/aI03Q+qt0KrJIH1NL9gJG92BKANdpPvt1D8p
q3cq5sFFniCG/aV+P65CL7BFH5zciGdgaKKdDK+IRR/JSGWZZAHCKWqmw6QiksVmO0CQZ0ilO7mF
JM0GqfW+k759P3rtcBT/wUii1VWIWVoU3L/5DrRXtPoPjD7eLu/k/ipxdeG8EsgibdCbmCvnLH0c
o2GIUAscDLRJURCA2UbSD+xSsMWDQwKUi0vasTSt1EKGXIk1OMIiup4LPFLdhMIfLhHZOqOPqhUA
e0nkzGf26zHUNVcga9Qg3EEwvEx+ZZskQhQEN19pZ8x5jc8AmBWygDQ3N1a7WwiqBjKeFGTK/Exo
Kg9aj5aA97ze29ykE2VU0ycnn6eXZDRrhJr+38VT4r/ZPRnvxWJoYU8nZzhU5DSF0TCi7/1ajx4n
qGGHGDWeo8R07zLsK5t3Dl6GQWuTB06TUFW6fz90lYPql8QjQ1T/TQRielvvpx8oztyyAuj7qUNq
nwLBdGQKz4jrNoOROfWDQiWfTV2rAGxXj8TQBYgF0hrJQt9uqkboJzl8UAHQ8Maj6tq5MmGk1XVE
LxXfCXmbJLBVmdU0pO8R6XPTo5D1MwVrkCcY5XlwY1jn4+k/mU0JNdzclA5cBjSRJ0ObwrkrQBc3
qU5sqXfldx24g8W6xp17BAjWTa/MN/oOQz0XrGaSeyLKTa9gmDuuYPbRWxSQ2Od5uJnXQ2M50xdi
RDYAzNF6hATaYGHOdbbYjAa9Okohme0OO6RVU0nsNwDUrPc9qRfY7iRfrU06BNaTBW5reONQuy0l
AYdNZSPJA/A9By+77iTA3hj8X0Bf1UgU4zMRiZoJdmGZUVWxpwLz44u/MkhR/0DlZByjBGQSIF2y
E3yRPSp0LxsNShoqpOoIs8FfnWzjmD5aaJfpNVMQR7yFKwp2BQAbSGTBFXQyPLJWKnsIa1OCddz6
UsWpo7QKKAZ8mARCR8jWdIQyfEbDlRmhKsnvALVMU5GgCp7qVsgc+3xeM4NQj37mMEb3GOX6YMBM
PB5P/naf1sMdlU/KQPOPbC0I6erQ6uz/5a3ZX4uRiBjsM6wadIM2mVjb7kacZj/ThmN1oaITUsL9
VymS2EimOCUEXKwbt8wQui4tqrn2Ao/QY50V3+rsYlroXg4WfgkpjKe39t7Eq16gdPMQVxo/sJ8E
4x4eomb5s7Gfr6KFKnXsM3Pzs4u0mw700oMeqYIlcUG+RfmCn924UfToeKX4QLLFnWYOoCpZw3gC
xnnc9L+Jr+asZX5Dhxyn/nS/h0qB26OQFOXosoQiHsKWdzXYVQ7AK7Df9sqG0SyBwBreQeXrx042
jHiR/EkiFqpkkbQtSa8Fq6rHs0dqu2J52Ndwb7digU6StWDcxhKq8uCCdj8akTCKRlJKUBxlgJaW
6MVSdORZFROekYzrxL1YbtAQdgu1NhlUXDOmExOxSny3tHd7FqQHqsopsp2sposqC8KAQrEfcw1T
1Ho6Q161TKpqcEER/OIElFi/Hd79LFxOEbNST+dEDm3Vsa6Q/WOHdxCS4CGi/Qyc9GRsY58qsGht
KTjn4u+w29MLzNn7GUZHI+XtC9xJQ7tDpMRo0b5/EUsIjHn1mIZxe5hohFOujiee88GrQpqMZdcJ
Z+klla3FfyK4QHva4a29zdQ2WIM9IQhQAslZ3IAhwFT8NJlqe9/bKF2XoBek+Ikf2tRgxwiJr7LA
qeBnABWuUz0CORk0OkRGAHVfjMNChjNYEn8Lk5k4GwgaB+KQah1EKLWd3VW0mrN2EQtRb6JQYb+o
r9Y3NQ6WnnIA3KY0ukPMG4QOWICVfhacobQ5B1UQpZ0fivV5GY/WcyH8l9Mn+Y60F4GnBiG1AH4S
P1XY1WJJ/47j8aLKJ0UP6Fiqq0cwNfdXa/8oUcWcTOBKkV4RiSVCc5ntSanoUK4Z99IHaxU5pUWU
wZWktp93jXviluoOEEHG0JSHNC+N7yC/kxS6B4Hlpsbd9BBQd/sO/cMpXb5IQVYV9e4S/xEwdqPm
Tlqz0Sf0GUQ//YyR8rVDx8sbzW3GXUuE9yYcxiOQaiP3mdSEopyYHSeoKyDwkkJiGb6kFDywOdJz
usEX1g9frhHQruoz7TVdYuyKAsR3H7SybvNT40ocNnOf3jAIzaf/ue8VhwE9PYiPX0kVyMAYj6qx
LjxrjPsZK7c7PWmigpWD5v6hfBv0+tb40Q0ijY+iu7bPWE167hCfhpCLTll2R15WhzQGmP/qY5FL
FpaEXoeTkxWtbIHMyn90heHonMjcDPysl96Kd0KC5mjuTpWZ2aZjsMJfURnthRP+1qM5KdJKuyeR
Yvlpnn3iyXcJ1aYPS3vEyCny4TndyMnqHB3WHgbndh8ZwvWXrTplcsBL5599metwqwRTUUuC+vn+
JKKw0hEHcADgXEDSkCXr29oIRaTurtpoa3AgJqyBciQ6j/a74JMy7OAMq/O8U9rHrHfLThI327eD
LCq3OeeuDFlloyrGrTTmfhZfORdpBMMlEJoqqG47NqdZ1hq/8HqAOAL+QdNYmAC+hdLwBQ2uIvUk
cdpR8b/z8soY1e29z9ir/bxx7+jYV2+XqyeOQw3V2YEM28G+P5yS2F0I4Or1X4xCsQsPGsGQYsj+
15fiy7T8qym/PvAAXffVxaW8/6aP/CoZvetJpBrAKiRMg2cyuFQeJDmFWA7Yf+p1eyG0pymxypxJ
fFA8qSMJU/rjhicw9jPZswF1bXO3V959r5R87I6t+VpK3NU0DnYhtBeRotaTAw8c329vtIOnEvMj
gURwr6Hq7Qfat4Gw5Jy+oOC62o/rIaYbA5f5gQrTGvs6ciniNOPZL7+Ae+6u0GUL3OIQrudxv44g
er5cCHcA3e+A316oMboFwBT43IWwvJarSc1Cjha5jXqxfiMkG+DIbe2c/qJvUl0ZiuqvP88Jrn+S
unr6Zt7IbK+k4yIRtecJl4JQpDqW5Y2BhFYmbOtiCKg8Of2kNunEq1yA47Af9OY984q2WE2Sl03G
2M3ueLRWSfnr44qWRzfgFMEUs+Ldkl2usCFCJspAgS5qBmvDsMfk5GNOoafTAIUvLeSLvL1LLStv
vdECyZRHNgL0Otr9OzYeDKhTEyIynL7lsIWnu1044PLJ6le+dxCIYAwJEet0rmbsuM5w7jt0eQ/J
MLwkZY8CC5B3hu+0sHyoME7BkP97tk8+cb/NyGIGgthUea36Em1ywuNKJRCQUplJKKD34dPjM8A/
sam9kOvyaPVngUytJxtTH3DNT09VCcADlz+VXsdU5jXh24OtW6hzOce5ob9ohpbMVX8b83xGXKxg
sxZQIYvCQd16UHHYX9Ft4IdVjXj1NxB9T+VqlTLqLvdpkktrqmOK1T5azDy4xmCTSi2d5Px6yRYC
LdtnpkVZOe5a/yyYSRj0GyXPOJNNb/BBgNckTtQ3urXZ94HzufnyPD5esDiTYKRMJ5oI7kGgPxmf
G1yclLlOFMFGo06YSULqgSqydjcimamdT3LF8dmimIIM4H6nKXhzYvlPkyYCxesxqMmU0M34IOQZ
Fcc3tf9QvIwUEUs2KJpuJ8jrfxvwfKlnYq85Uiyoxi+bv/kiSVpx50porUzSzlmEKIlzCZ12RwCP
i26kwG/RDRRnqtf5eEwPalynbsxgdsIbSAkaoS+MVlaEWG2q7QAMQGVfR4/A3BRLA6sYxZgdDnGw
yzMIHmVUyIhp9QDCnhr3VKjEf4WlPQeBNmbHaeIkbKnq2VX5sDR9fDFZCJl0NFV6O17KcI8mc8k0
CTCj4R7Z4BtufwADTGBjPQ1LcKYZWtKYxBusU4BYH+EJeaZhwgkml7UrXvFNWbkJkygAp8CRe7ME
zdaVy5mmHtCkRKrlkgtHSmpYYNVZgCTyR0hgYDjd/W5hQBpD4MSyh3cqJs1CYPGOBrhTMz2eduOH
h8FnUrBp3nn1tXdfmpDnWS6BjqKP6QhPR0Km3oMn4RxBp7YxB0q/iytQGX7BHjNztYgSK1vqenRs
pFoieZOIXHdL89G8JYAmpjE2KLy/6BhvK6GfBpOPZuZMAd1+F6VhutzNgMyL65Fd6nEDWTn0t5il
PkXsMtaU+m1URF/ml/MDiBWk3JFYsvoVwToFCaVhtVOFa2ayLopc4mX/sXF61gc9S28A3gD5hSfF
nYr+a9T6Q/jupzp1LjLnL4fEQvAPp3iBcGYsov/mq0tm9xYXm99/YFbV9D8NZ3UmRa2p/ZZPbUHa
0CTg4rSc8RRTeXieYDAlMxp1SvDupvRAjEp0nCRHqKr0VvpMfDfNY8lyqytlUFjd3/6qFJBg5TOo
3CYh4QUDIPLVm4fKy62sOpw0c3AZ65K+Ukvae1hLJElEU0ZbGBOlXD9M1/sNqkhEOSC58r7yGU7X
Zt2M8bShToitMwGRziMweEQg1tttYANgVpDqfTYpHcdL16+Io817PaKdyrYFEeUG2u/c1ivaA0fD
Lqj2RwkbO91Bg03WddIkIeSHfKGUIJ6BE5JdZgRZFTRdSsDOwgOjUw8q89IhWtS2PtLrADFPxMpn
LKpv4gr0YPE9ewvPCPaAO8XMmGGpiq/k/xRlyRdWt94jsyWtIYN2A8z1J3KnIZHPkFs2xUBc6ZN8
L6Ov6RkSA9WJ/3QXASCbkJJi4xhTbcAznk6Yo6zyKoCWBh3Ay/E15956IEJPs9ulVyyyRM4RWgRV
SxjkMWhH95v3fQzSBVJnAPoH3ra5+I/ilaEi0kDP/s5fiCOXumyon0Z4I5wKLD7DmzlWbsEs0IS5
XKmYy9zvKWjomSUFOvs94NdBI+pU0zaSwhvCYPTZtEZyK39eMGdofmfuFMJmnoeHwRgnFm+LdxW9
Y2c3iB2FsVaBRfcTHzwDJExfVrVr1xEt6XFIpVjE65szX6EBAtN3c8uLqkYDy4hKMCrb1N1ujsO4
Mz44Jg20NkzHo2MGUAZjIRRRe6T3V2rFCdGIW8FejzpZdAHzkOUiMaZQMh35C0+YLnhrIC/2CGQ8
G5gXwbhi/KxuODch98EJbUHJcFKvGIZYhgpz+7iaxUMiMuwZvZdH/9i/2GX0Cabz7flHNM3+pny3
ssP5Prr1uKsQ2xIVIH69Pirkk9WJPgvPS0WzEOUdw3elwyiC0GcFfoZ5NacdiFBi/egSBDZa6p08
0h3uRvYvaeRM/iV+p8S57ui7tLwyF8+OI5unJWc1JQAv6bk7MND/44sIT6nDYdtC8fpnnm2Llc7R
Dg1ia+W1LRGioyLYx+YMjrNE3vUHb6D0jIIFVvoycJo/jY4eSWZbBvgQUUmrqyR+QHdaVA/WqVBN
jPN6mcKbmSm+7spU2+GVYeutq+aiCrIbhdg8iNyHEEzKlj+8pDbp+IZT38whdYRTcz3Sfb5+F6tC
Whz0pxuXlsfdB36Lc7ZF97318Xx7H2mp6CkzI8H6PL6thIxaai28YtmpxOXDm12hp/dk3koeBFOU
SgXnDpxwOMnIRI353/u2WmOJN+pxmVvEELtqrte2AD+6fDkqkzs3T0HnoO/YtkGNfwVgS0UjDfMs
9wKRviFQIHuAGyEiLdsHWc7JtLJmASoLaHVDxYjq9YR48JZPCFqIPG78C9BXYtwRGu5+MM8a+DgL
4FChDfT/6b2vc3IHELkKnN/UYenywQ8b8e/EwzSWnkCrBJCN3C7enrIHNW+er6eL3N/90scA3RaA
F2j9u2SX2dfp2Tf4nrZGEIlsXzASVqK7nh0+F1a/vYkE47f6s7gYVXp8/zEsjheJ+7DuJLsdw1Fq
BiL9CoDdQAJeZzSwxvCeSBBGvprLo9ZzSNJGKpq+vuIkfMCFSVvMcS67ELtNah5pPsQ9R51rW69T
UXeICjFFXB4LvXMA4ZKOesOHp4Sz18Hezp74/uzh2IEFgGGVnvMva7jQ1/EHMfTELmScSVPxrSZL
JzGxG+WmE4QfgXvft8BAkO4KnhiQjjoqWXA44X2LyHpDO/7P5G/8osAwdUdjU9WHVVUv7/fLoCxy
IQavg0R59nou19z+vg3mHA6mXadn6ChqX3EjXyXhyQHOC5AV0G3trvpjqxkWWFYwZ+XGw+7VBVh/
1k/ah0u96u/q356NyOz/WyPvp1xGLe0zHxhH1WAInR/nRJteYFqOK3E6GfHcMBF9NIz9nneoXSIG
8WacwJgGa0yiGERrjldJ+OQ2yID4isTXe9K7KF+JTLj9+XDEAUSnjnzya6wjJYzk4d60yQqyyi5x
cZid6usMhk6F4BV3MFM1ZbVJUL+n1P0rZRGPCR8PUhrgDiYXOkcMPsuhU8vSmjHwhmaO+Q4CKY6O
R75srsYF7C3mrBUM/R+LRhuY9xl6laYn01PcFUtGe+7tIlY5bZ7WUtArnHvhpoPFPJm4zhOErd1a
4FgHuEcLazVBmUjB/wpFfDAOj5U5RgaK2DAqJPjn/yqzZFWcRgqPEeGJ5OEinbfde8CY+ukO3Rid
N3aio+IY/nqZueeuXHBeW+3t0dAeqpK+RPOrJo/WbGXQyL0jgbeWJMseZTCj02SgGYkGseesgJ6H
NTiwpNoNopMY2Bf1ZorhcYHeHirfB2yxjG1c/xW2vSE0r3w9OZyYUEV15P5KnISRzCYi8nv+gmeQ
RwNya5a+S4vNIPWlleeBIst01f8q/eNUDsj76SPfILQ/PcpEVrwqF1WeaNwGMlONZpHS/9ZVd0mh
4+cGNQ1n2BpE6HaakbQBn2dJUYb5NInCSOMieb3DTJVPFd82a30RPiN9eQrpAFHkgWzK+YqXKUel
3H2Kl8KsgeGTYtl5Aw+YrMuC6Lu0/AUrcN/1JhUbPqwJlhiEels/vZ5udBTnb7YDeKygHZR6Gezp
kyELx9yPy0ahR2TFwN/sOKvNut7GbAbCVDUM0qz7dYgU5CYsOYtGkLmyyZoU72ol+QHyCureFYu+
M8lT9DwyGsxart0os1Nql2jwXaNg7nkhryXG5wvgA6tik23BQLXWlsL4hVU6nP3AaAvbAICvRtY6
ImY40Z5fQmHfYWoOwMx06AVQDYAHgAr2HS6hGEUmHh7c78W1kXL+HSKnm/LbrTqdk6ZsoyVIYPlt
+eEbSG1GhTvdstuHfWaYwbhrlM9uMHR7LyeG5C0DMufB5e9fAP63LYOLqhy07akPeDcA5ygfeVam
wHTfE10YX8AiVgi0fGdisrGr4eQcR0L8yV13/j9Uf+U3NU8TiZ3CLQ1Bc/zNQgcsCRvdctAr8kLO
agCrWWqc4WbbzTidwC3zNB7OsOWqIbCPnSmKMUrklYZbnvBvS85lYkCm8RWT9HQw88I21xjNgBLk
KnotJ6G8UCyyXkWGuiB5RG4NiIhKG3AEgLC10xzDGOFn0SzQ2nQdvuNGgRES9DRxY1I4Q9k2+0V7
nDS78x2OITq3gda+oQasYsBXYGJZNrqUnKWmoWtMNeIqTNg9IcyErC+3TEKD7EpK+zeyNk/6BjKx
zhNOU/FviVgBd7SlhFLuiaPwaG2lrqHJY+VPRPgQGhRzS0rtMKoqLEkxJx/3ej2N1pinDu90tOMT
5tHHPhI1x0V9UyrpSULYqmES8TTfrkBssJTXTyo7FA7L35SPuRW0FRVm1hBg4/IhT/vfZ2hwtYkr
VwZHF6cNGgKFK4tWqL4vir88vwp+WQDOEiZBXbyb6/9yM5Gm8H7CHRgi2ymKy6Ij45u5/9pYIpkf
CGWThcCApM02LdYvUPP6FlgjzwZtvExYKnfbgKY+rMzkIpYZcaZNd2TgJXw6PXkdRdrbhGPPLbjR
ho/INjySOHFgS86ZuDxCV2R6ZYpulbMGl3XXZFz4HBbR2tMWfs5tl5PoixkhLaHZ7FIv+fRZI1lp
qdjBcNO8vdUR/AX+dRsZgdV3nmnCCnp7U0HzSOTfnjgJaQn94hm16ighfr38czf5Xp0V0/Q602NI
gZYPQ/hhd4fjuzcHzG+9dG1kfLfDLyyHjix1VR6jnyaUXBKwBkOZCpGTPTPatAGU5W0cHiN0V7nJ
B1QNn9/SzSVN+TSZ/vB8CXknQCUYonnDj3Xw491/bIFXVrg0xIjZPCbpJufQwtSi2DilRIYjYlsA
W8/+u6J+rnoiA2wsRl7sgMhuuWgpgWm+n90XoZ6c635sbMLJ+zcZPUMCGOoO7rycu/2fh2EUMj0W
MqpeIDCvUHzI/xRpNpecIF/sVqfYEVvomkgKscSVTLtN/23aEl3NE9LZBwcrj69GxSNIeCSyCjNC
vbMFjFsv7IJrngGPflATjqoF27YO5X3JuMo3HNgApningcpu3245I0PxnxIEvxfc1NA25AvbREcT
MPr00Lb3iKkP4MGHMzJcFZ1znz5BB7GCs4yokYOByKcTOAQ014Ty9ntaTPXZ3hbI4Qv4FTVJnrZo
fdCBBb3DBLByE27wcrPLnWEX2PbKtZoWfX6S+bKNmBd6HafxGSqK0mLpHgS8xYTPigekFHUO9nAO
jJ6JmjvcCydCns2GhQLqzyI6lKAzNG5ModC2UTWsG/XDUjGetFjo7XuQih7CVyHQCw8uLpzCXtNO
03lDNmiJU2Gu2t4zpudjc6SRkHaaH251k5NbIRmnlPM1pAtOw6Rn2hd7q53ab4UTQfq2JBM6k1eb
y+yt+83QEwmB3NreiClTVwmbp90CXcNwL20TXQqftB3SWQDhTc0tC7lEFzlL1K1OYZ6Z+Z7EyOg6
AiwLg8m71CSBIiZ/jAv/n2EvPAg3nQuy4DbZg3gy3np6M2xg8LItm2VJVKc0a4ibnBC9HG4P1LhN
Dw9JFkGr1t8XoeCTJVpERGT7Vwi/J+yG2kQHnBJy8a47kVsiHRbT4lsn535f4Gdc4J6rl0WUvlXm
XIWtF2mxt41Jlnjp0TylttoN34dKE6eAaPyFirzTHE/NZTpyOF/GIPR7ynLpUaf0Ea3GJyJw+WpZ
NWN/xCBvEr1+vGNa7CCOEd2LUwFhpEvvKB1qrhc6JmjbgU/4DjDeeunc5intSb7pJiKFDftM7ApR
l59pLcIHbfrSJM86i6oEr80lAtIjJtRiwiN7Ad5XhU2p74TFu2TtnZ72ofVFjFFhi/QyA90Z0Awy
HzWG6qRZo3Nx/oo6IYFlh5FCaK+tCfNlphnXWEDpBUoVVv0+ayQ15aAfx86A3Csqizo6pbuYyj7d
T2OyKADbTVIEsqnZcslooSMHpgbXNmjL259oJB6xzTa4IhRwUsNyDEAaUretY5+1jousdMsKvjM/
vsGe2ih1r/GYoP7PgV2joDR3DOlcAT4dh/T/PyCX3h+sLC2xjTrbAMrEJfxEqyEcuuhAAr3AF2FR
iI/ZtneEo0+EU3Bqs2NYEnO61XNBpFuPqE3fOVZWZ2IhLe39cZUg8gN56UdE+mDH8sYVYpPlECZg
EopHrJ+SOVLllX0FbnK5WgFemroXfEIINaRn2NYB66/t/l7CRvBvIQgPg0KIhOcnwvmsboz/PUp1
o+ARo5ajNVkkYBYOTKJXjMUHR6T81+dyjxdzigPCMHW8WCGN/liplQd4tVp2F3Gx5lJK65r3SAiA
twRPQrxDJpByorTEfZjdxKzgdRZu2o71y4t6rJ4HhxNfOmg+RitFcwu3WoiAmuLE+6bJMCXatwrI
VmQfKCEPAkIwjjd+Ci2x0WqJ4JGYpO51hBuOjeaZx3lINW/zIlj70q8aFWuEhnjvYJnxJHCm10nb
HXUR/ohfTSuWSaLTg/SDXsRopp0QVZuBJASPMlFx93njcCrS04w+AjeipqWxZDSO1pw143TiUrq/
n0PP6kIq1sZ/bjp78FuxWCT7l+wzMKVQG51clNwFOuQMikIaOt3cH9TsrzIpDzxbpVsN5jHBfSCc
V8ufhtIoi1Ud5Y8p84LV0vppuxBC+glkViKBfP3NXwhr0OFWX4Q5TK41Bi06KhLfJUM0ctSovD/a
tTj2SBPvtNpLaTYpALRUG9Nvw5mZstjOKcSFA+uAD//n7/IiLLoJZpuFyZzI3U3/LEoigQlhkFSw
1tlb2DAe9RIa8DJq7Zm6Oe/j/nYFrMXRSJYyOOKz/kz1Hifj0GOmhsfnzks4dlFt/v9GHhQBAnfT
K5cyEc9SGrOh+KAVxQE39WCrQ0wuPp24lRWlf4JwbJ73W4gFXJbO4D/ZU8jA9U+uMbtHCA5aNEh4
teBUWjXUuSosogeTvWI+BopEoxYDrnJEo8+KmCzEZZr9FBVBdFccpIM9Te06mNcdwXAO8DNiYQh3
SGmK0VxXd0JSj6l+QucVJdzrvjxpOY/LrW32hOwoHs63CnnQnIW7NAjxb30rfKlOPZh6h7pUhNTb
/79Baa2CGtwblbEOW1dqj49Lrdi6Qi+fvdjl+7LjluBJJWcAgwWrlGiMPDQ5PfwBQnd/VueFiV7j
EmUykZaV+rnZoDCrU9Df/GnJqSaT4Zcwoz0gCziVRGeFJ69RQhWAwkd6/K//Mj5Kp1afiE3EegAY
ArjSBYAC/7G/XpIugZPLGGAURjqyMMzwf15vBKF7RBInJGfV8zx74DBswqQlA+7KbHGBjENqaGKE
gcxGMJ18yYPeyiWg+qEsdz4qD9IIVmahDpKGyfw8eIvF3krTJj6MxEkIKG+C8D4uq9XpHKjy4mRX
aSMNIj19HDvhN25W+E3qrpwd3ejpJm86rmGSyDHcQ37tirYmoSubw3uMPSMqgAglrxpST+i9ZkjV
z3e88KaaLQBTkqP5ICz+7Z7Ry3XNBYmHw0LLpnoS4QbdrM1cjDS3kuJDGs3yuaZ9aByBYqfxXwr7
aKStXbeiOWNMA7mvIrb+MHBEFWbTlJ+Os/o3JXqHjv4OUBrXxBU0H2EHIGNdsbkodcCK1ZwGLNge
WetjaDBgnlrBfdXhUO1DIb/Nu72Z/ejxnzm3RCyeRqtl7twWbxfT7rjMf3QLAHZCccrC3Wv6/PdG
I3FZbY45LnVLzISx50NE5wotUHQ7cDh/qmX151eQDiOo3Fxp0wBU2a1Mvv3Y9Cb+dls9Ld9vDX6x
tCOCItDVg4L5p5lL3jV00JqFnVsGa9ScYJ3s3CSQOh2u6KEIuAWEznAkIU0KbHSENipJwq5IZKFo
i4LimSQyOOsp6/so1bvL0m6yYfld0fPI4fDsxHsoD7Kp+W04vxS8I3UVJMhfi5Cp2yszQRQSPGTi
WAS/dHwBzCr7QD2X/ya5x/tNqm++QbWabAurFa5QKwsyGX61mg5sa5/8lpeoSLsV2Rv+ihsHT6U4
I8MBj2B0LWtvo2UZSOlrNvk5NUTqFPCHXBnlJKrLbOeqUGeyhuM6NvhoGwCzpc+/PJHcojwF0/U4
qWbx/rMKdM/Kl74XB4J7E4YjApdduje4r5RaMVAyV+JPndFSMvC9DT8UDFp9QBsyOefK/busPmP0
aHD9AZG5uVF/Sq1dq2KFLxHqYZS3z1GXiFX2DhfGONnfTfPOYc1REllL7dEDV1kO2T3twrJ+Gdpy
SZpVx6jtkGc4pzp49VnX3suRcIRZhx4p5s+xPNLgu3B+tp7qhHamUjF6GnAZMeUinvepXIc2wqnw
Sc95IOG7R6mblbY7TRThs0EwDSPynxtWYaeJCejYOlGZD5YpqoUrdW4/+TZe0lzAe4ZgqQyTEsRl
qYypb1XAK/CRpYH4Xhgn0SbQ3rXQSSf7oXjipiSC0IlKZS/6Y4xvvGNATIY10JaoyeDSqhOfQecv
hR0/b0YlpejFYIlRR1U9t9J4gvG38CHlDuEVqMyIK1tdJWVFykom1cIi1bomolX6pRhcaxAMT50s
KbdLji4Fwl91JrC8ROW+YVYH/54zi+CWGq8GGvYOd5B0gRnchFwiNMFzbmVaSeyGv2ST1LVaAWw0
xTLof+DsdlwYIeipDghzdjzpvLru6BkwR4B0u3YxBSFLdTCTVjk9LB7p9TOovTCBseqbbCXLpEwr
lu5c5xZIQiQ17ErMgbVwHVOhCo00hh3S6+UyuMH1H54S0/tX4apaH2s0muA+4Gk3LcPC2cQwqo54
pXKnW96m25uHIHRql4dcJXT8XdjFefS8LpceMlFwkI4D0UGzue7uzh+zeBBNiip7nLwQGJpH424C
u0xA5kKiOnQjHWERh7gTKrbp3xHNJf5AzHGh3r1eRcsWWc553BUlLWsaX9Jop49b+MZO3lobiKB4
llwettv6KOwvbqMT3IkVobklKbeSR9hRPcLeghda8gmt0R7N3Fxtwc09m2s/Cze3G3hKrftKzCOJ
PZLwYLD0Yf63qAc8dlwWayblqo8TNjGg5DGL6miSAr5eE2M83DS3NcBz2A/0pB4U1MhzGplYxmGT
gew2IusYQNCQ4OadGifOpIvngnWZKd0S7T02G75lyQVY/mt+zb14HtOk9M78N821r0V16G559sUD
9edHBLqzYGjSs06DWvZ/6Vjcf0lIcsQpZurlaPfiUNMS01m310JDH0HS6N+yFBODeYsTXMMMmc86
VZhN0yur/CS1S7rCj1HJFIg0c4HHT8OTGLv29CjrQUYzbU9zZ0GjTHxxzY/GgzKCTrTjNE7cVMs+
3cB9ybQcCiVlEPdd2+zzlWyEOr3i2GyGFS0tMkmJpsEmY9O4lecYdWmqVBcAAsEIqkjLSMbH8ePX
TwimBMy0PW6KHYPcG0CGSbSnpUN+8z9OkSBQjEeQxQbM1QOEkemx76+nsOZ8TOLmeNc7Hrkf15MR
IqqCXfsOhPFpefJE83ktBc8Ouc8e8QJCWYPL7tzDyuJJUW/d0Jjqy2Opfg8lCnxCJEj4NaiYwWUQ
n1u2xGMogCT+cWdy8R9wnqtL3DtdhctoR7KJ5vW9UdVj9mc0+JyyB1HSnMPSTLTwqd7dp+A4P551
IFQkAppRrlNNmxSpauSvleF5W8qxy4ZpSRQM7ZL8pWc3++3SZkh1VTTc/FBaa9ztpcULIQNGUOi4
Iu5L0lT1eVP8KMRhF2GE/hpzy3m9KtkgCiuf+4ZsehfepEnimOcNVKghZe7pp71eb75rxkjK1kdu
UAYEU8DC0MZSD1UVdlCArr5v/tvbKRC46AbJ0QVRwRFE9b4NBOduaYKYNqqL3AxjXpYh/xI4Bhty
ZsgB4DURZxf70L03C0kA9kyyZsGN1tasshPW8aGwMclEUSHNBzAwAvspY/OfOB6btCLWmNKahs/m
twEX20/Se3R4kBXUUqb/B18eKsA2+NWf5ETD9Z4gxu2IMeHdK6C81CDVQIBybSbLll4DTmqN2VxA
No/SP5WMs3CvoOESXEDzCvwZ6Xt4DX5em1paH/6QNoyAm1Wb8S+CkTjDVXqDEb7H4A0nwULdCVgJ
s9x4amXavlqSrVxyskUJ4ni5Ci+Ao2NAie07F+z9C9U6e1QjCZOVNGRb++wzICRWL9rGkhui55w+
4rndxtNq1F4c2pnxEUmCTUBd/ZhLoGQropTSAZbZeARwzAMczbkJQ/hs/muu8j03SfY8dVR+MOe7
5bLoLVrpBbzCkNPUDFWj2BlepvHQuQqse4F7o5GkT1+NTW+Amg9//kiA/jM5lfkxJxNzMJv4EKUP
8BHmJf1v6wfjERyn5IrWTVPn9auyCFJkdlNAagZjWdSzsmoaZVbphIwBsAJg0rFjXMLwV4Xw7Lac
+MDXLQZe5l7LVJPiU6ZKfov9kYvRg37fTNnDiuwiadg4ZlfTh5sz9XwqT6i7dFSFBl+vFzk0KzyU
r0KOf/8d13aRe7eblYmQeNazazjD0lGVHGgAhBL14N7R+AlY67gitzfTiHEucMfMinsllRWwMVu9
cPjoD+yt1TvHV0DAkmuzzmr0tKbMJvlpyBKOxj0KVovn89rzr4bDgKpLsiHn0/Xfahd0DN4m3cJi
ssC6J57HnpbeE88C3e8mM9DMGAnq2Osf9U32/EkN/dguEZlUY2s/4i/lwJGstCkK8hZe8llX5TWB
YwN/Dc3SS68Qx1JDhoUCQD0/R6CfoL4vbmc1PYDJH31gda78ZN56kXheJroTZ7p9hOlIMJ7WR3Ia
88afLbCZLIEpICNJ4iXWnI3bEvKYklXoCnRnqTlTj6oH3bmXznPx37JedHKErGMrLJySwJOgYIv6
OZAj25cX3kdEI/Vn9jqiQcm0H8lFGAWfWKK0kJ5WegEDwzHQyyQqmzkPNtl7SjEBOJT3b/S1FUwN
5Drl3LPVx9sa4UdLghnQDLrpf49tdmXXP3z2CjkaXRcCU/S1xAMZcIH477C8YZ3jlr0mJ96D6BBx
RuZc6eNfiQJ0f1S5TIC6/MGvIsFMWvjOiUQXBlbQo9kAa/oc9l7TjpOFeOEm9lTfbEFAz0iSuCuH
ozHADYQU1ZrvkUCHKYL23P9Y6fPDNN8buBHQpVInh05ZmR1yC8UIb/xXJ45hsKpxnqN1OkOcKKX+
Xisem5FioljLtTp4dMJKOi55c9wv7f0LWz4XzEOIiBhlAecTIfyQvJPC6Rcjw2SBGiU5KXUg45I+
5302QvdQ2GrSgfPMPG3I/ISuU+GRdDNFL6LYDqQqyy3WPAAwkE8KTS/Yf4N//5/hOLfUHkT1Kk1n
oONtc+cY0sXNEcqPJ+prCB8Blbc7t+QeFfpcMFqoh67IMcFxsTFBlkei7awFUauw8kVC+UP8epkC
jkNdEbow2sr33jo55gEsrV6XQO3RYQbu4G2jmFDxzQCmCnWXgJqzWKELNtD5hpFevXqNtk60nIAm
SKLcHyJzIPLjMzzF7wEQQc8Nd7n9Gy76ZgxcTLilt+vdqiIIHsxDGaA13nsdhwoIXe6T5A88EwDo
5iIdWw4/NFbcGvawMJRe16xhUubhikOvwYvdtmAX3BYAXR4P5rxNvs7bHXpPn3xT++p1CAEB/kcC
2C0kv9jt02WqNxsGzZXEI/2+VjYvp0EHce+b6LTswDc8RdUymFw9st6QlqqraU7Dc7+6NzHtNjf/
OQJIqleogsi2E5PwdVjarmhGLBGPK2dAv3ZNsg+DDshRm5jCZAvGiVvsBQGc51SpT8sKNSY1bwN4
2gBsB7UXA3Txq8pQGs5BtyHCQs8JMsGd8GGWchQaZH63ZvB3IdhiXY7oSnsfBm+XtgoIhSGVzF+0
bmmEbI77XdnC1efQ9t0keV4EjZ975llEWTwx+q8caGuq7aUlbFznhsyHXoGgv99itcvyMArFJTY3
e+ajzMEeqFZwbRfxShQ2N1jh7V/wXG4NCDcLhiqmqk++BUEbokfwjyUVLrzxx1tGS8Vvb5CbQ2DT
g5iWioIN95V9IwNW0C1B63m1yVPb+R8cNAVUs8ij0oX8bzK2wftlPk5psGZ4KewpTN3bdYw2c9Dx
LmtNgqew2iSVv1Eq233aZp5YPQvnEh58gQYUUOZJMDKlO9kap3lu5jLTUqPKULZ3jJHloOjLYkKn
pPwGlgdj1dU9VljnLOvf4tLSy13KLGXYWzHKLMw8FbGDRSCQwd5nXXzWelT/W2vysHOuH20kUJIs
BEStaQT0Q3KgR09xw6OarKpeMtpx0Ng7od3+ebaXJizKK1YNoVgkhEMAQpBSW9a5vq6x2QL93csh
yOD39b5znndAVNsY3JuySCqAVImq1Jymw1tredGr+/eTdMGvqMBN6cTSX29tUhRJwFk2Xcq0VPyN
feOZ4fozlYVgWCSOLV1kW4/SvUXv8QmX564BuW715zaeYxO/0G+IaHDmOXx1CqOLAB340BMthw5c
XvXQZWcepUrvIOcRCBv9HgNG4roqUdSWDgxSyq6W0ZDg9NdOf9xPEGyWy7ObzTuG1MY4uQhA30T0
bLhj+xiMXvanNdzV8WsgXe4BnB6cutTIth+W7xRgCyI/v1kDt9nRQyah7fwDjWUAov5TKqBTdxZn
agledDAq91m6Smjq5Vy4s1Zn8f1HdXNCwsGzdP/ZCdYp8CtB9PIEZel6zw4c2I2so1cGBnDyxNQI
vxE4jNcBHhlq2iBYF/LF8Mg441T/HUYS2ul3dTvKalt1wZf32TWRhebtUgaxoTJmVzTTqWIWYZdn
Szfs/120+addui4JMTkFgPFd7LYMWsLvuydaFTnuwPmCOTx1rfqIrUWf9L42SP+rrO2opWdTM5lr
4bhImMdwkjKuzFZte9UWidDOoEowqMvLBomT8b46s/OMY7/ev1C5mGFtZISMBAlLOj9cOs9fSly2
zYm13nNrbfFYw82Pdnd7V+4Kb6Fa3XK7lPwbB94tpp3KlJ6jKpyjNUY0TChuwyJnUSXoYWz1EUzf
DQWZS65e4fHSexU+uI8RyYcxq+XAPhZYYJs6NYpoKPIko0rgOa2BQSjc+N4knsK8EpW8IRr0KlF7
fJVUjxIUwFP8qrj1lCLlIndKSAhyhwmv7M9ISSk9Aob22oNcmEYCBuVLjJsELcGdoSKmKcmkc23A
L3eakO/ds2q9ZSsyYQfYs/elDX9t67W8zcqHUaRHGgEteT2GH5OmznwZIBOCi3fN0k0wqP4SUr/5
TGRCLsBFVWvfZi3OSB6MkbFKY7Rz2qBR11Zq+ZF8F76GxPm0KV5GHs0s29Awbje9UH44zoxUtQFK
6nhZHZWUB/o6dDpvm0C44onKRAPVdzhEbnI51EZ/daNBN56g35mE9caL4O8xBQvZiwonWY5I5aox
7gx/WtzJY2t6RvexKpPE0quDna1C6q7B05yNaU6z4yegAzO3und3R5xNyn0oWVooYdpFV9USQY7G
QMQRNbZuODPOVemFEog5cr3Ggon12qz5N6f5lBnlPVBWsK7wGt91hC+LarLb+Hv5PrS5oxihonSM
ZP6KhehdzxEqom4KoMUy5u6NZQLuVn8CkZxHiGTlKXWG1/boKNtz5q/xoFUBdCWrWIdcXmpvsgmn
Xj0gpvqc0r2g1rEW51zK99H12Ap8Vbtl3QEfPxGlKp2uGL/zt17DzM0h7NUF2gaK69lRf1caqiJi
pMywnScK7nmJPtQ3AuClFg7s+MzmtnUL6RyV+1lURQ8Y6i+t8VqKKU+4AWO3pXkBwH0GVEBz6SUC
mSc+mRRdJd9tQH9fFt98gbxF40Uh6n47FPYU4Ros/QP1vCStJZjA7YK5xuGIBWHIBS2evCLsR0lw
2/5kFW0qiHODcNd6JJN5WN80BZKUUJMEoiE9PwPnTmWoELR5h/BneHkY8hENATRG9/fknvF0HMP/
HIVdssNTqYJ/xa9bl4DmeOOl2+G+t8acFauRKNal/xTjrMSB6c8hK/cfCSYUgsirz79qEMbkWfWS
9pp/iOdsJQHlgSjVoQP2M7h9XgY5f8kSJ/xTCFB0hr/+9gExA2h/o1LymID8BAedpIXmy+81wB4g
UQGGcGZ1m34PxKZ8PU1BIx5wcowkET4L8vvXmBAqAo4tHnKKeljaGhWdyG/zZB6GOFV8sWVrJnyd
hURxM0eCvvC9wFoEgAIinUlYA3rbPV9ZYyl9FFletkhJsFGSg3mg2RfDW65K9dwnjaDIObC63xKA
pBkrLVP0d8d4QDQGIVfFwnheJ6X+Es9BoyVRbgrLj8NvCJ8WpKHLBMR4SabUJZ7rEkLdLtWQo0kg
2Pcdl3INMgFcjvQvY4aYCKfmXUIptIbI/QxIwgySh/4CwN0Nm7GfsxHg0c6RXFqKQxOQr7agkHMY
swPqHCeiZLSLxJM2g2yQnGJ6ey7M17DImdW5S7Y4NUb3102bsivfZrddjoH1dC3Kckkt8zlNPtmr
R1RljuhpOBGLi7QnaPN96LP+yUH6sizcRH5VxzOXRexi1+78jQvSMGrI4nQa7LVuIn8EEocNPeKm
8ClmNXceDjzFChphYthwNhz1iqkr0tgiEm0oseRBF8Vz1yY8fHvwEvU0lV8bQHiMNsr2dLC2bZ2H
yIPv6CgHDWd08wmpjQDlDWUcM+wuw+bRW1+1DGwd+UqpvaZNdveQvXIoAY1iMbyH2MbNdxWFC2vQ
6vGO0hqWQ6A9iTqFoWdT2I2w6qgZkLT4fzRyiZAnKprhIxOGa+Bx96qROeuSJSHegO7SMC6K2D39
ch/J9y+L5tClhbVAEe1zAyGOME5IlUArTWAGZViZE6/76SpDbtiRzDPS72pxYer/X95MAuHPcBQg
j192QzVrRLv+rCiJpibTBJjmTQJO8oU9Je485j291jyB+mZxCU1eTe2EakpW3y52KD9BO0eccwTj
gNFHL5JTjUWf95m1i7G5EsRJNsz4cL1NBXSr81UOlmSLUDbbvTf6h3c9hdfw5l9qjDBLzGplFxyF
8Nojw/1Dmy6F1QzIHxHSVZQEjDAWvvXYJYKygMhmF1t8dahK4pWS5jeA6NdwphE+baHqSkpbXFIf
954XmdrwfdYEnCBVc4k1IA1/gcLnS+rnTe87FLJneKzLffitZTybMjiWDcdWN8ILQIEAr+p0ZjRk
l4yO72Zt5BVBkQ7KnVgoJnJ1NraP5uwdeboX0mwDDCe2zl1juOWi2TszDa+HXaPLxTa+eT3vaTIr
ysOYRd1CmQmt8ZrkyTtdL+NMxV+f006M5oI+ToBu4t+/OoFVy9xdFpbB7O7mrWGmNe3WYGCT5ZMH
NDVGCYl2uK5KhpA+L++XQ9U8BbcqSZbYQiFAvvFHUGqrEQJVUXpDdg6soiySsrn8v2Xl8kLX1nLs
Vf60svXsch3+ZkdbPYNcT3LrQ17YAx8cJflZzum1Nxfb9PL7kX3s02p6w+vVR3d+QwqV2UpRDD0S
2hm1FnHInYDvD1yRnyWovq2RGb/8koOI2lySgPRS/4k7T3H6Ex3HOytzj2OS+Yt88nVy8BEECCjG
+2UdWippFQtUY5Ez3e4ZTcDRajRT83T7rUDT+WCJqXbB1iu67zVBMK5DqMIpO6zBnkAEMzRXF41C
2GCbzxcYBNwrpKUoOYYNYZjVFJrkwlqslFa2dgta8WQu+xh1HgpAx3S4hhSztl7Jvti4+uEEa/an
FXF1SlfGBC3Pn1B6evW28HovwNzCxA0O9jFiIyrF60hrda6jJRhJzHdOwA8T/y/T6CcDEZ5ZCDK7
0db2t0lRC+3Hv/a9zEVae+Ztw1pvjIPvJP3dv/VcMH6WgQruarKpERvJNAkOHkGyNHKrPJCLdg72
g+CWbQXQwCoy+xNhQd4dpzR5ByIVakWFgJCLo+t/ej0yqKRNxVjAR8co+aJGdXrrvjxIDGlqN0/r
Mw8gmdDdHt9DV4wxp9eviCSFKX0FjKfGIZkzZzxl2gDhLFCadoaBon9ZmXCMzbAWZ6kR+pPG9aRA
+5dKGOAv/bQYTI117r8JC/fF0TH3qD7l11YvpbXMelHKdK5YiODbi57ZotAxRSQmRzLUKo5C5OfV
DDJwoYIOZYfKfNtE3ALzzdq7Ywh3jpeFaGs1aNAC1Knea1Nmr2eVBmKztutsyTx8twF2U4Iu9+8h
5FyDpXmvXTX0+c4P6cQ/rMW2IOd1o0+iPu4clQ+VJZXJaxNFWm4efu74clwz/WVVva4orIzLeiNt
RZ9p4RLzMHVsO2NjAhanud0QJwOLau78TuxqfjROu09IUF8fxAnGnekIwo3XKJtsU7Gw3IjJxEli
n49RSMEVg3KQWBS010Je0l0MjjSqy9axwIb+0t+U3COraHwVMStvk5UMWiitq4oVtt0zcdGY7rjC
/bBHMhffIx+JQ+/lJjE007fBXjb6/Nrb9rISAVGzEd+etUWiEjeWYMDbnVaOVtVKeSISXTsBaXPz
GrBGtocLMPdatf7lA+Ivk6Yj74IyJJLUngPYF5Wa/XyMGb/s0gB9gj09MXrxuvNFpGiwyyoQ7s+Z
pLmTb6swkWhMsJ2vyl2OZdoy0YX+uvpKz/qZWVj5S3kwRU8LuepRwuy3dPIKQMv8zSB4jJ40KSWd
/6M2uYU6gem4GAfElj6jdd0LwcxGl/4nzcpf3UJfDFlo7mohrP1VOdGxs79cdCImb5MdTvBkFyg4
a9pEgqMlLw2CK3rBXEjj7gZerzgcj41AQGCXe+UTFQCIruMwcjyRJ8DYC/9O0U4Y7ne4v4qJbHYp
c2k9CyP40kzcTVWUjPTxr3pWh5JUByQopep+0gvESnRxPlTIT2pg3PmYXa2TFZHsaDBbPVCX06b9
oC0aVjxVETnXWJncaydxxsQrmHPcT//Ei8U+CwodSV66xB+1VGCuEpsNOjCtsAWN6BsQ7fmd5Djb
hxmKwICsJH1g2imdsCPecfb32ipp+9lLOMbBp+TERLp29FBmwoq+F/TB8hTHILo+GGUvkNl0OATh
h6QXvJV3yRQei1S2P3qKvNffIM5QuiWcBOHZe6nYAbRq245S9Lc701qXqmsVBGoM8DgidKrsLa0T
rtFA+NUOy6RObHG48dRayZmXF5Z41+Y7tNJV9RPgQdnBCoeArtaGROVUdIpCyUy5aXFY+eMANZte
JjU7v1wx1YVy6bbtYbyFu1+Ppm2Gv3nCNFZLWfHEWpPZYrnApB0PzaHgdE4OhLN5InUO8XFlIUXr
SZxGz2RVcq5jfermkiGzGJwz/np1nwAW2GJaiHtQsK1jiWsdArFm81U20g0ygb4FSoHRZaDC1vew
rEG9zS+3fxH+A2AqgpMl2bttaXI4AhLda+Wi3SIYOq6X1dhvjz1ugYAwTCiU5Xv7s4qEAjhcOKeB
REBPDemSNXnG2zgJtAGHi3oDj0IbZBfPzEpozYZVxbBAyq7q/o32aSMcX9+SPc9snK+n85hrbw2C
goeUZhF4Ba1+d7H4L26vsyBll5QUkEW2TA0DXG2+MoVA+GImuWt+swimoGYyuesS9lZSaiSNn2WY
+7l/iUuw6Z+pviQRM+S+QAV8R9eSOU0gqm7fMps+5zGlpVqr+/wND5ux4ixU0mj0BtjetM2tl1M7
KrFu2mnYDs4mzbOMsjRPC88qNPbkMQ32Wmt87d3XMrwqQZwGrht9qYLUlkPdoQ86hKAWmNuPQKto
qwi/FSnwisp50nJY+qCsX6Dap9G3h/ILa7n6eeHtDP1TvP5VsV3HGbWUacaIh8qDpdq7gM2NWPaY
4FZaLeD9md7YO/ASivXEQDC4m+vt43JhH7+gswV/rlNJ5rYbmL+mnUJWDp105gQ/OTMIxZsX/gky
OCrV4e0ovXlYCqgwbUYvWwaJk20AA4E+exAZttrCrUo7PDrjwtJa4hStbZ6y7nAOq6rk545KXSJ4
MSGKpoulGt/J7o7ci054NIRTifNYt4Xwr1J3pXbs5votT1h2t0YWPmLDHpmOqJrSEfn5r4liyEz2
K9ZCNTt2aAZIkOyFVO1zhxm2kO/dsmaJUpF3O9h5iuFIkegQkhCfFMkbQeAVRvJ52c8STgJykrv7
NO/Y0yJb9HnsrlpMe2/L+fbbWVhQw6HmRYk9PyXn8p9fkS7VWXTlAvYDYiCVHcYaPgO/ZozHn8xd
20yGpk30zhXtjEW9cBy11lAHR/jHnsib3+Rr+a4ofIoh7c59ydlLTmaOXuroaD9vfH3trl0aajIb
58a+Ol5sB98CqBjtC5vDDvbUetI4bB4iSAWnrhSgrUMtCncLWnLumBudWiv6/glNw2cVkr+I+I3M
g2Zv/2Ta/3HLHvp6knccVgbVa24BA/iL7n6lVqclvu+g81bfd9K2OE8tLukYxiCTjnral1HBxG4p
1VBFRZqlNKu9YmfKqp6G3XAkbsqjPQlwSyeiN7WWv4B9Gpr5QIycIJ21g0dcwkwoC2bzugIMZO3V
UNLbea1kFpv7ycBCC+tO8AWrtSB1DAfU24oEmXwB0vdgcblb2D2vbCqMoS5KHoAnI2wW5y0/w4sM
LXqzou1HNlUx630tVm8roS8N9t9FOxO2tL7/hdqsO9UfiA9TFsSZ8OYc8CWF6ndClP5snpPBpbwq
dzLQ32GvbHjGUW6FpWsF6SpBa7YVJJEZAjrtHEsQqQcZqJCwbc95ZVhietfSvPUHn8lauhyTgo/j
u1zjQoZJgahoncDWbllbWIGVCOuuk4e/+PGPBKNDEHnPH6dZZ/YivCZd/T8q9CBWe7CGAQ4eUR8/
p+cDFR+adpEjZz1NNaMYs17zvZZUthereQ13bGl2YHlkCTor3ieKLRgJUuDK68BGtYlsDadu93QJ
efxpWgLfhliTuU3v4cQqdI0C7BBgwWW4xw8FSjvREpt83QvzX55rHfzeCx8m84RUivZXSndONtIL
ttSbbp0/3//Sc2gTiBcmZLADvMM+QDdqBsZvjTptmueLFN8PvrOFFi38aZFCXzWjEXZbx4AwUtmq
rJCUddI7+8NQSbzfYFv8I0h89kADNXbGNV6etq22oq/2lYLRK2b8HWFEhA/4ZAIFlFXlhyhlDHhz
yXdKfQ5X81Fp2OUKt61Gu148nmUcbd9hSb1UTc0l+GTz8Auy1UoQIxXxP/5Hxrq2JaRoSLiNKJBN
m+C3zom1hYEYPRON4pbsmokW5EvLZrClCQ5oiv05xYpIdBXaQiMZnTSRYTqcWvrOzLaMKw8gUt5s
oMmWWfj2SAG1I+tkAA7X2iMZPqKf7pVikH0FcDXH+TZ7MstmMzc6ZMDg1XNsWWygg/N7IKxLBlef
O7S126Ga14oFzJ7KaiKyJGeKZeaYQgud0hcEKI3QYk5tohqtD0GPy2BADgpXktw8iVP8QD4xU/tD
vxvaBSxYyo5Frj1oEq2iz8cC/+0OLgla55abajlD3HpPqA6EXXwMsJDUXeWYlUKqo7C53q9C1ugU
6UltOVQ6flAF9y+iMK4PbeJo28d8N3ks3705ujK/+Q2EjCgdqgepdrDV4bTvXDEQZ8Dp/ai/uDbI
jn2mXrmRmRO3XnntC06V+iOqxpdx2iEAJJ7Vnwq8fEmnuoDYyj+4hTOR2B+/QdhX4xTPiUE3TJfK
W1kw2heyZR9ThqwuseTm3vzEwXDTpQbXZGRYQdNSZk53I58Udr27nnOHJXcvB2G16YqRSiwImtQc
MEVTLiVOo2wfJpvlicymBZuJgTc12zCHe7YRMXVGZ9soqO+VpzZRBjw9eFPgo27CTEBxYRBrGsIM
kV0GdjCn4ySwpbB1H+6ye7UmCuIe3qGgkKpyuWAYjySQqVMEBJk/vEzxDM5Il/0hNDUaPy6EjUax
/2aUoEVKYlmhGpCZdeGFaRbCMvqgwDkNaFoQSGVCgomaVwpVJeN9Y4FfSy3NNoE8vW39nJwE6YUG
E1ODrJpbgPl8PV2HpxpsKjOP1sipar86mhG1DB1CVcD+WLTYJoEEMdNdTeqD4pOAMNAtIxkaLZgd
QQ9ePbyiR3WPw3jfa32Ck6v7VyueDt6aAEB8ZXlRqar9V8zJih0mGRhPerH10ymvR9qMcrr3rD+j
pXCDGV4lpLn7KwJ4zuwdZQsK64lDa4pR8kw/1T2h+3F3OIo4QlTe4hkb0kgOjkRkHE98TUmYBjeK
CgILFh8TioQrPO+hDz1qAiWoxQ0TCu5FSFcaTB53g7wVViEhZsJID7jtD3paRUt6s13R9HoW5j3V
8+6O4MgTwm10PciZSz5EXtVxf6OtmvrvlVMyHj9NBl5VZ9D+VK5i9Tk4S+1tQJjOsutReIEoeoIl
dcVC3lAhp26wz2YkrNaZ6ICeV+zTJ06gcifI6bvHL++zvPoJQJPASyXj4gyHk6xKsNg5mTXUINIY
sX3xXt6vNZqEvAItGrp7S3PtYc8jHJ0lPwRniSJhzwZAaenuyz2BQFmcFRr7pLXj7nnuoYsUh4hW
YRnuXYpao9FsgI0QKX5II8Y46ZrwBjhy6TAR8DFtccJDEJsU4mwKbCiOH5JnWLrxIjUDgqRZPJHK
MzEtwIPAUhRN6vjXSmDzj3Ik48WVx4j0zVG1ehSk8ahtUAiNhv/rGfmwsIHRmm92WNEGwDfocyIc
3WzXXm384iJYtdi7kg9D/usT3Jj19ZQ7tdKllkYE2pDrGGEY/MW3kg0OAJR8LNPuZNzjjLsYWYD5
qpdDSR9xy06Mq9Tkb18x4co8PAeWUzMfKXw+XsRLnjKC93mxa1iv1sqjCY4lqqaNTriwtrRsk4PD
bPJ3pAuIe95Y78/340+5pjnFKNOZLpLAm9qRKg7OcwsKW9CzLw418KW/ako6tsVfiSKt/Kdu9dEA
eUzziGo8F8jpnsgmKXnf+fJuMA1Rk3uvDJLvJhx2l79rqfx3jqUX6UXCqbfKLpW44hcY78koVNhI
YvY8QOyJnxmwBLdw9B7Q5rCPbLkWF0LxO3yPqmf1Gh/lDKKTBhZlrb0pUpyF+R/29K1HNJUQfa/s
c61E/JMPEB0WI9cUOYKpNTb/Ab8O7ng2j0MDkvV8e0mtkTaOXl9WCjXg/RK6xMoYrS/AVHzgLth8
/uFj6sFWSqcgvSV2JkkdqPJcj59J0Z0CEnNaSSRPudH5fXYA2EBVxJnBCScO/4SN/yizDUizhOCy
k3zab/Ft1H6Fb/WTB8LhZAxnqSH8KnKpaDVfKtHir9ib6BzGCGWgHDK/rGMkAIB+4byQywYQmdZp
s9EMP1FOFmPe5OsJXTUvRnmIcSdcqT76lmEiRNf30dsMW+EP0VXGL/zZQ28xs2zsSFr+DSa0qkxZ
r3g0EThC5ARd8+9AeClxAnDFaCmm+iduvwVH8zh2PWO885/5VWMhQBA0IOGR6p+BRoldhc5eDIMC
I2iMljTkeOyvUNp3pGehnYLJriDgOQjHj/EMdDz2Pq3itLrKYMe3kbRPzmNjxH2UUwx2TYEGa3p6
ck4ZYt2QcKNS5Vt5Ww/4xnhsOMT+8ltb/RRBSO98WVFXU5pcYL6bGf3LmOMpRcRYJx18K4105PzO
ezxk8BMt/Q2ikUeFhXWhOLUNlwbo8h7tgPxmHceq2zT0+EQ/rJq6mfi5uZ2/KEFqtusJTMfcY+Mv
9MWypkldLwSW9cqVjB4IXJLMGXvrYFf/FCSAzcpR5Y/K/yeZyZbk3wIgN/zgidlqfiYN41+3T3Rr
/IEcPNR+HYhQFf3NlRqeoJKJk7Hs/EycEQZM9E08BEJXpkBpSnS6HjiJ9YthSUVIRr5YI++pAEcO
uMr+qZtwrCMyhu+PGxGfSlgMlN74tIlkUzhys9hQQPcDLnAn0z7nu/+iwqkZn22C+aS8S0t3LVVA
HrM7FLYwFqPSfu2ygYQJjevXgZAbXqpECailAQodQb/oAjZyclEVXb9su3tOtkQNhvKk4CwuzNht
NIjn1n7tO440dYtpikHgcQaoF7heHvd+t5Ua3UJcTd23y3L1VCHHitO68QIQIyDvBZFuXg7v0+6t
n9gxTKAFrOwKLKV48OoMIMTuaQA0VhHrEtOEnXc+vCDST1LZxgT3Utgg1oSiL1UfSfVGJRq60jKR
J/SenH7K9MmtBcrct81ilew+8r7UpZRnDfTrIdYjWVDkyui7Q4zadvRjHXs8LHMOKN4T0Yzvrngm
17zcSiwit7Wt+UmQU9ZKRLcGutjIqA51t97d8AXmRmBZD/3061CpZUEEXFCaJXMZ+eStwUbxBpHL
4Fva6kVrXoUD8QpD5YT31DA/J9/+16Nlk+Pw3Z/UfotDEOTDD0t/Junj5Dk11Ow/NZV8AuHw+YE9
dEpliBzzb+b3Pg/xnhgkOvOfHeFD5qQfGDPositWSobQjuPgaSIO2PM/vKJXxGo0cJLFEBGszkE5
0pilfi78baTr14PgpF5oPbTfod5vkDbGCDyDcE/St8ZN4eSv/U9I+S8uRHMOCahNPaa99ZjbyeBw
BqEnKBYahuc5oEDVHTirSIvvuUkI7pWbGp3fpsHnOsl2wjelGx3oI+LS3mOdjGwDslXxoMeHlcs1
9CXZNobwHfcq4RV2bG5j6yA/BQ+SVUBKdH4Ha+89D55oz9m5GXzRwT+esquAYALDa5lixjtpnrZX
QeZD/WstYgo6ZNGM9IrhrcZTR+X/0G+pwUD89ntsHTdxM7dy1+vFCC+tm1UNxcsrJGN3K93bbl7b
2ayOzIcuX0XQu72UN9fboPjOa3bxN/p3UPjebRKq3vbcxYnQetX3JeTzL+JwgtFBM2Ia78dAemEP
nXpR3dFba/7uRYRMg1L2myFz0CPHP1QM55fwK4GMea5gad4SXgW9JtzEefBVwbwIW6YHKF6oF/Sj
I3S1VKdWZmTAdUFFylvXhUsShSS7rrTYhT7kqiEeL4QfWNgFff/47uJXX48Vqu0QUNihoV/SJwgR
92I3Y/aKNAfbKR5RP7n1XNSvd0eGoR4/3MCxZ3cwVe3SESAOTFVeGDJo9mniHvGskzooFVlJMYdS
XLzfiUnxLYLhcgcKK3j8TwU0lAPiMQMBsTzrLGV4OLv+GWJwqnN9nKHYRnWxu4hiaqu+D20mzJt0
9qn6efMtSuklvP1sCC5SECdjiZEAqg2q5tNkVUNjPpQlWvV47d1t9EoiFPzco/5mpC7AwyzxwiKP
BaWaeQoMRLraYV//YUEZcZhFpAnGu8vcWF38OyAekTMZhd7SP9qWs9JiZFTENNGdX37BhXqy3VkS
LW3iQOLdxN+EqM1jBQBD4QXLVElBBVg+4zO0LO4JaefGFaFI4z/1MDTxyaJMcPK9BnBFrAGVE4wQ
aM933Rd3kgXQUzP8EZWEf++kRVOj2m5H8i9voS0EVgM8T53pshLTILOHZTL6bw3NTjJqvnAEyTLu
yatnwQwlHtAAlNRM7+Hs4ELhMRsyGyTvk/r0azuA/E4K3/ZpX7Csqj2EvqYtAo/cipdNFCUep7yb
fpzt+YMDG86Pw4WJ7Qw4vDsZKeD/VL8Ce6n5b0Q1w4SDIwZurM6KtxXN4F8hrPloPh4VBsPvzebM
4q3ExswGVCu0fXeGV3r/xOVexLA4q5sVAMkgj4rzh0z5A2tdUoV+ftF9N1OKFFAHIyzjDNW7boG9
VryUGuGeAYLzu11SiskUByp6u04DkkHx/zsszkLqtc42GisO2eY1QoNX9cDkNlEsjZxt/4WqO/6U
nPeKRiQdtAHsE/a2vsD17bccQtvXuLSXCJKQ8dbJjCZctptURBdkHbQjdFjWuXwfj2W2snG8avEC
yAl7OfBvjp6r3nxIM4d2f2Z1w3p9u2clZECyTz9c4zLgxVxrIZ+byftUmv13l2wfXJ1lfQBZo3AA
UVEqLo17z9YIFnE9pyTv2EHIfcaMrOxilDGCgVN9642yBOXWhOkLUaGVaERivwzo/TLC4LxjJuGy
zAaNNY1yuvZuPmj+qc1+tOW1FldWuU1ZXfrMYHRe53a/Keztnkeu4+YSGZIPMX+tdAPy5+GAxXLJ
fczIcmCTKDuYxWBfNpbgKUmfMtJB3f6i2basAwHUwwieUlc14gTJNCIzA2bBNu7B6FKaoq5wjyXc
W1Oygf5mnzQ6iKHIvM94GmXyWV6lQ3OvBZdW7TAO5DnFbqi3jnnyiOpZY2RarWEk5U28PZW75OHN
DKXJI5lhp7Lgn9QTsXPfk2anypzOX2VtHokmWH/zdEbEJ+t13rjd+QfAwDlyu8o8nJo65xLEslf8
GuECsiTRLY20uVLbO6O/VVM7C+O+i7UWggvCS7Irb/ol5BGCk26k8Yue9j7swfcKhqRFeRH/fUiL
xG3OQSpWHVWCbG5mZKp7NTmFgES/446S6pzfT0wv8xBebPjNKb2CMFKG3SoLGYCqnq0pCgCovcig
O1Ky2P9VnBjlH4EJnY8d9trEJGy06iWjteZH3IqLxA9IZB2GWZenyziAUw1e3aJF5e+OSEjudWYi
qWnyPUQU6wTBmminSjzq/iePsI0rPlHY5oaWW7bJmwYOekY8feXyqegalRvokeLMwwb7eJii7/uv
+MrPzin697HbI8RWrHRP/CLCM2xJzS1SSIDSxsGgwQkLqN6XNhSWgvdWDMdO8Y/F591nR1eZAsDi
Q+tQ94ZDYtc44aBqbNqR/bIyPkY+Ofg1c97Ch3OfIMUkM7imDWzwjSw3xCaE8uaWKJo5I5vH8WaN
UjCbeUNwDssw4E9OK/lJAbPbPX6o4diTWBbIZIYJ4RlxovzoV0SCWj8ys8GUtR6U4DTwDXMtxYxL
EQoyYBNvwIYqEVT/Ii62HbX3PE80Rj1aT15kYuw4w/niIyj+a0To9vG8Xfw3vFThs/TNrQ6j+Wvf
wQtba961NUdFJ8dlqqMHp2YNaCumIsT0xqoNhF6Y7ZNIb3Aq5Jg2xkRvPjhipZeUC6FGPI+hn0H8
f3AGu1yXrGv441NDTjn8LLXlXk7NNZheshd3MQaRqZAEaMlkMXCdtM3kWPUY42+ECwxHkRrwO9h8
mv1HTB0BPSOF49jGFCwTiH87oXVj45Oj/rZ6tMEJcOnjE6FkGuH7uKQoZi/7Hkp57yb1WVQjCjd6
dPL7iazT22l3TNiRxjVUegNsvMVTERsSFdevn4+8zal1zpSTh4/blDYnhAgckIUWOtUbj6Lqn1iP
CbXL4K1w/4Ay4jdi6PZu91QuY4v7jA6ZTMuScmGXS8h40btrKr6VQ6ufF6t2iGwsJL1zyqvoqusQ
dEgQE+cZ5CdgvU5PYJlDHhQb4c6axW/cdahZlT5+hcf/PNYDwSUDdKPc8P2SK6xhUHreDNhcYgkF
lx/LWEykZ6oFB+67TF9jiCn4f13Tsmf5rRIDa7Y4Bmhcm1P/rJVk7fxOfrCBE/INcoerkxf4kHbP
bc41zlj7RinVq/n9HoovOmhwMLM3D5SvtCU5p6PfH5rquCDMwLSxMtjiqOrhElYi5E7Jhqwg2Nm3
oyF1DRnBEaG0UVS9GfEx1W887W45G+YVCcCEyGZOByll6JAzgvwVhn5VByqCQZuK8K1vT4DnB3Qi
yI9aYWFjxm/WqiW4ndAI1ysluCHpanWh0lZSSbFmMC/HzCRhkjms1lBlD7yXTwZCxC5w9FaJnhf+
Hl9gQmoCvmlO2P6ay5J8HX4PO1iQ+0QBCLPieVzxtOfEw3x0Pf1jVb02HXabS5ElDlEjQueM00RN
S/0B4DmE4GRdsmc1AxFxm7DeaPcrU9PLYWW5IGFBqUokyHdIV6K0f/QY0r1n/vnE9aS6Ceubt5H2
/yxxEik5xKmX/HhlNhxnIY+LMs6BXUoB/H21i3NsZX6LB2YEzyWHLwaAi/afO/OmPnNRLg125615
wmk2o/XMw+ZgXSKSQdQ4DYnLEkbFd6IQ1MVymn+nNhi+xpqkLYNsNqYG3RbLUB9f1vtj3BzDMUWc
ldDakpyaICtWbwVp5StStSQ6inDWRjm3pGLZKYLUGElK+uIK7q1dAk6c+c7h7V2W5QcB2bhDBLR5
bsntM1qtTF1WiRpbgzTDbWKBySfhg2WM5IyUZHkgdZpFYC8SPbWsVWbLFhTRcSbIn/ORqYZVWpTw
/CYj/U2EeOWZo8buksAvOj/Ua9cr5wj38ONUTNuCybOmRxbnM+/rP8SOYlKtV+knKd8xtSnxvqYh
Pp0An7Zc51vYOZZM6wHV0YCknCftf6umGNGfJz4KlurqOTBLZC1d2DrfBwXiM41wRCx9w+Sw9K4/
ZAm2nbErJlZDbE3V39bLURJ/4YsrQ7q1v1y0/EJU5meVXNA8eM+SCjOqGa8ViwmMtGalnDO249mz
BFh9N/cYiWoP3yvuz/wqMr1VIIG2D6ESMSx74vtx5w+QMmgzI6jKaDnF8rhle73+q5e4cIRJG3Ub
bpffH8qTF9HcvtTKjpQh+yyOMqoNPlv8ZPl5IrlbNrPEC0KeehXdOUz+yBR2KbJlEFD5Q65XBZ6P
Cp5CMufXP4z3OkMVwgH51UWrzoa1ii4QUB4PwsTzW4uyKwo/4P2H8JS9+n6ni61x37SBJn03Njaw
Pq8BUHwx/uuXx97W1NAe6AFcg9V7nvNz+LgwdGcCH5Y64YtzEodnVusiDM5bAcxxOkA1RHIsAsmd
bsTT1mbxaxaklrL+VF8nmYhZIEJQFHDfw8uZMyYEXWAmv4hXpIpMqFoUXNCDsbRji0Uzb8ZZQ/x9
iNHWxgiWcelbVYoIepjFP36aLduwSvKEC5BABc14NstEQIeqGYH+jSwMq0R23jS+m8EUSBJNrMu4
juK5U6iUgAX/lMFId+UbMuR13MrL3JO51mOyl4s+NOPJJ1kOAZ5kkh4/uVl7uvTz590R7teJ+EiN
2zfl01zKymhEzLzIB6al0q0v5b8H1slzNrtkz0x1Ha1zhC7obohw2Z3xJJ29jg/snGB1GGa5umOi
dRY592y1Q8RH+Eos23FHBNqWNMzBaNziJp660roiQngKuIPVObw5jsiRoyinEtl8UQ4jm15Kz4KG
bYykjJvirXxh4vwbsDKPn9Gk4vOjU5i2mrTLPBlp/Bu8Oojdcp/ijZglsj2rbi4DwcEtieToubAy
gREnwWfWqA/H729/qQo70lx3ulIp1+pTMKlvmjcMZ7Ub5On7JHtgaNC4dmpyFXuFm4d+VRSIEy3G
P3cq10s2jucB92MHpmW2/vNylOv340c+t4DOZXpaByhc9VpXjJWsN6l+c25FdwOwI3e92Bv19ZB4
qmE1tmiDp71nU7qk4VWAq4NSfA8x498/v+KxufRHchsQyfh7USEEqi+KeQahknWQq7NZLoYKsiNn
J0iBJX3EIoUoE9k1mZNjv4+dSbig/J6J2sDPy9vrTYccrBiKJ9VlqEd4xddDGzfHQxlaXMIwnjMG
vRGTovWb1fGDqT42DAiMf0e6bHNgvDyOwRfx39r3BRG4mqnGiP8dyMpa6FA+ASQvZZil/Xw2MgJi
hDSf16xI0SX8zCFukt4t9CBnqwXVeYIabGoCQlmbWex3dr7g8BeX13R4klO8/PUgqYW5oAaxXKZZ
q8wLgqkjV9Q5wgz4uSAbojrMIYsj0cQGuNvkfqJnWG6B2/OrUjdS+ADgmEYyGjqJU2kcWjPbV7Cz
QCEHMoRzXB1DoS6/G0GJrDbuHX1Md4kEOr7p4fG03JCl6r5pVkxvSW6bPJt0PIaCZVl5J5QI/qdQ
48GnO6egpcXZym8jg5JPC1Icqpw7nhQQB72DW96LimKydcuPUYnGz8pvhMJktKn58ppGQP8muKHd
fKm9AZ9Oolp7ZZJBryc+MB7mg3m4EohWCBA9mwe44fC+cziIrA3IpikaDmnwUqxHnd4DMphkHGPw
S/xDTpKgmNu9YeBkZLHRqdYmPADSqPXFL4FmszF9zjRCd7VDfOFlWic28EOOtFPyKsllpRbxDLjA
8Xrwk7fk/VK5uVIkDKXA54JuNrfwWFvuWULPFZ3opvuSTRF0Rg4XC3rw0M532F8mFBfDjtgWMBKc
HOt01QAM5bkmL/fC07xkUfLkNWWVlsUSyNy+99myIPOQAPuUWQuHRqqJhKSgQnYuL3JP3YA9lPgg
cKJKlakxbF6QpRLLOw3cTxBHbHdezHmrWEn/41+ukEmAnFPXgNVon4wPenGPxVyd3My7cgPXiVyv
1TK6GVeM9G8AQgl+rpEV5y09AfFAyhAYdMO1nkGnuuVHENyy6i9Suv87K15DrI8kyjJO7FC3gTUt
T0yNug4iGT137DAzBTb3DeRZqybho9pu9oM4xmHS6byeVTBItJj0+turfSZiOMSG+ltZ2HcJ2npU
ZyR2Bgnctf93qVg2MTWyxfN2e13huvY7Q76XU0lwV1hfY+HAMmzHU9TDB7+RymUEn32dMNZXbAIR
SAa7X7v5pYuZd9CUPSP6/C0HHz2gHCiq4lCbKVhRSo8f/2aDjB3x5+y+Ko3EjhQddwe1c+3dWwfE
maMmOdwGSUykwbp9mLWG6dozkQ+EUYV2KfR15UOGmChLXt2C1w7JApvWyPtXYh1oUeh4UQtCTFWs
MNi/JSxl/GkT//wzKrq6z7ffGj+Y6AyU1rZQ6iJaAGz59v+QYCtl/5VwkwchZTy8NRVhbuqSPfzW
0sglnkiljBbPx7pr+UwnpGE6oS1ELTCOOtesUePgz+5f/QTT0GR+KQOVV7oF+1mBG1D5H11qYM49
MuG+mF5dFWXyt8+ebtrukK7DV8O8uwP3pGBP7xQWguqM9phyZOuJXIkaMgbtLY4POCA1jTrZK/eP
ALRMtF6I033HFXS127TJTMvfG9Ky4cS5fKW3IjyhfiDb91QkXR0UaudjNKwvUKsxOEcxJ2ppOi0i
8SYNxTdTqbYf1Rfb6fRRHNzL4uA1kOhQZb8FvJQWmUOHb1VGUPp760kQvtwEdzmcXqY9BZzxMw09
KNa8cnfZdh7m1xpCBYyXATdOzYHPvASrEvz6Vk+hno9mCQdjoFaFI5LRDvxMj91mOhvt0J68CRw5
Ow69/AWYnOJ66Es9GsIxNP5Tzn7t/kS6FH8mUFnwuqUsoiNciFTRJWEZbcK1T4D9yvEkIM0Wn8ZC
CwjmmuRJrhEurQ9uu39Ojnc853iVe+47J2dsdnwl596tevxHTKtEFVkEYznoJoNq7gDCfRufLZvE
r0Bc5uSOf2NicLAgEkZYKf8QwKCTlSdAs1P4qWFTaRvQWtFATHK91POGdQt7E/B1j57eGuTyrM47
E5owL0J8zS3PpechgD545dp7MOwjmcU2MKBiq8JwT3tjD4LAZTrwX4a/W7YIjHx0Tn9lnMXcvKC4
KzKLLJ7JXw5Ls8tO3/XqImg84BkwxbzRhiRfxCbvfqaRRe1QKxJyOVncHVr7NYk2eYxpXPNNnS2W
/ZhYm5DfBLnVk/J30MsnpYmzCyETh2AEtjKDEOCXLTky5udDXXB2/8DUIN0Gq6yP5Kc/Lsi80ttz
VgVNbw3xiQk7mg7SKKB0Snw0gbv9DLRlbRNPC1JZh2FvkMb3M5cHvhkM6NLYC03/9ExrxmI3YhCm
Vg6taGCMTi1IVSJDGWF3xL+A7fUi94DQZqJBL6bUtlNIR3Xkam8q2tMb71qzbKetaC3XB0o8qmFK
PL452HKhVs/WleYhXYsyjzBeENmDfL9A64nXcv57xeUhvE6RnPHVDGpgGE9fjk7r2eq0Qz2RFK9D
XoFcLVBZq22WBarMZJUrqt9MJfIz2fVQJTXSb2RasRngF/fmhXlHUYBriM2yX4t3o2yIIiPqWRQ+
KCfib3uF4u/8ZYb2WkUtcxNaOLOqQywhqXYINco2OU6z4VzSKOH47/cnLspmO7YI3uZ3QuoCEL3T
QmARbruK6H8hAkWD2LDz6mdpPeUyIYYpsZUu3fhzvaiUHQ3bSHPq1JVV9kXBnwh0ODPEn+0mtX10
zAQMhtjJ1FjNkzOQsK4M4Gsw9dF3nQgsAjBHFM5oORdtkh/dt9Qm8glmygAZsrVzz5qAgqNg+1w6
pN24au9Z1kXNl4Qby1yhzwr68nubq/POggqNFFvlGbak0vlLQkvzSFbpYndK1ecDFFvPYBkkt0XR
toN8tQi2B9CntkzYi1XuvZuqq4TXsPEnsbUXr1C/ZK/pfOy2lQlcVT/R7C68pu+rV/ww86C83KDF
AtjTVVgrHVYYlXKVlZIEDuXoongtX+C8U8qMNkQ3LBicA7hE/5hR3ipfe8pJxkRoI9/geBfEqA2V
+0iiFRnPBEj4UU9S24CO1xOIirjgnT8q3Eykqur2sFE791eBxgkAd1VeEdTRPNl8zYu8Goey3C0j
hc0MLb93iwnt/KjrdFVEtGCcM4PQq5cUHv5Dy1oX277N7ugmW1kRZLL4VyhQANyFNABCQkDqz6vv
TPYIpLVCtwcTwhOBrLuDpp1L/yzdHC/3SO1NIJUqOENBbt6eccX22MO331SxJA+Scyn23R5grmg8
MqEyfgITd+PWWdjs9Ki8fuseXFCcdBXXk4oC9E8yBPi4zek36OASmN78toik8+g1Bk5/p97pUATL
DsCfWXZy9JrB3GPLwJdgeQ7wvQgpOwdcyq8huSrObJHqthyXQcJIgVsUN+Pq16NLwI+j686KjtbQ
6/JfU7PlmjznzFtR0NhK10zwrUWXA1YO9YZTxUsphktlGGewdc99Is0iMUkMeWEECjwHXaaKzht7
k18nWdwWtIxFy2Fyp41Ybxpt/aBKP8666kDzeUlTGmQDX+V+6fobCMX92SFelHZmZqQ+ghiJ/Bt4
JtYF1VYPiytEBabGRYhotzQpTFNbVfS1EcmgAklHEWW8sF43Ff3tnuSLXrfyAQiPaHjO7rjIT5L9
XIpPNzdZkHbD1VLwM68BRp8u1u6zBiCXMrrcC0IkzWICoszEUggL38OxA2RNoaZ/cdM/bZaXOKCL
980Wz6YUqi9a8kIGjPtm2zyMKgZQ+PLpAsSYAfDckxSXWzR5wCvMdJh0QaOoH5h85HjuuStJRcx/
tswDJj9+ZA8wXdi1LGKZXaMERAaotjjTIi8c46TAMz7ny2Jwy03pAT861tWA2RRFDbN82gnzudFo
qSGc4wOaZSHBGAffxSjUZJg0fpbvL+2Y5+HBPVMK0OZ6GzB4O7ZXJhfPliYv0VdTrlxfI0fjtVKs
j6ODebR7V7B2yg8mSIpwYxbpx5ZpSjs0yPljcGQ3wiI12WcN7e9Bk+T0NuTAYLP+y/awGuJ4AFWN
3YiCUzjs/i5wKBE4IrKNBYjdIZJc7W5f+ha0+Rv95qMILUQDeS8imeI6GWT+mD2HltrooGSL+xvy
XDe7+b9XsVMFS3Ls5XqgeSy59ElLmZQa83PtT1LYDsGdfoHV195UrxGHYvcILWiM0FNL0kVIzWPN
bU7TFMXr4BSfu8Z0aBkMNfuiRvo74losRvNvil3lYO1mMLuAbae0YJ3JtVDB/2qqj7LsZY5kp867
RQht1LDwa7EOoSvU7jA2xelehO283/3zuB4scbNYcap+hxCkI2Q3N/uvZBYMnsfr8xpyFWKMmdVT
y9a9lTobpanocL4dBmuZ58IczFIXhdlMIjOiuXm9pZ0sCV2qCTBiQn+BPAVUufZuntqFkwB9GC95
PCu2BH2FRU6E87W7o8eQGPeZOHv8oQS0Q+Wb+h7m4f2agSSB1dIjfRHFKJkDjW/0ut1EqoweO/cC
Ko2scH48XxITOyFNgc9XPf2fnqFNG9HEOtBNjxxyeFSqXOL6vAjufL3ONg/qGJu8UyJJx/ddLkTf
wcW4sRBNb690imnjWiIx8eNix6sXi04rW5inAzzgCfFXmMuROCo7xoFvZSKbm/Gwuv9eDk+SPhl2
OT79IDmGODEgqt6Bm69w87585kAaEw8LdEJ6ln16Ex/pg8y+W0C5ULCWBoSQYdo5tCiIS/drgeRh
CqDxFXpLVZoOrogMnuRnDyozCA6YGos3bq189jyu9/cTq+iEDpVIvvWXT+M/o6Aj7UTUYzMSaz9B
csAe+ICmWBKBm1DYY6pNMrnrT37AlwV/O9nCNSuj/AifZwvs7H3uGgn7/RRWCLvI5g7iNauqaOag
RS/JjD9q/Q6Kvn0WQKwuFXF/X2UJocrpHAshdkik5sf4/VYdnEQ7outuUqzlhRyVUSksDvLR3RJa
a16KHkmv1anduC7qhOi3c5vh18G3VzCx9ozeJIuWwRcrEGknsuP5K9HCVLq60S1+8uwuXlGq76KR
Bnz3Xfvc1834eKtoPJOujdIhx/s6kJ11WrQe6eLCYEAXWXLVxyGjLa912irngRx9UrISkVVlKGys
YFnCY1SrfEFWKD2x6i/q5fqJPkLrfVQCkKWGceHHR8wnp/di0dfISnSQq8/+8rk45JlIV4gKPUdE
suTjdkqMSa3xp1wwR0orepetjH2voNreh6rRUwn5X8HtYUvJl0onXcJg/UO2UG4zNsCPGWyM0ze1
CCeApkGDDIDQEYV47116Kc1zqtBeX+4zZj2PZR1zeXyeirWct4RTuixdfd75RU9OPsAEvOMzoTPs
BMc4xadSK3B6h8e/MXHLgdrB/YNhWiEI/LLOMcIQ5klziTKDY+ahkQ/VpBHK5345C9nAf5MAheZr
NN7uKO5bt2MvdCy2LjvAG6HjgILJjpEYpJ4FS3sXBAiMi7X3dwOMu02RUf00o8cA+y7aWrFg1ZIC
p5nXqFTenYs+S1L9EY4s5oAVS5emmQLA7oya8Dj3EQPLtKqjRVx6hrzeBcNUkk0mmaJGDCC1R1Io
lrzi0lwym1wijVdCkscVNl9/d0jHAlzYXcLOL7sdLpl2gthjZYZqgqvvQM2XCQ2viCPjvpLJHuCG
H8si0WCWGxk2oYOhPslXp+6Ub2jEB5eEhaJKhA/6DCOm+z+Oi8Q1F2tOWDhMX2p9E2hTEUtYId3W
9gIpDrN8NHwofm2EpRQK7OFSQvMBmnL/cXuY0rUJMkrp7bDVUH/uykipqc4abXKC3UFZ8GAWBEDt
LDBY2OjaDYxKNvtgUZ6/7daZISWvybvsXDyhmAnqhFi3Bsf5IfikcmXw1daNAgzZHlarXe/3mU8d
BeRv4wAowt6ypzSwlGKWVmhvtPM8MLdNosKMhUqsyBiqO85F0AFY9Mwj73si7v8IpbJMiMpZi9qH
vNQoDHwyxhk+2ZLTURagd3DdT8fjn6Jl7vGDnjwInOaf8zJ1vQZINdtPJp8tczSIsY+h03pQevQI
5D35GxTXCUf63WjDQeCcHYHoJUct3Qr2f3VbZ1rcKaxlrarSSgMAtYrG5IH3Xr0/G1mx/zhiismu
FIRjFu6+E3EF3liq2WiGKARkvC2kNbkqeRoRo+qp29kAfY58AH0/GhvrnIccQhQaF247rKl48k9h
k7LujUS4MvBugVwln3GG2hzFPaOoUMEztwljoQzcZgWgXbqXceMgfWe55WtuZhhheZBz5+KDZmjt
K8OYLlfkNT69zvb2ZekI89xwihykxzD0lSTPAa+VaJNuG3GruoQMpSHV3xnHZZ8DO229XhtC1A9R
KoyOZ2YgXTsOit9LS2FWku6NFQL0CC4nvzFQfFnZWQIZhqmfsYlO0mhib10+2tNr149v8qtg8eK7
jfVL5hpmYfl+W05zcE07zrBSpqXd+1VUcu1EhSOnFlLor7rHzzVmwg/jTvAfApIpg6CtirtIUG+7
BGerWqMF5x6e8W8HJThBxX+h4anrI0CKl9EKNgUfCqhr+Bl53t9s9mWlaBPrp7ecR1hBlKd7qajV
eO9z5JKHVV81x8mqQVkGIE2Eww5P1VTTog7LUgi21D4IxlMPBLm79/cd9XGSUju9LJcYPx5QipHS
lGa2pkVBAG60be3BNjWiHUkUlqF2ZmwuR2Od/F3GrhpkbKScnTioCC+r4dX5OT9WpsFPDjLOekGk
2xme6/JGjENP3bU4rbAyI7CbDQtNFpIuB1hRrXLYfuS2TA8IiXhMg6tX21O7xepvAZEb16ELTxPp
s766A5ip5z8XBYztN3Wppx2pSbF2Kw0gPeDPaa57eUX5qGaMTpz8MIPkD6blAgOnGAE728FTz7Dc
TrFm+44jlLuBX0PMiA93swvtEYW3yGhs0jNfF8+YbHEIW9EEHbZF09l2jf5tUZIEfmrU6qTjcobm
vCU7gS5pby6m/DvtDAH2eEuffTJS/kew1NQxwoMTZq1CmBTiLMsZ58VRIYgRDy/7eaz0aSxStVgD
v8j+O+o+18xMty4HXUx57r/jTgn/xznobYhmrcz6FtzIcGQ0Mg7DwnQm9T0bpYfa6Ca1ZWhkv2BM
dPv+yua/L0+qkdd3K8RqVbaToVIDipd6c7MMHwLO7QiBbdTQQi8GOKwE9samU9TYM4jGh1YF06J7
petpI3+kSDsl3rofvFV9seH32gGryV1PEjjKkGPoD91spuTPFRg4nLt+J7YR2ptyMh1X72F79bso
+Unu10aAWeNqscor0GUXrj/GFtkbN438aFg9vLIfG82uUUWYXn+fxE2GhmKHOnQaB0dHyrUrewHk
3tjW5bmATZlAdK0UNUB77MKQG/Jk8T0CaJ+pBy1zSh2+md4r1QxEQOgWHigK6yMTfqnO/pVNaED1
lkjvo7VCQETdgE74QkRgNvKdQVgPMyc2s45O1FtYiE4a7DoGYu2eFzE2VcaExFvYduYqepH+tapi
hLwkCOAmKzusTITbAwEarOedibyfV2KSTQIWBRn5V3R/MkXgmxq6nyR7IM90iDWI7lVpr8QldoH0
1nDqDE4mies5irUmQofMmjNPXjGEcABKPLkRODBkOAmG0P8jcYqiDp5IcQk7ZgUA+DZ3BkLzkGR4
zJLLcw+1anrP508Sbh+rpN947Xyfl8LhFSnbiUmERIu6rm+ov9aeaO4qOe4qT8BMktwUuHpjolBp
9WKlJCUkZsvV2te/Y8VlpGsRuBN/Sk2dzX2t6awDWwfg238f34Jlm90Gvu5p6Eed2jOwnMB3EZMH
U3HEfQLVQejgX2tOS7C3G2LsVq5yICNvwl1RKGwT3ChHmI6fQ8cAFC2AaI9Cf6n3MekyX0kNnWxc
OxKz7C+/81JV778V4F7qACfZXccBJTdeYyxzYsx464iumOINCBzpf0BwVoebyeBl/fb3t4jXRfZm
wuovKQzGH5KZE9IrKvrrnCa45eT6BjkseA82diGZiqKM5XqGmBHtAkwnSWVJ+fA2dvH1N4XsNsn8
9ujsvjUT8MDXgvqs8vNyZBF8zfZwLwi1G8JqIE/KiSZ2NSg7lLEoEeE1c/8WTsbGunadj1DRCXyg
WLdI8lqiy2sBuBEyPmIMSPuuoC+2oasn76WYnXrSJQBTFAgwQvKvGMDEorVQ9fwaDNMlI0OFfdEz
HnZm/f7TKAxzu95L5BPCOMBOdm3+P4neckaS2o70Ridz+b3d/lT60P6RZ/D0Hb9dbeHNPZbiZtoX
gu3ZAySPBoggeW5dj7Hi5rz6FzYOx2rq+2Q5dHgHKPWCorJ22XMOGVKo/yshewLHjvy/wglPNIOX
PXBnt3OlUeSKIpheCQMuVjwnU+++/c9slvS9utvly/oD+JxlZ+Mm0Dp6pQz4P1itF/pwmGVweSOf
a84DMMPKKnaYgJUTxd5ZOeVB8BGZYuWTyarLhv0Wl/kHpxo4zgIlKl9eDjNETZ1u8QUTclWi+bdA
nlsww9FBuNVqDz7npnA6gQ9Y5omUf0r33NX41uKYWBQ74uEvRdEL3wCgcYmZhMbtdq8+woRuggUA
kiX7DZfJTxmQmx3dQGfIPMXHRgf3173VTTFl25szOulNTJw+UKh7pyUWUKWkZ6hX57mO8UGIhQ1N
iIDdpbhkNrujLwl1w7vGCoEtRgDKSxKxooe+/QzC6uwNa5G8ajrsMhVGMhBU6z1i+6kszNfuPmBO
4gWHO42ZeuJP5N9so2HZaiuaBgHJt5xJv4MNBw5+hP59dQpcygBSacu5+lclEjQVNafxMgFN2iT2
y48P5UMGN7akmp9GsENGCGLqxGBPc156g/OFM4m1daKYeWaFOrgqeHV348K3O2JA9JVGD/ZlyB2R
YKgGYgz9hX6YVUiBqVz1WfWBULRhJAV9uX0z569wbt8dKdiEaipLeCR4jKsW+Lz2m+QmSX+cXxaZ
g6ECskKC81Sj2RTY01P7vIrlqJtF3ksy0EtzEFFbawPU8OzXhfpIddb4qw5xx6/f5UIjlbPqNceT
yLNitywuxNXXQJzPc2KICT7Y6PrPkj2mQjuk3foUbBm97WI5LBXcrmiwKfUTNRlxZxyqqN5ztUhZ
eS3aK1d8J8iCuZLCOtSWeF5PvJ8gUEv+RokuT6h0UWyqjbpu3qMIMvX54mSVydmPXFpxGM7byX0n
gioFqySqfcdEpsxAb1ySv7WrCkguTMEpEQH3Xfnj3OS5dS+izkCNdYG91IdPzAkwyxIsMaZat3OP
+0r7xfuiAZfSKqOAE7dg0X/usdHmzhQh5+mXffZnIq3jYeghLrM0wcoJ7iG4zesbAetqo2Pp8nX0
K9DXqMLHS5jM5nAy9d/AsARYP2ofZT4N6gTJAUR5RyVbqorOv7b26yX5/K6cRJld6SstpygnZb/7
zljfP69Ylca4EzO28pqPZQ+ChAIDfIeXGjBB9zqx8bdllAxB6ecgt1lwFprshv83l6zLNpV5ye05
0c2mdC3LdyYcfwHPsrt4hBCp8XdZ32LQae5dt34wS3RmYUNbvDKJ2OwtIVM5jqoZle3GksBqGMRA
HGxL3bmNVez2x33SzMxf8+5VGjcjaHqdYzllBzmyGSTLoH5MTKvTOX6mvPIkeI+0Db3RnZzkTyA9
OYFUBrZRzTApLBNZwKY81soiQShlMD2SVFidlxjzcxNQiVBt9DJMv9PCuiOkFghEUBN65dBLm9Lj
a2uPQwzs6l/JPvCrmA7Iyb0CL/B+Wc5LMRaxkMO8BCGupp1CXHZYwPX2O9w5Mpb1EywVZko7JujS
GSLp8+LGOIP//5GXmFhYSPdD2ZGZzHqxIYZjBAd+M6hBUiNDCKkBMhTPneEOAu/+h3MPLmFf1eBD
/UmSxwr1utKASOxCVY7J3ft9dus7JVDrfLqZ/G15MZE3lJojjJb0+DxlWz+CIoFW1FbGXBG+dbqf
eJ20hJRClk6zIuffhxJxnUnoc6qSJW2YTnHcKpq0C/aLMMuYrFjk0c4oLQHN7dtwO2UoQikSqc/H
OgqW9MveSnHm0YMwXa3jyuet5I8ELXi2+M/oKU5Lza76uF2JHPjOwtAKZNdGjHLa+8AGmCZw2XdO
yvTAHz8m2HnG7MqMu86OAaCsHK9OrWmYucRkkLLi1GycnnZgrBHG2YY1Mcu8lc9x7FgcqOBV4Evr
oj9JdvsiC8RTxIHLCeY8+6ETr0C5k5ikDa/FwjDjZVyqVFlS3c/15cRgU88Xc21F4mKcb4RmK0ZZ
hBNKmlbM91WmLfxXTcM3v/6QNnsOWwovUpSyH291kzydOcYH8Y/106iRkRWDAetLZP9bBvPnnjy0
VR+f7FBy50bVT28iBNntOKfpo7STfau/oFBdqoXMMZ5/bOEZk7n/usILrGmM8XKczJtJNimFCvnS
JyxFBgvDyh+tfptMzEMTLg+sHZOjFcB3cUCgQT0Fzcjna1Aaa7NMSAc6Dw5XsEbVeCaTFHQ/1jpw
6av65mVDWSuu5ph13YTIV83S3DkXDOilMucqrgz2RYPoUY5GUxHjYqiOjKgGvYGc9KccMYUF/vOp
csErb9+05cvNUC6Jl/TaZrBMD5Qg4X7HZXnlsilGCLU4gOttpMRxXpzNF2vdAK2cb6C3eO6nCv/7
JJ11uK7feF9htZVGUT2nG7nMq4S5lyXAAq11KkHqym8XK74ngXkXP1XSocVc+Qs+XWxo0IDvrZHv
BMLfEhiTcBnyuoqYD+hWwIM3V3iA6NqrSWqRx3VO5LWr2YbMapyLCKvrm3fsvNdpDrS7lqvdb5fj
GWEpYOuf668x+5JQTKsW9Jyn0wBXBj438lNokrYSZ47i1AAt327rW7xyVfp9a4tK5wyfgX/Q0MCd
wkXbKZtDqsZv5Z0OZVSZ166XPJRIk2X6pVQE2zwHQ4u9PsTJXeTnIeKwhK3JkUFl3IAE6WDNDNHi
9jRHMjkgLDUAmJ0qXUvdYzOnCUpfmC8m849Sr8XCDfE5qawNPmbxWXEDkfeeDS6WzLkYAXBdK0S1
7mJmmJaslCW/hqzyTzE00E5HpI5XScjv8jko5jAj3c/wMG0GX9AVFGkibf+0SWaMVURYxwTqq30/
Cdke353pzN5alpMu6bAEv0AxQR+QYpfExrk5K8ENrZBLuhff2zOHpZ3638+RRYs6A42TpZ/AQKZD
OlygayvQXqVk8QtesayATVELrpoQ3s9nHGh83ib9ZNOxDqHKA5Bi1MaW20GDFAaeHq22ofTXaFqA
CX4IYr+JM2AnSikbffuvby3AQ4SokpH0ZuBKH5/wAQ9m+bSXd3cI4PA2VWphVtoMUT1n0HI8Pmvk
n+SGPA+sNT1TGLxNQxrYmsDFSo2ULh+hME9yWUYjLcyf5V193wbOW/jtBeWi/AJ8Toj4XxhMvDFd
2MV5oA8HQLQelN+SiXYIRgbVAT5Yd90Vst6vI89JqwhnQWqnz3tItzdbS4PPGyKnR4GyPxVbQ6hh
WkynZKQF5ow3HwNC1noiv+KGGqL/Ulh6h9k/FfjItIC7bTmXTUCsC+VZOEiIj/Ptxk4zDbKHkOyk
bh2Mon+oXQYIEdMHrAxPEgYa42CPjZOLBKd4oHQFbGuAlfPAJGa/+HHSZ6j9kSdBlaWI/qG4Hm6o
sMrD2Wj4vQOasRO1/VsGawGxYT8FHngHCqJFNXfopaeSFyVadzYmkQpBfRMvMzCYi49wgzQiHs4M
MTack1oYdNmQhZfLFkAmfFBTbSME/yic5jUMLXbUIZ6oY3x/3x5hT60yo8OgcoJJK/GkoP4uBFSm
UW5oJ9uWqQEkBAARBwvie/cJ3+KlNFzEtrh6yZm9nlPWPXNgTZQXBHRdjcJJ64/jT2wIZ7r7XR/W
7HCEpVmcERNMiecufb2IVaAqCONQUGVLiaPmfPlD/jEBF/juiD5p5mLvjGmkovQxAR3E52prM3TJ
uMBl8zH6JHmStZVEQbf+4XWeHosz8R0RDlo/fJXaVUy947pl6vNTHJd2aRl2acwjLJN3cgY/Nuxe
LgBs9T0RiBdZJf7vqCLfuotj7Lc/pTIEhd/sB3PrHmmB/8U00JmbxodZhXjLsjJ+OXZbqc+HnLoI
T7hxJrz6ZlD3p6hKMpt0NBFSJzkflcSDWKMuNRsGGi9BQ16saeqC0zHFzQXTmvBKvXtK+n9+B9aC
3B4iAW4xNvSg0szINMHzn8mB23K3q6k2Sfpn0zGVHD+yX+QGm6DRsUTe7J6LZ+sMMB2DdvseYxha
AFmByvrOdmmypyT0UJkE+bxVTIPOM7gevLcvjtX3lw623YiRoP7MLnNhN9Pk/v11I0hRUc+7Xw7m
mLszG5JSBCCTNB+mfNgavDFRFM3sIZzvpFs1v0TFULaro8A3ONhzEFJeDp/TEOdm8UkY9zc1eanJ
mujZc5L/upCSWhf9gIc6Ib0pVALuNEV9JPaRVjxG+jEBUSMmyhxRwn6yTLgp18CzMkm50GNG5oWM
7RyrIEfLIl4M/Ir5b2hfzB3An4waiXAiobmNLH1E21YsdMhWb4yY82lrqWJvzM9azkTBDVzDue8/
K91EDNckGtVQdxzR15ET6HE8TQb4mO2w8lOl7FJ+wYu/B08mrH/zz6yNxuvZVqTLXQbVfuvHvVA2
85kVGeaapKBRNP3thnIfCNomhRpamc/QK2bVFUr0VdHkXn64CbzjsMr5DE/rF9tM/cjttUVDHZ5P
aN7cC5a3NvYuyJoyWu+ih2GGAHRrYGz8vIg8c/Ez/BCVIlK2fzJrr6ezbIiwjoHsW2QEyCgHdyxP
scJcnfCBrjOry2kToTlxI7aB8VFhiUVmPjcXh44vHdpxX8TFiaiezOjIGW5AF4R+VsqujDaoM8UO
kK7XUqnH+YLaQoSEu4MuVG544u2CTjWBYyQpco4wK3hGAaKaveXgFK3Xhe6Cq8ZQd6QcwHVK1ANG
hXjXVbbWLckfru6zwstPu7+T4tl9MPBBqrJQcMXwLxb+M27I0Qz87SpFjnjL/HYqWt+vy+VZl0eQ
hLhAabRFgbEYffAskJ+KyMHpNwjIJ7y1KkDcjBZDOSAit/BRG99Csn9+TTaWvNfNAiM7x0DnPVD7
Nqc5prXS4rFZoreo4r6obzlpkSxkIWZSLA9MI+ZTdCRL+FFhPOBGBtCV51a1BEFRxPU1efT3iUX9
rlIUNd8Wv04QK9bmZocgMvFHiWPl4R4/8oRiRE94AO5nWMvR/HFBLWq3JdSz4O0cWNxbXp7ww6a5
icJro4ovLSeKSxvF5w77Z2sFHeLBhSJMMSdAMdgA3BX7BOSvHQgdgWv3gvAKLkDnP65+26xUpakE
UM/r+Ld057R9qplwUyCQP7XDcOdJgmzORI0/5FI7aHvrvSwLq1TgghQ7K3yekLJHImwnPOfDEl3E
zWrY30KLjwUwvCofI++3E1XYnEO8S3vJuK0uV9Rme/oH5S0KQ2bt1dWxksXtu1TmKFBMHPzR3WD5
i51zqZNGs6ocDgSZcV/k+VeQ+hpSFVjZ/4UJG75hUmSQS1+KXHYGbkOPCsGYhESOoTH+v6gFoAwZ
IM+4jMF5tMkFAU+Vf7/RHnFymzn6vb1cit2ORLixTA5Etp8BcOsEDgJYliB5uVOSknWrv+GDp+Sa
nHFl615ptFB5neDq/++I10YX3R3KZlb6r6KdC4QsC7E2qyZgdl+gETjEEOF5PZq2DiJtseWjw7qA
0MIhgOL+1gaNRPJclUoXsxFuqNFxFvj0xqaJxvqqU2ZmVhaSSjYFw3Zt4It1P4UuVFcpgzfOIE88
dAuzWrY0ELCSmpH48aBrpT/5FERnw+aKCZZufYKLhiw4BE4n2Yk28YSFz0xn+qr7O/Jf1I7EHQ+c
2R9ZyYWThlcBqY4HeuuQNAKH014bSVBWHAgq5b9yDv/+YW3a32Ee6KaS3XOzn8Zt2srGe2BbeyKg
U3a25gR3pn3KUliFAISFbv41aB1/Ged17agBkW+2q7ciZ8uAjRNbcebJLtFSdKWgECJZ4sODr/sZ
+mv/SBKoGixuxu3TZNoK9fpGhZrdBQXgYS0B7SW0E6Wv5NXMaefF2ODJAqAMUZBbzUStK9qwGg7E
OXxkD7Z3XY+IiFvuBH16d7bjsfzoH/Zlpfnu8hkSfE/wz/xyqJA09l8h9iEMX9vTTFV9rvKOryEG
NmF5EsD2Q5uIOjy6oHD6YfojOZXTPViwls7QTW2n9K6SLHuCEzwjs196t9KNuw8EWq6iDm81dErr
l6/UTt7n61RSyz7PNEkAdaq6jgpb1XjRj5hzMbDc1tXWuN52IVUa/2xFR7rPARRwH2NZihYKugRA
vH7VT2vzL5MtsdHcA2xABUHiJEUZjF+AOifS/jrzZyUCITAXb5YnFITdedAVx8TitBt7fwgkBNga
wSDZufHYt548mwGywyhFdNUvXuOmTOOLKuEBYTZabGAXhormmUUc+8MUZTBcoXp5ShFsw/uFfPtj
QnMYcNQ50pyvqXFKQNgyqmUK2ZaKIipG3HRMeRnFjy4n/jwdKPhd3AmA6In25TEXsuNsNWNLMExa
sW1NoQWorG0D4mLBnUTBrOyKBoiqrnj+bdlvy9sKA0GXY8TJDAkm6PhkntxWCSznJktvIV8dOuEb
LecAhskdUMpX80OjpcNvr4/4qlygsnmAYaAPHI2x5MgwJNA0M6amyEqRltPRunzO76Y78n1hC/DI
+RNuTRO+K7t7j52EG7+XjYxMgV6b5XYcF7gKBJFzyVoG4N8u38MbWrF98iDyc/TDpHkEA5ZtW7pH
mBM7RZMncCq5GUSmRPkMcYpM39mAa7qLsDtvSrdzLeEc8PpibaBFy2EJyJdfe+GSvnpRYAg5LOjg
VC2UsC+ocOM3RVLw81ASsRhvKvJqd73/y6pVaMtP9K9pT8KsSssZ7JkSIPTyLyegFH3Pav39pgKu
K6X4Qz0FW/qxChJ6Xv/F8urqZId0oYWsRLgjPsNjWTrTDzTMI4rlLQvlYlV7f+vFUy7vkGWrzd2Q
DDpk35cEHtdwhMB3ieRi6/9VvouB9luRQZeU6bwLPt5g7VMyc99HcPENeq/G+72p67F6x1AuB39m
M5z9RpRmyqek6MCM6KwW6oNceuF4uC7TCt9gUxTRZuDLxt7BTCn9jeLxYIHFCjtVP0YcPMgrA6q7
hSCNMXvvDJxpNAzHU947EVOn/X4Wsrn5jlU8A6zlueU6TU+V7XaXX1Z80LMLe/5sIqHIQk0fWHh8
6WRHawcKZFX1wMYnueg1a81Quoe3n7UbzfmE0UwvGk7fSuVuVTrrxUr6X7d3uwhqkeENbHDIoHli
iXQgdNpzqcZNQg9HkakM/YXYJrjD7S7p22ixv5IWS1RSi4gZG95hkWtk1BoWfNBBr251IOU8WXDn
TRWxr9WUWapWhyk5keImlGmKLZ5YGMZ2De4pqzUR679WqKR7hOU69DGkn1TK3q+2tlI7Bg9GNsbz
fy0/94DnBn6wAIJbCiXpVplGaReeb4oSUBs6GIG8oN/uakP9vy1vtVVR8Fp38i/r5NVceJGjJa+h
aiC/GdBZ6IPSkpBrWBFnmEI5/ZiIp83YwUQ70HZKLewf2tdiUgYJKfDhOzTyRIUOg+NsAbCOhaEf
M134uc+UE4pxv+XziZdUSBb1EI5Iml2MGHGCR4QVa0vbGUsBmHAz3PZ/S5MO8PQD7UH4acXxnPFU
BFe8UL0dmcmdOVgfFrDWYJrcSA8HyaDqgi3MSvmLz3UuW65KsP/+N5Di/4gP9cv2QExTJZ3Y3KcE
9osQlHo+n7oyeKvTiBoo2ps9JVF74yS/ByJBNUbh8mOGLtAzcstF8AFJw7MC3l27HdLO90wsdZ8J
rq1TB8jO1KYM7AF4ksE2hFjLwZL66CkeZKa06ALVzPPl7vEAJeg9jB1Q2pR2rnZ1wrPgQ2E+Jdzk
emJJ4pw4YYpaz0it9a/JW/rrIJC2EJh2lvfMeuWYQj89/sPykcwPrs8FUYcYsXZgfSFCGGbhDKwm
PjLH8JPR91g/oZDqiVOfdjgb0GfbXuVcSMf0GBEFs9cUcRpnHJMjj8whn/D2hPtvKjktx28Z8hv3
+0LG+r87lY9pxPDbNJyyXkquPjXy7m5a3aAhbvgrtRttWkvBfUqbvzX4zg2TqkmnsfJ3kbV1/jRp
PJS4oGUguWEkWu5Ve6KVdQM7A4qFUWwUhkJOlhxsxIVWWBs8z5zmGLjzLVaZDjKAkHTJ4d+Un3e/
nKSsxV8iTOaCGU+a9nmWDJOlE2DdQcePQx0BEJgq/X74TzKERP6exdZyrToVzaY3SZ5k8/HnN4oT
+YUyvkKblJqLt/GKTX/Ap7qGE/PlC42LkAvv3qg9VTvy651R3Mi7B1wFoO8aS8+sGePgooo9uE6t
6e0aIU9UxPN5QsctV8dyNmO7hJtRaV58QnfUgHDeCZtXe1J2W2T0ITBCANmHnfT9xtvvSII2Zq/+
24oga/UnkCPxqm6hFxrj/V7VZlVRvo43DSM6+heVDzJiPSGwodgmmrhCueIP6T3MqisROgIvIlWW
AHRvQ6ImbJg61vDmkLqpSVa8W1ZCOWndjNSiuHeLrqY3h/1hndcPfkJgnZnj5pqT5oB6gVg5S/E7
gVnOSij/IxGPqH/m+9/E11q3jIdUFVMkae8bxlT1amJHpMX/1VDIqBuOUv/ESTjgFGIiWMSAYu6S
YYOvaj1o/yWidDJStCX+FcqtRWKod44U45qY3/rzYcEMP6L4HVxa3d5rgPSUmAFqdv3igZXVllbM
NJ3VlrI/ZDWAP4M63uJbYxt0/mfV4Rxe1AuiBo22rqEx/A3HvDhULsjPdEax03D08rKdxVWP2sZJ
e7bd6tAbwlTsuOJzyxiWGfJIORSNdOcVzlV53jnV01jB8xKeYVfvH0epYl1ZDNXlLOBxZ8OjQ/ql
tA47nt+WIozWuJ73vQntY1RUmHQO6wAzayONHBibayH+91uJP8ojeoqPyKeSGB+7F+/p2guIK0vj
u8KuG3t4ohvZdst4d5vnVSafKvYYTe4cpzrWFm4uufwmQlMl/RbV/5Blvp3b0nnKru4TM95ROXRB
2Z5ICj6zckuzFlCEcCMivnXXfvREqMH56YmLzMczKZsTVjsmBQH4dfFjViSMzIXypRIEsV3P0u79
0XPZAwUtq4kkf3g2DhRblsulucSoHKOUUOg/cud4BYKVmQB0Mw53B8AlvDD7KEby2fEehNwC4oQx
3JthtY+vbs6a6hC3H7eRJ4MZav3a/TEkR6W1Fo57UwTopLQv0maOiv10jGGa8M0OOHNCl5QXMey+
MarZgQwqkNOKNoqKS6pacRsmIVtynt4GuE9R66R4u49Th7UX0EeBFBj2jpyuZHJpKl5D3GJ1FzqW
ZdubRSQl9hRuY7yAR6Q87i+EEYPEmAf8JSIzxTTgp+pxJJ4ZH7pzDt1HOWk7BZhrupkomaWROOa7
RnRVOTlq9Dg4pn0kaP984jwURpt2en0GY6bEc4uiGPYIDg5b6459fTyMAsCnXM3BGJQs2CSpih+Z
aQh7CNZbNrgW026qcXQGJfndcPyZ33nBmdBUeo5/OMvjNnWnG8qHPLv3UWiV7e/tn+ZQjZrSnWrF
RTbYU74Of3QjM0F3zIdAsMaiEghe2LZKbAKEnUDrfAow/QFRYXYDHsrg7Si5vo1dQqqcVpxUSCXt
XXlMggtB4VdDJQu/ZLnbGkhvdBPR9h0UeJhAdNVoWh/aqs3gJgV8nj7ilGSO6NWQspPHPcUCSJ3u
twQjSvAeZfQi5n9upZwbnhZMaxNEtWtqVvg6Ks5SgG/c5j3qyOHfrDg8kKR0ei9Kg7iUz59LZ15z
s5cj0Zr81JgPj+pcQrk+Vjid1VUmeQ3ZiatgYuOhKd7+vpRQXyRL6rRCKDUuxi8AdEWV8Y3BwyXI
fXctPn0iCZqnrL4ho9rF5R2n3Kb8kLUg6gYStpC2bVri6aoTKI0WHHI7eth4PL4EZT8/xFo/hZHU
KxqDNqRMedHjplHFUsXAP7BLzN/1actEBDw6pNEJF09nZuKcjeQeQeUj1R7AEML7hgorXsvvvFxF
lfCQUOBvsuVE0ZBUiZ62oaxL/4ek3A4/zYYaIBA+N8LmrwVDbcQtyoYSc+YNaoPLFtE/xZnGiv2H
yRlNAxs8qx7jrNhqPoPjmhOhBrKzU6CU1Tm2dr0gzwkZVMWNR19R5PxWY9qlUB59XE4F7XHrtlg0
XtDxg0sW+RB0/PKfl+5fcCAHg8w1dDrH4jMBXucDSfiWT3nwwwM4UAV7O8KYJmPNXMSYd6pssiOp
J5T1aL2nT/SXS1lvNGJ+jPGNbBK5F0uXiHJe1PSz74uLbJRsPJGhKXH/IspQjVL3n5+0inqZjFf2
xZ3q7LHVL657U4HNJZ3kvHcMcTlc+s2FP+b0iKHvwxHBUD8ZA5dGKnvKWtpmeYtYq+EJhwtF0ivc
Mtejxhgqi0E6h9EPM5Ct1DZaSF3wGtr1yX+VvuSmox8B3WdRmwB7tWmfvCXPgV2+QwCL7ZPgygUp
IHdm7LQlc0i7GbfsX7bxsfSV55o5rze49sY2jPV0xglvsdYjw8NYGnAO/194K+f3xx7LvS9xI1hg
TlYNQcmwYHY/fU3Vfr3j/qc+QlyhhzKzRW1dnwnis2lA2LPwbgSc0UCckju02HoEMB7sBsJ+F9PM
K7vUlEAkum+xGYGrxk8WCZHKqVYBpfUoAMct+2H7NXDLg4ba+aVjwvqxwyr2F82Ihon+F7W3elxa
6febRXWBOv9AZqyaLHDefPCFVP8VgUWPmtBD685rX2OjGTdlzb5aM4y0vR8fMyZIhfZYuRqvH401
GNt0cC7LJsvQsoyocPhlS5iDELhG2djX/14x1DjhgMQtf0I876wJWuJqHnucVniGFHYTDwIY12vN
G28rWN8DfhpHqvyqj4RK/q2gWfIImt7pIbyIH2l8GbSlhkM0mXRPkke7UcadtB1+Ttg4YCbUCvuO
ps09bl0XiPukLykI3rXO9TD3IKJyYdU1jTC44yRKedxc9yYCsV3RQ4SVtF6wT5ANNbLhPNoO9yWg
fYH1BmrWRVoBI/JMPWqD7hFs+eWXwsEIZn/NI7uJOtTOi/IslD5ey9yrCwIPXMKT7yRrA3yrIFFr
BCfplDt+lA+QKlqNGZeDDI0UtswHNu5ZPWxXgh+1OiQsF/nu6TPiI2j5Dbmde2S8JBC7tH7BtapU
exdKKDk88TqBtIEbdR/5nSsYIjzbJw65Aj+n2Kr+rmzraAsv3/uQd24DcU90zwmIa+DZIP6cguLz
P0tuXHlfAr7gOQrYNKX8ITWoFu9phu7fD3e0ID0r8Rlmwyyy3QNU9FHI0BCUNSDRYZxHi8zkoaip
HtXsxbbShj5hhQ6C9tqQiyIWwhhic8csQFYm7vINy2TOz+c5FK7a4hKEyqIIfuF25lr7gijcVg4p
TWT5eSMnaLIJQ1oxI56aqoe3avQ7jSVOl2O2CAyiU0VocnTHgmKAaeCTXBG/79gwp0o0IjAeri1J
1HdSiw10X4eBV+5f3ORPhRLjUAOvIHXCFYRKu6hoLlId3d3YOqQctzp+emzJzYAlZztAG2gooKo9
BxbSTQjI6aqVOxqP8zZqF7JgVSzFkGwgyNmi3OGuS74OcjBRtpcrwak9M3kOVpK0wPVsFHcDl8b5
5BsoC5zo5SjNzbnC5Lx1YD+H9PEoorcjlSrhtABs/BRRaVL2IPRNeVXkJ4WlPXGUsN6lqm9vb9HL
cIcOXs9Y7bWoSQ6czcVZJHkADDueqChb3syXcheeBl8aykUQgbP0+neTaOFPWF8n3ckphoWEnK8F
Duzj8pAljN7Hwjp1AiaT+xf2FcNA44MCC8pFXPEjU8PljIoy7Gz1BI7CRSudmO3IQz4yD3JYldc6
l/hGJvKDH8uA7zdsn9zgPp8BPHnI3cE2+hfZqvQ9TjJRbk2QDSiacPNZjwDFW6Z+3vwDS4xp+oVy
0AhJn2UlPNy31edTFwfEQ3r5oLc9SuR3f41StU/3xx/s/ockm7KyZtopKeXoGEhwQDNxQZyeynx/
g/tcyJuW3jfXv+hUFPIizgwv5Y/hsKciCapFSamMgTA+Jaa3lHyBM95XntecRRXTgNbOCpYVklre
IuJJW5iAwBq8QG69O2Uz5/jP/F6vv4YeHLWUMReThwKkqtUZtHIvAVjUXeBUQ8kjNhv1H3f/FIbr
YcNuLbLhLnRsPx23++/FBVXbaxx/6oSxJKWx6+psAratx9J0CEZIJzqfHmVmECmEPI70aKN2Evqk
o8jLx6mFeF6VZtJ1Apycd9UaVoIWV/i6pD/C83XRZ/XP0ZNm9E8c8gk+G+LlluXkBxbLaXR5y59T
2gK10qNn/NOIhujXAJJDar1/frB5gXmuich3/6Jbno+OE9QDfL0hRm31a00b+0jlpqGZU0+Vr1yp
5X2/ua6KmJz1U9dG/JlUboCD4g93g28+pFV0+Bs8l4x/GZ8171KFCormvQzbr0bQgIL2c7WuRll6
zGoFJ9BswkPrMwiSp7wf/iTPO3QvO5DgyYDgRXzyTbnW1cR+qMm3zUAMuH5gfHuy/3H2rqLLgpEM
vmJYTcIWuPINeveGkD37EJZ4Fjwo9qTcxBcxpRy1FOJO6lLtZyijwALFQTu6jyzcvapTXKSh/BhU
cW3FMlDwI1XAmKGpEp6XgdxC3/XA2hDEz94sFB714MJh5x7Dj2zcgDVIOhA1No1jESLQpPwrTIH0
RcYOYzydRJC86wp4+lUQjlfVdTKz9/8Qdg5WsbEt8jtDdasD7D0nOydZvi94ej+utNLbMNL7na02
btP1d1oiMBDzGC1VYlq5MpiYDIbioECyP8MRVtWNGeayaPSqqs/TJLYLTdJcRSno4CiI8TfzFrOD
jUN78g0z2WpBaGi7OVFe/AUPCnBZdwqrACQ15hJUqeVjksvOd/AqruaR835nb30c9ss20kk+M0ES
gufh7sALAycGloTRzMux55MSeqhN9NpZRtFq3pIRL9LA8kgVIuyWSGur1rWJCqiEZzfpPUdJtnem
e3NwpKrIpEPNlTcWHVMy6Fq0mr/Y7qfK6jD4O9URTs299MhxbW6kHc1AERhgKvEXP/waeGWgpoZv
ZbJ48ILPXxTgL1OZsolhCF0Yuk+97ulvhjpUn5zFIEW+qetn327hrZmhaSR/B2/HIrYIOjbTl+39
UluLYObmo0PFI8e9lHywDpCKw3uJtP2eMJhVwBPeVFTGr2htpCp2rImJ3J1KB1nR6VxB2jrp5JOH
zcSTHMYucR4mLg39AisEMZi1cSgNsJCp9d40cN43o/odXn/bC1g/NOD2TWQgCiE2SV8HZiu9SP/S
ZL7GIb3MBVeiJzZ7oOS7vztjZAVtZtWZFpbvRnIKad6JdfXq/O4zRB0VC8bJQsbYElArQnY4jg89
ZM8RailTH4pP5WcWBZqz0P9ESOL6k0/34oaNeK4DnbFxFyA249M/1MXhk/i6AMY9vsq0SZonHlVH
dLRDXiLT23VRJttCqiD1ALrpJ41HiEtjmdeZpFvwVghGsyOcO/5nViQ+LvI4IjY9qErKbZtWhnlA
u3YEWtHWEDMwUgfBqubNaoe9ENEtMevqzno2tFDqpVzlsnpasDbEOv8mBYSe9A/euMo9F1j3zwep
yz09dQexF/OOxu6UrA1VD/r055o7cqhwJdfMv6p0HNfPtDbyZimabJF7nwWeJX6T78OcwEJeSZzo
MRZiYm+41SFi/EH/uU+8BAhu4fR15IAyvSfnb8hF3T3ebfXm59Szu4foJeUB0qXxP7zxC02Q1FKe
aQQ94un91H+XYXmEoI08LGw+AHFkUV7L9t6irz4CtABPhlD8moGxGmd6pCylLvnhAzjzbsoup5Q3
M8T460P5I3EERdpM5JC7FEm0mSOu51DfAlUnoKwJUZq51dnk73q0aca2tzNzj03sNDzoXPpedtE3
aSrQxM5cjJUSF2rJfCjzjmFcWgp/vpDic0j6coGvJQnWY6cQpqyVMaixB+4Gt4kQsiIPSvt2I7e7
4c5qprpQJBsudijPpVTARv3rxGtDUNb/F2Swt8D7WgC1UmebDYzytB8ukY5Biz8WqZjxwlIG8Quo
wq9IDR6VOvW6zg8CYUBHqr/Tzl8RLCpwoapVzKfntB5x5RX5nQFvRqou7dFvvfw04shuFNlZWk8y
4ec9tP2bewz18EBm+4OTJpbTiWp85gWTbKj98laqbJnjGPTm3WcIoUI/9C90GdAX7lPFDYzdTdV7
GOVBCd4aK9e3QIMNj4fw+xZaw4NECG/3Kzw0yDIhP0fflEbMb9ja86Badv5QyztYrqesCfG1kvBM
opProvN5RsoUx7Gomi7DV/hzZGG/4TvMkvR2dbeRp2RWiZxz9MA00P23WLHDFYnULlHgI+7cwc9s
ekya1kaHFraAHHTXYeGEo9PuGf3W/ZoPHTKBuLbYdfjZ23ZC0pmwTcAJKaU6og6M0nGQSs1iDYwl
hllK6Fx/hwYVsxW/aBTnlxvEh9KFRqnpdJ8xiy9E3Tk/JDUAkhhGxcuFKeRMeyLLgdNl9cAvJ2Ay
OTQef+SoUbz7gMOYQZwG1+NzJYJhb6kEQb5Vji2atwwFZI3MD/gaaMTfDAqdAJ+RhYiFG6VmgORv
vNlzcq/v+VrF2M6OPlJHedTxNZxKtsPDCQBPNQbA/Bh91iTNfAr+TrGjd+kqL+90nRbK8SKnKvPN
DtAbHXXyY7sk+6knkyz6c3WtBNRYn98yOEVs65p5RZAGsl+Hh/YRmhoomUfLMN22CmDFHnp5+kbW
CpFx5meekEGhoUPCEj6G+g/dDs3+Fv4iaWz0fgQDfOvYlp2onYhQeWqQCfFf+kK0McRB+hhOrm3x
zvrtlSCa9MTRI1PkTkOEMGJoOzOJpdv/x18d1zbFQjFf2h3QjabHe+Qr2AMIvM4vIsgJ15vWzmV8
LqkRcn+C/vp25IvzYFsfUh+5vdTRx5mGkFPxyDx+dBnf6GpTh4n7Vh62O9x5wlEuzTHp0/0Twckl
XrMOe+weDy8JX0UHSJLCSXO7jWRz8s65f7yhKGNsvs//GVmV8v0xisnXzAoD12mp28V5wUcvBRQL
SmnOIwHj5K0NvIk89JZqLXGNFjJuUrXkFIQikG3nVnM7Twf2fThU8Hnru4A3r4D4fzVJVw5HJiEs
5Lm+Ap1zHEqMrTDgKTBabj7GzpJJ5FlGuF14IFDaMdYYKaE22M0Sqg84ehb8LAsIJb9cB9yWwPiJ
17VqYYB8ACubvEJrLp1kI9NP9tQlU1ztbWK6QU9Xy3jbod/XpskCmaA5yU4Bpeyhet69n/CdMcdD
Y2JUMIHCHYstGr7yous6Za3r3cKe1yG5EXtMU/zOuy0rNdT1VmrEGtFxGZt5dV3C2goOU+q4ap1r
zHu7/5iQ6oqXLwj7vZItVMR6h7uk1FZg/w/QILaxZ0PFPyaiEzvSx88V//5WZyBBqgqBLGEiCzW/
7puXiT8cCBtkD9CJ4MUBZBbIyC5zrRrGNNKEdIz/Q2v0pZZ71o4wvdBaZpzaGZIx0ODOM1b26Jyh
1NzRWr5zbpSnLbQ2UEbdvQ9VNT9A+wf7qAkePCrkE4HRf8NSbYPaxV7YpMDh6rUFjG098AeJ0nGz
GMRPbTf/bc/afxxuR/F+f1bTcsE04mJg5Eq/1CAj6/eGqgaTnpRpcpESqkC6tdpn06WNt3Opwk+x
JxCoFpTr0h/k8aYZPk4S/TecmmpbbeQIozbBrTe8weG6K4Ub9rL19r+4V9qrSZ+jZKrOcrtxffMG
kqNWPT4fidk7vu5l45e+nlr0fNLJXTfkkgSdxFxEANbnOf/GJSV+bSNEFn8XRvJ1GUYzJ1XVEc1M
j2KEc6rUqkzwgSViPgnXw0iOAHI4ZiRfFCaAXFFSMQvYuVEukepsMNwGbrTen1eDG1fCGRivK66W
l1u4w/my4gkoT87lLcFubd7EKHgPHatxIC+/LeDhQtnr/SL54SJ6hG/3zgTEkAoR17gUWbi2m6d6
IxGNg1V+Ko5LkJCA2YnEGyqD/EXeRL/luBOeFbCeZVpc8hvsrTXX5dEeg5z3F6UW/rAnN1SfSKpf
GIwKZy8+kZrkyWpkGEQVzOvXxhWb/PtnZ85cx5ohl46tfTZcNnFqMoZSbfkaJNqwSzrspVcbLtSq
yX3eK1Nmv5PgrQQZs2l/H3JHtkxcrO3Ln7Ug79/UBxUFOEdW15CJhDHgdx+GjuhJgd3Hrok8Q30c
VYmnuY2sYcmZYROFGXcVcN11Dm2SAgDSgwkdWAeDm8PGO3jdBd8CDcaR82n6RXN0GwNWWHE5mbNA
RXolApig5odcmTQm7eda1wCMc/u+cxgbp0iHhcVsCk5kD0cmr8su08iQPEfL/sxaEMreva6AQk7/
PhA3ZvLzTSBGoPhqJ0UzdfeOuEqP+Npop33I2mE2kzWhlvY0WiOgqePet9D3FM5L6YOUkNlt0YgA
1nTFXZQm0t9gL5xfnHqDYF3iFAGExx0LWkwOp3nAkejVWWD6qnPiUi2lteEbT/JtLA7On9s1NL0u
xYKeXIZZxcuJmVuoqhvd2aralGIozPxNAdJKpfmz51XFR3J+7lmAR+twMhS3GaN6LGF0LLgeV1Fh
hYLUd9Sj4ds9phbrrTOHroZvbYZzt9M+YTiC2xGdeamUPXN7RzGLCjkObOSHtW0Z9yLtM5++KPCg
efEkAwGd3Wqu8aTraJ2+rhBY/2mZPQFfAlCaLk2gJhpdDTazMygjgUPES3SUTLS3uSTUjLNwy4UH
ZN4N6czMNMjPQHjTf0H05y2lYPOOt9hjX9YmgsaIH2Y3GsnIUWhU+7Pf+7Cvd2x1zqhh1DZRk3Zc
URlE59DhNsowDFR8F9vN3+nLPFRIPsE4+lhm/1jsBNex+65Nh4t9sswBUgHlBLpX5tWvAmG/hr1M
R/LUSCw24n2IrJVMMccRWKhF+nZ4TajwrG6VVSf1PcfZGob2fByDwhYV5l8ktRpNZpZ6mg6rNu/A
AkO040WW24iGLhOlzy7Yty4F6ZwVAx2kmh2yDRGn+N79XPbDGQnwFTIMax35zJgT81iBaXomv7fD
XU/1i6n/PrDt1SaEutnVogbfsorrJCLvH276zKNB4NKSD9z5Gm9rAotRY6hOZZuAe88/SKvxmZVG
/P2N3eKDkl1n3N6zEjpKAq6wbo3hrl0oIaMre8vKB8aA3whcHoZo46JjFtJPAOBjF/ljvU7H3asd
EH71zke9pKcm5cL9fVuQvj5GKvxLlWlPm0ABmWw5AG/cCqWjjnmVxGiPWCb6MfXDEcAgpXK/JsQb
GMEhezqwrYIxnNJOqEqgm6AGUOSib5O87a6d/ciMHPg4AbW6GPsuqRyDmwATsV/Cw0ryoQOgUOdR
GqWWwAdYVgwCAS7PcWDe5qXAazip474SUku/6ie5uqhmg40Z4Zn8P1ujzLvObtu1Qk73ztOAS3Mk
g+23aYmhNfp2kQ5TzJuGGCTqs1CaDq2WiMV15BkQceH/yqF0LNgIORW3xWYY5zvbs8GUiWXppJ0y
nw6n8p8sYVcdRof/Vab+wksgIf42j30dCPS98s6B7B3pDXqKtQdeVuYu4CpgkqNzopnYQDH8atMl
OlbaMR2GK9VEqvfRjWnnY4odqK6k1Ii04biqMyg4ykiDL80YhO5ozISgWP+uR0B0dal6U+kG6INy
5ZQSRbck4seQ79U7l7sZ/klVGjVOJJpz95xcyGfw/U8ESHvsKQEeX2bK5DkYiQuvmoQOkVeytF6k
20IzyOCbUMO3woJXM2F+SjrT9TNu00mdrxDKr1nBAwlB72LRmKRSrajCnhhhS/XgMybd62WQLbn1
90FwVEoO8hTlkBpDgXP5sVgREDU2o1K1gvPZu4xmoIiGMpZbK3rf6Mjs2QZ16zih+jHaAuY1iDrD
8e7rX5y4WHYBFTLPla5nhSaqoEg5YfhV9c6h1zxOnF3XSxCPdYuiR4NoRQ2rUw12jI6TluZc8uhz
isfYP2HF5HLBpLfIJd5wEjwm7ycZ6vU5wnQMUsaFRCFA3oxdIWNAMZUcpVmiS8PzxSSah06ynrCS
WsrFlw8j2UofQuBmU/GmChYuj2TnsuFUY+oeTm2unW1/HWK1RfIqtfHOK/Lo6mclpDFCjAU+HFuD
IpRfqzgp4MyuvCDToIOa02fZDQw6lbQba/mGLbhfr8FNyt2nGBVyI/YovSo9hYa4+zBTdDjQ2sXT
SuuNPthJePgnxOKFNvxvkTa2uLubSnSaeugdsy8OwVdOkDgKLIr4CcE8d6Kf5LRdVfstZ1++YUuM
3kcZ5WaXR4ni3cmCLTUtSwk/RQ17G0T6MyfhOML3GskBvyvqkYan386OHsL/1+/3Ttw2KhTn5WRF
wXvtHIuzKSzTCPKkTYqKIzUsttU5FpBZypsFtxkIvLMDXshA6s5/qV9LFKIVmTYHjrMvECB9EprQ
eBOFQEE9XaRtGMJuq/uAni67I1B9AfFQBlAr0dcesIFPHpJG8uVlwvsjyOl3Q5R4xcT7/hOfQ3vn
IzM8613q1EQ3GdiJnUAVEl3KnF0mH36+dD0G4TpLY2OXbjAF4/QHsHTvkrfUZfjDPBqKUQLIxMRX
1IzckgJc1THiiPd8EV5aztujft8GSdP7BVD+WUDFdU5dD4BxC8GpoBasH0jyJ0nYTiVnEx0gYb45
UGokNNAPyrbMT/r/D08Fxe+LEjKigJRAqWs+B9BiSlthf3yI5cgD5ubnuMCXZUKJwQ0vQXWwJZic
iOJf1RbvQpE1vby6Cwv3YC+nkpdw17A1RSyLaMK9RxIXDOt3T9CNzJ3a9A/zh1dcGWi4Sr5IZRgl
+bsImjZVad3kAsrGFy/HZ8Tv6zAW8asLxMJBCuVo6T/BjskQcnfhsMZHr8k5HuCPCEoFyn/zOJCJ
LgDTMvbUpZ5DIifz39vkaq8TttN/EmjY+u/at7vl4PtqHqhJ8WXwqH3nRKhzlIgyZwdIT03lbqxq
mZLrdKhF/AKlcbPJiVxOIB88wz1z3gZyxZ6aGaornHlu6tlmDG3hz5bL8qitNPRqBIi0MQhusD5b
HNcseg5aQn0p82jtoZ70YUOogcetYdx4jYwak1UUcxLPcDZd1j/B+It4/YvmNRPUqhJ3Y8yXvozZ
9WkkfLoQCB84p73+G4fz23VwvR69aPMXLMWUmqkueFyr+aj1bhwk/sGJd3eykWyEX3456Le/HFiF
NDXBoDx1GJkw7Xvy+WOEz3kkALgDxAvCx1Q1Vbw1VUddIhT7rXf7EutUxdWmSFgTOWZHvfgE2NpK
L8GrrapPSfDnKD3pyY2DLgiVNpvXOCIJdxWat4ITeYbPqy0yU7/pl16uU4XmYfAxk2i4ljTDTRH5
5MmGl9wH+xpBP5okPnaCSbZjXpwVb/qXAHJRnR0lGKHqPQ+wbOeNnEJi9jidbcf7eiY36uNHrfD9
77m5gWt3oO2/9KLSqucDnV1VsPkeWPfdk5cpmfI/dWny7dP+r5Br1blkKqJevYOwPUYHGEjYkyaq
rJvMtisEqMYrLs+iag9C2eGC9daRZdkjpcpxK4xetLLdXw8qXGc3pcd36j06XqqA3iWJ3CfeD7TW
v/gfmUrzNzjQi17GxePdrX3RxRm6L+HcI88ApjIul32KgCNIoZay5OfatrpyNbYG53ZCXQn7p4Rg
2UVpuJdTMpANycIotJQZVzbIv5DjbLHFvJr68MBy7zWkLBKeog+nOCvoV2F4Dn5Vnw51bRXPlTul
wCd0hNVWMo4mzXfh5RhYMaU3QWJk98qnUSCo2DPKcLnkKfSs4uiwhK5YwVVxI+1cbwVXScmQWh3Y
+llt39dinCG8SGBKt7UUncc1dwpOJGeHvVp5kGeJpFRD7ziW+sS+yrcSQLthqIIydOE/odS21wCk
ciFBo850DYR00MbZR3Y6JQM31pV49qdHCeIhtN9OgSpASrPmxf7NRgyTDE3IPRgBfBuTaOgn5Ku6
oqvH538RFzxucHswZNLdYvMcTCOQ1LorHY1Yc5MxQbkQAByAJhxYaIFfLX8Zw8AI9prhZBZ8gqYM
wDK/3R5lTAtm0CgPD/cGZ3grAZLfWnuGgvb/K8V6s7hwiRys1eo8s9Sni5f4RVvfHfAmHJMh8YPu
/FU4o0OV/qsXZRg0toQ8lYeU3+736BZpwyWKk6eIRUYJWU+5XzJHTVh9HcJI9GXcSHetuUIymbdE
GuRNG9poOxT5PMEjPG6e68shBDReamhh8z0oaBXvnlXdTJsimzZrnERe1Ba+sI3j9xEaf2nUjpwj
lhbr9BA1/d23IZpjKQo/0oXuGrYubqsYjyW92RpiifglR0eab6R5u0g9WBiSequ0jhArm8bI6GbL
WGuz6qQp78/zsWLrieRmE0/mH2LtQCVjLDP5EPx2VvrMtatgMJOEt980MZnB8maM9hOInCqjROyW
pq2ssLJEHT3zc5nV79jPvNJet90ORJkv27COcJXGPHZ1myXCGtdzUMHiI/37GUBiVychHPbgQBkF
wxMmssGYe4/EYX12b8ODZSyQv2F3E2aDWzPzqeQFm4j9f2croj28fyvheAddYowO+xqnmgzRwtdA
+jGwUPNEMRIhshLiG3tIBzv43XT6CKE4rwqLQ31csC5eokV7Bk7rIKcO+7GF2WaYWnaebrQByBg/
efmas5WIMt0z14n/USfZynLNJbGuLBP8uK4nVl644QKuDW3xvX2rjChU2IWBCVPz6/91jOIfJWdf
GlATUvs6nAGav8x5bjkZls+iyEaJ3G1DS+XJ+K9IWy55d6km9s9VujzlNbVE9c5oFk66E0+tgdob
NYeZsUt6z57wYvxiHxaIX09zKgYGpeu7SqNWK57IGtRQYKMnUs/KLPxGdnMUqtDST/TdsveBivi9
8j7wgBbWrEFD/OcXXh5VSuXCN8k1q+/zreQMBUvTfo8PTARKHvN7lVRQ+i7lpcx7l+CzK09ibleH
1VdwFffip/3dStWHZj2UDs5M8v99j5MNjRe0401JYry6Ny6REOvVbfbIZl4nWiTTxDX9M4ZDKDix
pcVI1oPJAo0CHgUedj/kPLVBoUfozZhMLc0XIuJGM09KXqltEqkvzYHl5FuVqrxkh/h4Z+MGuCIp
Bhrq2GYPACM82D9wqcQElXpitMlJACOgZpMB8BsEbxQZqysl2kc9u11P42lzvauu5hte8+psAibc
gw4O2P0KDg5Sz8TOqy3LYZNX5HXGKJYNVh6Il5FVRhkNPlUqkseCYaACHBgIXYPYzeNIR3vVC172
uOHHzPsN94LWhd+8KvlnTnuSB0pv4tmYt1ixk5gFHGP6r5tJCOZJNLWG3RIxyZiATfCdUq8cgjx5
a1IyNT60ntLHMXU0vaCf1DjLNFww6JxuOO399fUyh7l0BusAhADmqllC5AsKEN+FKcOKl7wGCzh1
0/7R2DkH8lDavrxoreKfRjwKh/9Sn19cLQ17rmd9yYkLJ9rUfqGdknX8HpuZgiz7UB9cSy9jFXuu
3yjrPewe+JpgshgC1pySEic3VIjRSVLUfxywUyJOVJ5l3ZNLLcL6u04glG2uK8ppe76TDtZcK4dP
luf+Ar14oO4nE1mxEuBwECqQOYL+rvjqpznNPSuBIwe8xL/mEek3dQkakIRfD/dLPECTi1nmXC/d
zkRinpsIIpIk/tpLO1QlaCohkrEbcx/sD4nQj8fFyY8+NMctiHkH7DzMJydFam3BVXIt7hq/ECXj
T68c6MAQ78Sjr4KeKJvNKOKjqnGt2QZXk0HkZ02kQlnqe5ECN9+l23BVaqhNvB6NX8LJY1TRoy9o
uxZ5KGrdR5+w3wBiQU28ZqxbVNvU7J7O0m7/H3MPjPm6e2wHOQuA0r6Hz6cErUd5EcWgeW/lT6BS
ot0efaIjdBqydLg1AWMo9lgoe0rT34q8BxKxVLws2wA2HRVZEEwpLczRqs2DJyR5X/yCcR/yzu4j
2mvOMov1VLuH+F4Z0Ws0gl6LIMH7mXFTNt8NMqO+oG4tfCjT4oEQlRGMqFw3tFNjcVg9WvSXmJMm
oK1oll5W4KUuZa2HW07w2QxJSIgpA1HbVI+QBpzLMCR01gm4+reJ1oAie9cHjCWaGPRoVy6HVVXf
KRDWwgkuZSPIOpiCDsbQeC1Dmc0pS+qJZkfOWpo3a/qXrP34ZJgMzq4seqhDuuzMeAR+boybQbWX
w58YBq87W8KZwCCbBJJtWCrJkAI8xcIpzPZ2oG7THoYjoBSdHpr7fhz5jChdbXm8RUK+FNaEtheu
VqjpCD7z3DfiA9dHLvTLPd6Nx3wkybtI0vRJDF/pB53EbfePzU9fwN+Xepm8tfk/7ncOzJB3APKg
PorkTR/g+/mxPi0A5Sy5yqqesC3LmWzQTeD3TDGVEQrrTBb/hnz8y3vn6y8uwDRYZW016Gel1uCD
dXeIB/HEWkq3jjZZFEq2xjnp6HVHBNliQ9TANGWu2IjfGl2dakzkpjjV9i/f8OGxMEcRfyJQSNcB
1wS/hwr2RPCpsXE+SqvGMtTlWJFKEr77Z/AYz9TF0Ljux+9L4XBjQ9hrpMBkXnRpCiuMqOk8dNZE
c0MQDgAjLQGSXVLkl1aaVAHCImbmHoPp+Oy+m7Cj0GdQntwlDRCkwOUYN+FDf8yAr36zswpF1YEs
/MBto6e02ZKUXi/Mg/4Uiqvod9j0oWYziPMP2v/lI+9c2bKni9GxvhP525McU41VKEiLGWvwwJFN
EDHp8/YSfB/S1G6MDfw/TmVAVo6C7wmILRL5FlJhG6hBpjPqtHfT+yYVn4N138nKXaicFPmQyZqH
AMsM+uwn0xtDKFp6UC64at1hFU9uUQhqU+KMes14D0eOxJPQyeUkG41drwFKK3ujBlxT4wQjPv39
jacRWy1xuhUUOuR9lMdk0t9eQp4t67NQdcl+vEl95XMoDmFCwY+vPp4TW2VIxG0i+LvbVXk36+Yv
fHYSyJHPiLw8lC3aVfEOF7ceqFEjvHrwK4JtGeYJB1Lj0UnGh6QNpydB0bfoaotGeqd0OGziVgI/
f8A5fheIZcqshnJrp/ZXucAJYgkw+1Iy6vQn0oV8rxEBa4wBbHARMzJ43XuHKcj94Yp8xsw4jMZ4
6FsOUkUyLGOwagd7w4daKEuXx9RWSzs+UDMM0m5VglWsrIUg6oJFvpZ+UnMEmbQZAmLlGigsNoPF
rzfsxfH24lunUDG09PEsocfoV1bruACnyw+kec8uHoBtNwzaGlmKMor6kCFru4pmbyBwmH8fpv6f
/6vQnOHqFPR1wNlAKgle/VYNxgaKjdjG1pU0Iw+D1Z82cHJYZ2Lg8s8zc0ZVJ3MJIMcasKFlONdn
TLDWGahZX5pG/u8cFEMGQ3E2KY/x+ShjhR7iiGu24X9z1U/Cd4Dy0EtmX59nU7rD7bJr+mqtTqHS
CfqakvQcnLn9Xe+160x2HHW6yyMNvSf53UEaeCUSipJIidoBLKH/eAAR2YXu/dg9TaupVcx/Frh0
ifWlhMixHa3kuvoT5TPcaEjM4hWY+8+Zre+6ELH/EVNyViDmc74iwxNDe+ObzjrWSBmnfHjFXKz8
44ZO8pk62z8byXd0aiNaeuclmbQ/OJwM86w/UkmpC5qrRAVtkkerSyqBzcZm/bTGlgWKZLtpjZ7u
4Sm5h/ImYmOPfaJ5PjOPUo5VHAUqyiYRfWU6C1nLcQeua0yM9MaYnsgUIXrCGtlbVBRW2fR4lQy/
IfIt0nESdHiXborZB0LGj8sgnYLmwvVwRd0zLII5TrX2wv1po9TON9Qqk9qrUHslpKPCpOxnziwY
NnxkN1HMqjIw5q+68ogp4IFUGQDpMXu9kihp2o97+ApqDNqD5vaiDB5YOemKiv10WCFVr2YFhmgs
s/KHXZw58/8FqFLRDQBN2Ohf4MW4Z1IF0dn5ugomuSxB+kzlhXkzeCHKIrbJOEDGetH07QCqd1z4
Z9gXHMOx7QbMLLLgkJLN+MBG6a0I4kKEDhezIXBMTc1QDQcPIw7c2g3vhP01Li8Gj6BsQXhWoltU
2nWaB/cEhmGy1nTvuv9T0v/5q/iKHsNkPlJQ+kwKgewZbED2A1Mo8Uzm2eSRZFA4Rr8Snq4Eav7U
zW2njLvQacEG+jvPQ0xdLKO5w+6vpDgqOLKa78OfaffvE4h5iBJhlHfVgl506DiezXzOJYUE411H
yy+QzDBnxm37RZ0CCVRa6eFHNNcN5n+Me0r/NwF5M4P9qvCGwSfy2Phdt9SWJK1UUHYVeBkBNS3c
MnUJRcYN6OShxTff1Dh+FHEYwXpseaPPlXqzgXtfm1skia/vyYx8RgfY4iaHrCIaCOXG0nqSTf1t
lecpm8fRo2s1rAUKkS3QG8bHhOa3de4CLkTMnJZwXuxuJgYxUdQJjSfxySfmW9xQseegHz6aAYWz
1tUhSDn2YzLF0WVyyZ6nDACck/fmAm3W5hvoWaldvUq/5s0iITuQ5lsssyX9359Nz6SlaGSOVX20
GZ33cSY/lj+v1UNMjkzCiQ6JF1GUgchGE+QU8mhBEoxn3jZW35v49xrFniHWC+fTY8DRtX8V4SqX
Wlxp+H2e/HZBi9oL7yAuxVqOMc9lp18e6KLf+MTBdspMqvq2a22JNslDNtTCkeVtcFpYF6v9bc+z
yOBxHu929pteVYiVxPsnp48Rvpi16vRuFmsW3enatu+UG6QHStckozcFxD5E1QSthLbDvAo4a7ER
CWf1QJOM8Hm0+yeG53xmZQHNoI+oOfp7lleQrPqgL590E5I2th6UZsQ5S9xh3FSO6e5qaKNIf2Oo
wgm/g4KERExrb2nIB81LVN7a+TAhwGIzicvex8qzsRCDR7esJ4FtN/m1phPW8kPc/ojR+fpD8I89
C1tiFCDPtWT3rK2Cw2kYa72yP0aKvUpG4zmAtZszHwUFCt02Nt9RRgiNo4Av4X5MKe9SO5/VVRyR
YNfNqyNR78jLwnGdj9weNtZW9/1CsarKec3dPbDvnE0BWngxVxR+H8LfWNLoEoF3ghQnEWRbBayE
5Xg0BRzZVk6tTDYX89kogNbl9VIaRQK5SU9CRSUddqjSVV/DWlm4v9Iwdo+WpjemQBDmn9sgSNIB
Df0JPWgoyfgamO7kxYL0SQfBK/fD2oIeGVke+ZKr9wKeM3zZ4dCIH2l2D4OgZg2bTFaTeMVU+/z6
5/0USGyMsvhMJWAwr5/NF5/w+ti9/49GVxJDnwhGAEi2Av9N/D5eeIMIwoKSy0ot+OhnpBsg5Qp/
mMB+TuhwFrXKAmP8YrA+CsYXyLz8BTbYfXNaCyxVhUvqfeDYq7fQx7PTAIDR5LODbbuZgybqNVpG
l373c78gKDBrTFfD8KVxbsCBqc4oaDCz2Ihq9S2SE19M4OodowEu2IjTmNTLBuRhGBYoqwj72pAv
V619SJtXsfuvMSA+Ds/i0hHBY3O9RfZzYZDcBs60+cq/JUABFAS6nBdHHDBLLO7+mpFTxf7iodF1
qRVu41QYdL3JLdyRCqOmUwEF3RSbmFfFEKfpGkD9n3jKl81AWRZOqZ3nlG1cZyTHUP32IJGL8rZc
NNEnFS9gUifL46EIqQKhs25b67sS/Tv3icLEGLGCiuoqx8cAvA3c10KkgsWy+osdvBLHXa0bquCp
woxvQQT8z/kzPTUKwyxtfs3wvz/8+zzs3GTwCED9p5PIj26XjRuEjay9AvoLpOiaImQ1h5BBACMv
YuKd9bnl/dhl2I2dwxgXwqzzqN0gghyM31tXvYmBXZMABBY5uiVAMZMq8wCp4ayJrNCfuqHC1aCG
rJ5FYStrYuSBYBJWJDnBXGxg5qhMDQ9ssjiYSp0EfqLEVkNeeaJ5aNZx0F88WqBiNXZNPMPvQ5Vq
oMkzo92jDDzLL0ye4Tbhz2y4uu8yQ/xijd9k5+bm1nTBUwX1K3/dB4cYl4xr/R+W6x8srHnkqcSw
zI/taMnZwEqcZeE680Y49YoOhVbMGorgMcla7wJgkuTgkJP9Fx/lO4p1+e5NM0LfgQzM0UAkvuge
C5w7a7DT6byPT0FpoBcPadr+9mGDJFxZ16WVNj1bz5Xg8B9hwtpyjV3La/MTM71QcqCSv+igtQwZ
v/FsFBerIu3Ia24RNVqJRbudpF3UC8KaAuD+Dg/12rT6f8fbEX9k3L3S7TuUC5EGQpQQ0roXMB3x
jNjlJg2sOltlfMnUq5HuCuJkxtMz/Fwaa2OvAUeKjXy31s9wJJSjel+sW6xaxgDd0CIPr61m/Ux7
QcRInYfWf0E+ROAqmBsFQr5u1XWgCjsZXaX2IN/S3FHac2dc1EOJKYmqQtIk9ZaBI+k8vnwNLtZf
RQJgMXeEUMfwfGjmmYgwPZJlJoYhNJKsEtwMe2/iPGYffJtnew57HM7vuVQ+loCCiMnyiDh5ozoX
Tpoo+bGQX20QSL6vj9F7Q8gB4GBhw9hWiPzO0iEB0btL3uTrCA3EakshuuCewBa26Dh3olAm8cok
XdAhhY81d6TBbu6hoJLwrXiakbJZG5QV344Z70LpVJGOEBHO2jJnvUXtCrSddPplJpzAVPPL4i1k
+MjBJty25srO2Jssn6MAitjRTFHm3Ext17YUrkJlkCQUr321cE36MPRHeOroizpCzLDeouFXzJCc
nUuE4yj5TvlldixtY1rPb6lh7LZzQ5fjNn3wUq5IQC20JP+58OobkTA1z0WWIb1SC0A0cXbMtZdR
kKY47oj26mIoT/B4HxQ4ge+VkJcTNPh9k+h32Jh5QNQgsA1jue2QRT9jdWiENpbyaoLRBWHcEh0m
5L5r1kYTBffuKJH1FQ6X0h82t1Kk2vE0YZTzR80uQco1daT0EfeXfFb+RkYlcnp71+UjX+/fXUfY
mrkf9tbqm3yTOJSJznO7VBBTcJpU3LCYmmfcuidn5jtvuyEyNzQySdB0e6pRyqX7MsoR1+yk2IyG
ykRGnDI2AigE4WyLa02ID55V4PRVg7nY3OPndpKjKDLxt3xytBI9F03P+xfwBKCPmf43DnoQ0kOV
u/dKp7qOb758E00qizabHGZKLEp6/97LyMTn0iaYU4tx7EFgnZnNDjE3mJyRLSgKNqJbnDmPGWcA
Vx4BoHNHp7r5WLjMOPixiO9Og5DHE8ncByaCteuLtj8Kqimp9ANjwnw61c1NRT0JWkzZo6TBO/0l
OmZyILn4QHRzQ2i5UVk1F1O5sehtE9JLe+OJpDwLFiKe7IW5iVa0ZN4x8GA8duG2bZ+EEtOcrqWO
zS/8NwTVvKcdgwZOhnG7HQfDT2xMbXM33LSWTS8c6yZ1WEqeo6tNiiczHvb/2NW6yN86ovTaFFkZ
zHBGOhrPYYQSo6D/GmkUnXa/L01GmQq7lfdjUknLGAkhEAs60VxP55rssf9gEYTnIqo2myHb2tMV
PxX3UeiupEIFQnR+E5a+h4qMT2oHn+rAkIa0ZBL+j7Hxc7FX/z1NLpa+BVz2FEhJKOX8Ue7w2+F+
TUpzkUifghzSwp74rFsAE7gkVbfT2tccpb4CvY/MQPLAcc+eJHXG0/BImm0kWFJFqf1s0wJKNYqD
C40mWbv93MaC1MH4M6TAB+GebZ64cM2tbRQtFi15Au/nLYT9yN1COvi5s8T5NzHrUqbKHeFDPqP9
b83LU7Lwr+lWTKoRpSHuwm833SjXyClZitePC/8nTY1XD0NNTE0Y39j47bDEeYY6OAk8ucMJpeUY
8+meqrAPDfkyYwsWi/e9UZXC8lq/TsMx9zUc7cAPfj+znHdbf4QS9JU9lP4OjKmm2Deiaw9sjfHH
6aKwQSM+oipaVFAcmjDkPRGXQnChde4LX6/wJ7/BtwVgVcos/2PgSo4hgUvLa/ClRkxsT/3j5gMH
A0oKanc7P3Nz6Y4GVM0Jg4wpTeBK/tp5YtCimzoZ9WDozSTYKhGDeMjgT+Ur7Fw0fNIJnafyiG+0
CX/DQ17vBOXvc14ipfzYLZLUYgpI6DrSUVYiEnHnRefhFtcADGgRG3AMd+yZOYWuD5OLtbAnAgkZ
eBkA4PWUjSW7q5UZg3wQfvSZif67Jtj6BAEESMnQAs/NuOoUo2puSfjnOL9ojCY2LVFkMIBKg88L
YQtKXDTbG6yZ5P6wnPLCRJYgKIpRUAmakWz9fhcDLulLSIU4u8EQZ6ehjZeSLQq8c12oXn9TOmj6
G5F8v89xAKqbRYWTgvmrtGdkLva906pzJXbcBxHnqMXFzu/7CSxUkWm/KtQrgE0wrIXrKCFOJI2p
OV9NnKk1oWzKbttoyzgfqnIed+3y9ii9w4P6RKFgIeqQ66tE8qSrH8WOcKNAgXEzP1xhXL0sfh8s
LWPP7U/OoSh1zSHBsNg4OLHyXGwHSsf7rMvsXjKxmn3Do15utH0wlBq9ORIpLN/XMGQSRACj0HYy
FijmFA31hSkRrOxFBL+Edd5SyvYbjMogHQOdRljvZHyEX8y+JY261zNf4Xue3PLdMwsKhEURmbq/
MLBWPb1qaBqzmTZe6ngv+FAKeHBGkR/QPcSOOpyYdWJJga2zwyUpRlFqisePqrWcBRB2C1ma3OJm
w4NRbfVIO4YiJQrCx9pAs/pTA0CVy8nRl7/EXnJQVOa/pqsAKNuEAtKfujcxRWziUGsdYEJqvsYL
nS/kcJpe+bW6myCxCuoHncrthRaY6BgDyYOevEtCKTsbiaKI8rneuC+l3O/EBXGgC3JR6UW4KgSF
icStE1/p3zHz+buMsv26tBidnlMPzv72YhhxkFHJbjg0ccQhroZ3cCZV+AmLrdsNFLapg5Ru0US1
BCHFAs/qDe3FVbr400gCvQvwuEhArpX98f8JBmYpmfI/XRwuG1Ao2UrewhM43FZMoWe3IRLLAPlA
gh+WfkQ0mrVKetM8r4JSObMl2CdDs0rV4NPn+Bx3RFIKnged97z0JCl9i1IZVKklynE3ItwNOmNi
uJc13mwdSDFy7Y62I+eq36A2SL/R1idWH2VzsQoWNEl8Ij7rRJfdumITjmf6vwhk+0gC9mAzHchg
jj0capZJLSESE2f0UyrWXkvxi146XNEvPSvp/Ro4wxFyL2lQ0ofP2ubChljKO1nLycERUTFearyk
G6BZHcLmliuZFs8jIZsqzICYl6+sP/YFz070b9HYTBHXHf8jfMAe08XCVIt7JpXfb3Q6M5JyqTp2
lJrQ+Wrg/AU8hhrAQl+rUlQcRygK9XCNaRIRTWNtRDfPVlYHfYvNTfA5rn4D3XPsdwUvbEQfwSHA
ApF/DePQVKKGvcmQPwgcwT6L8RUh8mX/tPA/95cMcBNh/MBk8x+RXy3WxCZlsBY+TKA3EXQj2SaQ
zgyUPNDgEjkT8MGsuYN2BptzYr8O+PirD0Ovbhggz7oMoCn3MkHgbMFS6VQA7jtJEj/B4o3B/vm7
Jgb5s0BhHIB50682HCYZ530OohZVNNafbY5riBiTemYRKqP9QogE/bQ+D4eWl87SJG1n/OiHXLJ7
ZMf6w9eVc9Cs8KoHvkPVmtcFRVKQ0TVW7/lZpB/XcdJs9/b3oe6b8xPLaPAKQFjoJuCs3CS+//mi
x8yv4432wP9LpyGbGC/07SQIZ5WK6v+BUfj04Lu9uGGX+ii+E3MvgSsMUmkE0mKszn/b63H8cZfG
YbLjUr7Mb/NoCDyIme7BeiR+AvLK+TZjzkBjEhiJ4t65A50HI49m3Vqg1DEMut4Cq2pGUqkULRA/
VXAqLJIVuYedBkEFKoGDE4lyBzwie6bmC3u1nawXAAShPfmETlgDCnUCRKquN9n+crhgwNZi11vl
o0GqWemUFz/48m0ZXip80QuE8vtAf41AwDZeUZnWKg6DX4dtKFX595K0tXCF1Ytby96MDjti7giI
SYrNbhi1jizLppoT3CXxOWH1hxnqAC2Wy+n1UW1lLevI3nGbBxF1Dy3I2q36eQ8OHb2Ayunc7PzV
Vg+e6iYzzNmvRhzBbnyWLDl6ufdhnfqYMy+WaDTDy4BZB0r74WyzpZ3XCWZMbWKzvOvHzSECpklK
bFzR24ztS/XWx5ThYcFRNjq6hCWCm7fPAbw1eAk4wfUaQTJO/0Ib7dFEgYBhy8zsK0434oyKhTny
5CGIaNw3tZXmtvBfxOkwpedlLJrcSknNE9sTU1Tr+5KM2TXmslXkzBeSoKXtLOCYJQsKKKMoNPAV
giMZAeaLBVbrM033hz2xt+otc8ujrNysta4jOy3VuNSRh4fEdSffuXjkD05SShaep/arASarCIsF
YoHVHaK+N+RDu4Irghhs5cCQGcJAf+eF+TOZ5hsYRMrJcHq7y9JnknnVHr6U0N+gIzRnTiII9S2V
wWP4JtlnqUz5ikapszL5AHQnH+tPQr7/sC8TedAZ7r3QY93MkTI09A2mthQLey0KxseM6Chn5UPC
Cud0HGtml7HLc7ve7NETEmmDpBYlHT55gQwGfeQUoXh8Kt0bBaZ+eOaDIYhuvVkIDW8bVmlOFQk2
RsT6idK/sMfqEl+BIGzeYQzIQRoY4BmnUtw6YdoIo519DqvpPDL8MjhaKAaHGKbSkTBhHjzjx0aB
9q34OhfUSsjIyqKu+IiN5/U1qCOvBDep33RDURclKSw6bIuy+Teb44x5UjIaqH4uZFEK1Hc4w2H7
8O2r0vWVwS6zp9AzotUdzJIU030+F9fx+CLM/EuJDzdPXi8y9Nz6IvlZ8GVQuzpOaoVCU5l20PHN
kfrqR60eRn2CLXasJeXCr1zIwq+olcPGJr3MGyU8wFbmID81H2axIQOsz71s1uelju5oG4f3gtJU
gxPESrAkJD192QKYXNCJiZkzvuCZ/2kuE5h0k+DnYqQNIA2aJ1pz3P5Sa0OYwjsBKaf1o5SEfM01
9D1Yu+lHgz6E3aY/zwKDQwx9koEjEJKRKWzrUMWpeRJj5e7JusNzGxxrkI+oTr/p+J6OdOWCA6NX
7CyvieftMyLmAbiaz8+sVLKIEf32JWSUQRV23wxJmfQpR6ajWrpLQV9RUJrE6H/ae1xKcgtCp6l9
OOStMPkyJGVppJzjIwN0J6mv3iVa4eqez6FgdjwD47v5muYRBQ8DqDxqK+fwpLtBMhx3b+MPcgv6
/in77lkbiX7K+fGuaTOyun2xxVRR0mDYpE4oxcILUc0XZF6HjvCGR9nOTfsw7IV10hyMWpEKQFxW
6BRY9u+XZELZuza5K7Ncpm3y7lY/lsIldqpXVEVTJRcjIfhGE06JlguIK425gWdesADvTWOmZbWw
JpAImy94vKDCpLlalHNs5HyfTzMis9MQV3rPhQ/1UiQ9oAMPNoDCO7hZQLmqdwX2RVP17kWNIMo3
FBJrr1uKyEg5zb0k3AUrt5Xq21a6C12ZwZ0xvU+KX15tlQMnnouVMJxY3sZnywabK50UqZWTmXbt
y4hoCFpsODOWSLfrhiYNRSZTe9yehDGZ8Yu4g4IsEGBNEgm1BAxqDyzNv7LmLMZr7+/j/mo/usDP
i/Du6q3ibfF/8dJwFwqccZN1M+DMvkKOeNW61g8e3N1avFify2wi7V9z0qp7oSP60hLXt3ZDIObV
ab1yZlvq7cBOEqxGY2rvk0XzKFviw+DPgC/aODp1JltAWx0Yfg1N2j0askFSzNO6HvLSMEyA31TX
a53CADv8FTE4OpnTZKZTcT5jcuk4UBwUIzqVfMNVli59GIXESUjvkWRf4HxBm+/uYgsdsFtVQp1U
tbG6D9MT6svRKAEEWSyi8SJLcAEHBzHTSXccQmsuCRVjXhJKyqVKpVbNNAhaswp66VMENURsk+6Z
O6PPqDbrwSBtZN11vBFu2gOMfhxvDe+VNJB8b9NhqB6Yk8PFgEbCCPa3DdLCQVxkFAzZFosbeDdi
P/TLxF+PMdmhChPlyy3rvf2+h0xZRDVvTvNH9EhoqYKlieES5fIXPi0iTLpaRjwLwvZo5H+DJDtW
Wbbj7wroxwLlvTo1safBc04/SfNbh2yDjpV7eJFJOOint0ntV7+thUtV6U3ir8meAnd4dV3GN7EY
CA13sn7RnDO57m6LbDhlo0xTevm14yh6PiiNxjclKpK+91U5gfULie5Dg1HKtAmIT4BQUW48lF2B
3TA0u+tvqBRyvo7nA7frkL7Wy8eVDFWXktWSS28gK3jzVJAmfb2HoLM4EoLZ/Sxq5ewUHGla7+oo
PUPHLSbECGupZ/jAKRFz5uC6YJGroUtG9jxHdaRiJXaQWS7gAQ5PVGn3Mle4AdYYWr7QMs0YEOiH
1XHqm4IiUf0F/vRuuWZw6fk/q2L/DKmVBAzmMWC/hdAueRUNWqe8CFBq5WGFQZC/pJ2X/m8WhvcN
2QK0P0qDN7CMjYL/HWuW3qqzVseY6gr2vVroFrsdWNhUmU5FfYp0HlUsbjwz8D9WlvPlQfdzXXMA
YBeo4xrD+mWy9zqvG2q1cZx1T5rZjZL+vXP9iIJq/P2bz4C6cnHzG4r9+jsaSpgTzBc9YHwG7OBb
vPQuBiuf30e8Mkp/OX3DL06/vGFz9MQiyGMc6Le0Y6v4OTZA1YzvcGN/WH5x+ahv6Kfn/mmcJoUq
CmX1a9AXSaMdjt9WFi5seFXijcfGEKxpZyuhNxvNoxgIUCLNL3fsyUUf0au9XXi+eKlwcISe/JK0
Sd+x2bMSSaHp8lBnjQQyGeifpV/M7lvAoywNg8lImlgijNSJVgfQXv462MHcoLsy00r0oKDpXpkX
nbqGzXbU/xxv4Y5U6Wi4hgc173HjLeNuWv+X+VK5Wp6a8s9Zim10D1k30vybs+S+LmAS/Yw5UEOb
7Pn6JRPpkly7XJr4Mw41kfpApPI0NpktIGBKuEC+2s167NE/1w1vQ1DoZTsYlxpO6DU6zHn0YIk6
3kAiBg8/7yFa/6FggQzEpOrGES76iYsyvkHfUfl/ldKkfcmZ4+ex9yXuCWE+NK53u7SIpIdAkOJg
jjHRjoO6+jFEg7Af/YguvoC845mMcjCsamwCDVXpAyAL7N24nypqBoXfweOJEOvGvyIgORoHzZHe
lDP4peioZXjtx7vBLf7NYRj9M7XdlkKIlPoKnuwa7VBRmzBLiWXrrz89GxoG3lJNQ45i2JotMTnd
OBiryYBhh4hCXzET+suwre+ZsMTxTMcwFnGiM4Bp4ZBclFPPfVaYxQ0pE2Up3A/m/XSYNFMmcbS+
Mat+AHy4UcME1KaQKir5xgJ3fAKfPojpu3dwuJ3cJnTTAwpY3kbgOsNuA7l9knfJOf2rG2hr8AKA
k5HTFPn6egzKq6kFGrFcMOJcaLXDU2mfFzfvp7i/KfPF2fApi4ayKe4QbNKVNR2xQOH6B6tm0V1U
S9vBpBRPz6ly0hCmOD5DJ/Z3R9SQu/tnghdEsCt2y4nluV2yGBHb553/djMP2HMv491DHr2mSBpV
4AvY6oSO6fL5K2pItr9KrbdybsaCiyTn+aCgWqbz/CeVaX9EE8OLrJ1EYFm11qDVSP75x9Fiwk4o
DvDhzXd+BGSPdD2253IFWmbXsthtLQLB7LoSlgLZfStDRPLjtYYXF6Eh8NzriZpsZX++BHUsDLGd
mMk+PfmbiQqblfqRvEdaQhHJGZvgjrL55Kqvkt72pi2Y1aH//uG0gm6c/X9pzb2ddEc2RCRvHwkz
wqrO5nKU869Z6sDNSbwld5dstodeLcR/pQ8RsQQarO1ApGMcVEmq7ul5k5/GNrsdHWAvztZ16jMZ
5TCdNLKO5KlLCjupsXAVDXH9/K/f+E0w7toRvHlphrZduo3i8PEWXN7PTASXPOgoiQKw5EuPpfd4
Vsd6vpsnXfAXlsx+irr7r53fYsRdBeZdJsTrYFTSK4DIWf2xX8FZTFp2hbmtBUmGvrIbymYhHeEN
T85wCuSJVYBHiD+Oag4viEcL0aaqTE8OQFXh1el4sO6HpiN/qxy7+FIIss0PdVmDkQz0FH2MbVVI
kJ16h0V9y+uUiispHGnFKGgk/4OfusfCjNeNUitajifzfKvq6FQbYBQndbu/n3/6IR5TmBhBNarD
eu7RO5g5fXTrLG/nj0+5Ohed/s9DqIOLIDopB9omoJl9DrGNlRVf63y+gwTW5pd/SYeLM/r58dgV
tu+XoaCBXp6YtaVuPqLs4pdo8X89fkJK7vbt+hp+CX1vdQVwt/m0bL8++9JYhZkdKU6TlKg1dxCv
VZfXSrYP3/QVkgQD07pU2gaAKapBFR0QjLEZmi0jWXRS4ns5ofKL3yH4j34PNS5wV9V0mc3rBFuz
PA04TljqgSPsat3FTARJ2SWZeyxXzt8J2FsjET1rDoNnwv2YCyWAsBBa+lSmPez1ZPurG3oeyibV
HW7cGkdydtTnnw2UAiwA+5lizJZ2hQn+g8kylds7aQvzj1m3X1Tggb7MgXQoT4O79703VGbg+zL3
aaxa1vS5tytCf33G0Z+lobKdiz72/sbRhcbKukOuc1iLiVOcQpHYUk8EPOWScIyts7pSX3+1RngA
18OtG7V0/Xe8Zht1bGTR4W9Y6uL4fj7ZM+LOUD7S4GOaaVKKke0RMKqw80bIOKAxn7vc13jlqnQz
Cz4UJCnHJkEJWNla8y1SvvO1xJoZ+0p8D2ljY2gRAWPP4w+A4IWIsufziPmlNRTjKR410xCcR4ws
QcilMN1Csv6TuslR/vZBpgUxq5P39x9rO5tuxZeL0b1m6ik2DiEWjOu7qc5C7hJix6SfbchA/rGi
KMU/YBbNK8lFWMYkMR3xO2vTphUdhvzd1MelSnB784fKptm2P9jzI1ggK7IYB9H1PtBBlstKpX7w
nOmOkJMjjEbLzpk2oSVpyGPRckobBA0Yy/C3D5q8C/OE2caBByElgI8lAqPaHu2kfkz4weHVqPpM
Pl1OJ0qKyfWo/DWo4x3hTrammBL3uRqGC0w0f571EuYfi4avQdtDAf0yfmuPqlwvPKGMn9R6hEzj
6F5FgNLtUpnh2I+XJUjr4Gf+46zMJUl/nEoItEsxQrXr68WBUGao5qh6GDGUR5+7z0kob8Y2hsU3
/avkFSbCfiymv8ZmaY/0DQh649WTjNFnUWck9p81JXC1aqIuBgK7HnVFb3vmc8K+qO72tXYMxEHb
djPCZ0/1wwJruVwmMYQ/WQYEz2sS9OEpxq4r8ihNs2ROhbwVPoeuUqH51jeYK95zMP87n6XaQR9P
TpbNxscsUK25dHJFDOS78VwiMFmlivThVMpmNtNoegaYpgsRNlYn7+p8pJpkmCO0bB6IQIwpLztz
aodJQKt/ZIBw0Bz/sBShLoMOoELPYuEyXM3/cqHBvobQ+a3PisD3VvAocC6ZXdQycGdjkK8V9y0w
aDn+HHHVknB7ywjo4SSokfl/GV7qUrQOb81mmKmrkM9SyJn8dqDL52Hu3jQJMuKLQvwRW+OBpMff
nke1okqBnc03eAslb/pXdtcE8YldPkCyi9CTHhYWIDtfzx2m0nzeSFgz46/v01DRMnAl6WWk57Wh
YVcecyqQuavb2mlryyU/g+JaCofBqnMrFBLyfQ/DvPMXjmxARm9RGfuCAt36Xjfuj6mnZ6vsvhy2
LFP99v3pqPUpA4hMBYAnzdWLNS3/9TMYN964xJNCu+q6nmmZvy9wuATAUG0Xo44peZzIuKYDHORc
DmIM/TCqQSSReGP+D8wzGfJF8TbFfRtTmpFaTJxofkEoDgDmf62jrFUfvjbHpKLsHxdPxO87ndlK
VJn7L9HTi5yzpGTKbGl6qOMwUaH/iaFYOc/bO5WyAO+BYSBSE+Le0FIRSjCC2fFjUQYEZ56fWE6t
eHy80HjGHx+O+yRhEEgGQjTePCBLHjE+H5yquTCwCccSCZaCosAhoMsOsk8aLutZeeDlAYMQqkWs
XMoVtShxjg3V5YToSvjl+2XIQ6Rb2JtoW2YtA4km8JVZgXywQwBhr3cmoWU62D1hxi42ud2JW7b2
sAcY/hoHg/DIA7OJ/HYx0WHBy9NThIrf+rDjhH5jXBP37M/HbZjTAtCKUoCiuAj/V+leQxbhBWyq
Uv5wqgceW/h7+5SdbjmMuHJMv74tULMbUL0EQ/t5uDjqxSfe5ceS0FPlXcz9JdWm5nKE+uEn2Sm2
RqgUpfWBrEkjexlSbqZfD7Z+mSwNBPVa+ggAJcDSyFyo/uwunUe0BpI4fRAtwvjFllfqL2qardy5
jqY+M716kYgSBF52E3SlqVyQbXhFt2eazPU/r/IPQeXyqe1rgayIVXbilw/CClAJX8j+tKExhqK0
+kkOTRrtl7P3vmahcyyXd81qK5RyrvPYrXb3oEtZ67TrlAbRKTplMi2Sc71q8wXLrHynj2z3ph/s
/goXqTGhz/FQXwUBOEtHo66E19dDldY+a4bmkTu+27iJg/ZyY8S6N+20+xofc0pZV2Pt7RYsVrqv
UWSZ886ZFhnv14euYkmVGhQRFQ2t/Cd6/MdCslABp8GcidZJX7cyEVHcU4avxsBdYOyHYPWhz3TL
ZkJB8n6AYvckTajEaLgRioTqcy+4Bg8QMmjeshlJORyLbofeblBViHyvJaEwf15n+okM2AndOcVK
8yPFTBdI5aKH7Do+FULmf8i2FNBNk8Dn/8dd1FSnEGI8k2iUhgxe8ArpPh73l1jD2Vo0GftU6+ow
6V79MKdGGdk85scwEdoEPFLU47yZ9KvAswTwac5f4GJvGfL/JosbrBYydZawuiBS6dnWOpEyw7zf
xDxfG5eRp7rrd2cwhyECRUqZNSrZtc0HqmV8GrMCz2lxX4JM6noUcQ5sIbei3ppTB6dUVj50d18B
x45DOn/xNzMDh+VutaH8EhOzYlJrbhzmCjoj4BOCUKFUiQSWRyQnLEvKMG5KHJCNz9m6wtTHIjEZ
zA3rpvram+30MVjiqS/Z13xufU9KnGlXeZsequXgQRMEqcmshvpHFrZnxi+kvQt7x5kyQgmtyfgT
kXPzL/cAGC9Q//p79aHW5xKDUYJxi+FocUQvn1C9hnyarhF6iXfojCZDrcaFSO+E3V0KyYfsUaPB
z1QMbub6ndHKCvlQO6400zsrhNOW7aOk5yiJO1wsPKDfOipjCaY6p2SIoCHChuA2UCHsCM84PcQQ
xb+2sAGL6buR66WpbGUbLKo47xc1uqPXqKSrRXl5E0RIWR2idM8vAOESUwqdcQKoYqhpUwB8lIlK
sRs7M9W62xHhmoUSJ6RtwIxKo8DCb6o7dhHwxvALdaK6eyRLhMcBrXAf2Xzbzhc2k58NDRMesbFr
VNUjumdQV8B2GojFC9octwOILS5Yz5u2/5uPhmvv5sMkXHtTTQCnA2QAVp9kPPQFVSnAZKELAeFM
D3hBcfNNfcZD2/v/VDqQD5n6g1v8L1uqW1aXTx3CkhATsyzt3IaRbdFo6xOh82aE7L8pVbVSJDvF
FidWMinI04OqWYNZd3DpNOoIuiXR1MlGf7XAeE0IBKzqxhpiUU3jBZ7Qa4X8jjFjdgJzrOus7YFS
+ltsVr6MELbxpfqOitl4oMF/MRlXWUr3oyTKAX0KHWXhrr9cYtYAPjbInfQW1vZi3Le48SO/GLcZ
BRKg9nDg3ydqQjgDI7xOZ/S3jnm3oJFvZbRhF0AIqT85v3lOr+dsVaz3aatLTGAWXZMkmwoPjhne
Xq1PvDeMraNMQgirCqICJYRicMcMn4Lj3gj2EtAbGGq8wJhLdJDybobvImWUB7u27Mzqu6zX9nVH
UT5N/DXJYSzOqHIEsiSLM9XTt5O36gzg1S7fx1I++ZQ7thPd4l5C3tyOZwMmaeaN1A22ifrXn6hI
kOXAOHZz2tnGzlGbdWDDvw+sVhCSh3waBeyXNqfWGbgxWTqK7K9TZEy1pKGOE1qcAs5kjop/ztt7
n/9uwSQUu/W90U1u3NGvw1CqEPd2GtHbO5FUnZtdjAx+SJpDexqe/8qcLxKsyvE5IZHjTCFC5Ps0
KPrTZ/T1w/mzPCxmNywvHuV3WqFjrsn/yNGh0P+fX6+dCVP4whR70uGKdF73/grBFMgEJUeB2Zlj
nDdG3mPeWUNlNCeq6eJXtal6rj0OsKv17WAEc3Q5lqnMy6k10fpXkXiX3vWjZtOdOd/tBlGPZiv4
PIQ8dlBXl8xO22uMEP7DdraKYRdZif5U5+EbGjR0Tw4vmfVP8ADU/cK23OO076JMJ+SVGbDP2Mf8
pNkIawDfOzY2dl6ndX1VxdL9jCIyFCGMqc5xMLdNZ2Egpd0OD/ZJENXtQrXQBgjtlr5beiwIHBIh
vahcjKz2dIH8iyWPwiJmiQJS4vygbl5/2x0X1xdnmcVQJcGt4zdrR1PPyauFwfCpOqkB+79AfGNh
9YrYnvDTnbenF7+8Efb6aaSC5qsLcB2He53Uryom0SO3QK06CjFJNfh3aWadFtkde2sjVUAFKW1e
I9CmDKRd8Mh/Qsk/gP500cmo/knkey98/g4naHvlfjYwrUVOLVVYnWwjU6cYmFkvkvONiotKHljz
h++VIqplU85/+lgq/Im26ovtlg+x4K3A0TsJgLqJoDwpCEQGrRmriTScq3hMbbRiumlBJAU1Jhi5
d9I47eezkpPFYUjuE3bZj656spvs2/QCyrx2uRNLvvH5LZcybBuNyVci9X/CWG5/y+7yCe8NYkzs
/PgBpcAB+TyFqR9R6AF3WsKGgrKtA/8h0EBIox9HMx1OlRw7LU3UfllFnBrLGK5D51WLPMatuFMh
9oOqcUgWCQeuQPbanooa6o/jZYOvN9Ml5OwLSwtDtJ9Foq7hob/lxDtzsM5UZpkb+2tlpcSc8M4Z
nOYlD4bOLMaWHEEQWtM+otGFOrFWOwHYaP+ieWIk7QExhT8L+T6uj6OeOLKf4YB97zUUhTi8B5Hy
+ibQlZAStlP1tXcVVD2f9T6eqkSR43jKvdLh/GvGvHAIjAuSxnLENefQ6knbb5UMRJbOLd3BEEYV
Oqn21lI+fffqlHbnbOt9SGmUIq+rCXq0oQTLmH7lWwXdXoRsnOte54zBpua4ZSwR76BSqqZXSriu
8RvvBGlRO4SQ+CMidkU1rnIjzlhLsZFSKFd+CN/xpalYcTuHQev4Ub5VNHRUalHVeoFCut1i8Tke
+vCkFofrEMzN6zFzqUGQTL9Kz0JuTidZ93sIhDO05XRd4xGic19uGUY0cVx004MA9HY+PcNm8hSq
6z+WPdxNE1M5/VzbXB7lzGb7la1/vQnOMkCifWvzzYNyfBX1PpuRM2hF3HCj8wj16yLSHgMT5dNH
EDDuid+QeqsYcrh+0vg2vvXyZY2AHoaoLzWQJfDMyH1H+IjXDc5v/A+XnIVkKcV2Fv0yX+VKx0NQ
xJ/ZHNQMtFw5NF1ZXBiZ2UGCMMbuPo+VMv1DceO6sgN5bQ1N4FE6/i+F1cHkZ475r9KR6/jgSdMf
70tl4eDDdXr+j1+OCiDHsHzoZzelfBwCyDmM30hzX+73NBj2LCUBPJNXSHhzeqC5/UUSQwYFo32x
RLHGo6xjaXGi4+yEhEGV0sFDnR4dSq4VnD1bRufZl/6O84ZQ/SN1xBPb/zVmS5kxSiMbWbmp9oyB
4N4sUX6Ri+RNy1nWr9u4k6bCPV0sFcC/LYRbcc2OogUszGd/oTS09jj1PjZHZQ23YsmorjUukjuX
KgCzoYVlTQDQTY6Hwjq3miBznGomJtgJoXvJU+hFVZYXG1XbJSq13vjvbe1sEuVpeYGFh6QeukfI
MbgAL2MxgSRgNZ8IZRD+OU6Fg48bwjXWH/IwDlFQMSnhPjvTSzx6najra+TuQiun8N+Dh5kP96Xx
m5YxVjeoR1xOniA0zxk1ZL8m6s4I7S8bCqmAAIU/JBy7JP5IJIEatdunL82JAMcgfKGDsglcp2Gt
EGFxgWJj8oowstlyeR7BmhJTzTnrV4BqCtHER2tFx7Q/h73RCO5lBjhHPLV3ggoTweYjjR7AdaZw
8J7MZ6C+ijNTbzcG0cTBjRIU+RsiwqDWsxL2MMq/Dt8jz0kOk8VsXwUGbgiK34nTp8ieSs+edR5E
lzGq8NQugxw2g2BglR5mWlEYRaRD1ZK0DHg2PPo1C4EmqMCAKL19XMwNH3RgKrBEtOlbTVrnyz+O
oNgq6bjY9/fL5gXLZlx6YFlW2Nt1HEoaawcBBkzq/4imefoNAPoFW7ZWTEshKU+f5Lt+YfKO/uB6
sCvqEGtCxr1NlR/P5tYPlrIpVhx0T++WKcSYkOf1Bk28g4sYwAlDDu/+jTOT9LXwiDxAIx4+nAhb
IlD2XncRVDoqFaLEzHFBtwi6GkFTJGnBZBFN9AzB+q0arl94a8/P1rflhUrow2DNJbjaVaX4/26O
J3Byur6h9A1IH1rmQ1z5BzSdB/8s9sWeAgJO/dW/IWs8g8SA/rB3BJFjH2k2gzsTTu7/lJd4sp6I
b7xcwWVHQTyjxxYdl3yx3qOHOm2OVdGSBn1VfzI6Xt4m0nW3yEWmrWGXLLe+gv50JVL2vjM+Fe5x
JVx+2w5TXvKPiPpltUvuawhglN9RwGuM0XuNYypF8wXJd1dyDIwslyZcjgk239ShvI84C3GwYuA9
Y/QhKVJFVgYZKlTQHkRCDDZh3BxAbyRH5R98fLrpIh5tLMR08nwvgUHHkEYGHUq7Cd6CRnZ8Lwte
EYdhxO+ULRRqfJCkIJ9z6QvWStdnKUr61IJubx4BwAQWq8WgAmzHMTZ5HS6DdryB1h6PK4+IZ/Sz
Pto1AoG4F2kkudmYtkQlkcGx/6Hfhe1CgKi+XbC/L8xJJm2tg64r7l4EPSJyGu7IafUDxnv5AhLF
fEUP4B/hnLWa3UhHkIPi6WXm3s+ek8sKsV+h/3P95nBRbK6DwL56UhjOc9o+6I4HY0lp6oDlm0Zo
u2Y9TAD0a9nTbMXd0+ORSuplJu4Ntc+6HWIFE13SQeE876h0xX0aDFMXA85GT4TINuSANFAEyStr
LBouJcfdMt7gERSskntUEvK7uXDjeg6rM6WXA7dy6q9GrH01ynWQ4CiqikIQgH+D6u42XZwMUywk
tia0gX+HUS0S/gXROoPE8ulNGTbfDu1rGHDaX1jHzglhVfhqvP5NPVnd5M4pF6K51R6nCwpinCtv
Bozy2sWkdOaXV5uxUrJeCEpYasYTO6roI1GkImbEW4oGpUc7qlpMz5t5Z2mGGypEQlRVC3yVhz2r
OigtGeb4Zlk8zagDm+rWPk4QOHGRryf1Yt1WAXtG183Hrosr+oUjimc+CA9yXPr9urukf6PGI61b
2O4dbg6s5ptgBByMGbrroLh8tWkssMUUVuF8WAlTtlgRLCPfH9comLM66pkWbKoO6z+rXKF581K3
A2QLW1YT5NMeQN74GZbnxR3sOI0qZisHVqy8lQtRMenTLqynoWO2m6wWdj2t8Wy0jJbnpm1BDfq9
f6TFVTPpfCrvtujav2HKaglaIbyRPWbKBKrDEdnJUqifkaUj5i/fWzmKs/H8gAXfey+4/eXLCDyJ
pgBqdGBi9Cyqb9LJ8IqzpnKJwprzN735O7o+wiDjIr/UMoxZl1OGQoqhdz0AX0EnYOnR23wiqj4Y
kVFxfP/Ny8uDVWWOldw5dW3azQKMmWklEqUQbH2VbfZJCehkpUF5T56F+mXjyzHA0PAVMv1UB6NX
dLt1HHbUV+6y4TqYTqBMSgwtkbIpJ0qeYrA54Ss64r29GBXlqX8wBDSyM7na9FeaIutMwGdA+vVZ
N6nCnCroQa01H3Qkb4x8/Vx1PZ49J+nJiNqroaeNwHY8+rDAlH9pqUaLuFlqOvm7GnpfxwhJjR7E
rgCjNGsF2Qa8hnxms0XqYzB9o02aOnTN5gvEdRZELmc6VkFhOydzD3ArKlhbmPncQ48daPTjCnDp
bjIiRLuo2a1viK502WKR3OEZvolFc0WysfvEG1kZhxfZ1UmG2E3xZB0nKl1oXd2EDQ4Q6GZdwfae
/1NbrCGGkuTWkgs0wUg86aS4cxbU9vEJFIrymfcOuSEM7gKX+DizLc6cPbEwmFVvl3eo00IwzktF
h2qEIE0/sXxuMdBBkCsT+RYyL0QuyP8nB3pWVqW86nTGHMM0lBqubs3YMDo8tgC5tF9BU+otFynu
z0CNPaU/c5m58zwo+ZZbyTsnGIQu3RFYYfR8WlRb5ZAOtTgSSVRUF5v/noaqLPOi3K9I4j7zNmtl
yEAXPoGSaajvyatXPSeX7fZ6PhRGsXjkI2hTNxFsGMkbQLKQ+bNo0H8f8FlQ/CZG0LF5t0vqV7lc
I8qKF7NfI4FCE2M+likimu/WW6UURT50gnkbt5my25rtnmGOUHiDUul1IdOBDECm+MlcEpJJnI4N
dk6a+rJcJ9tj1xpYqGDgxq6DT/Yr/xbkmXOqp+K99wMkKvk8zb4qJxHNIFA1sjp7JBUmhS5McGCp
9/O9Pazvy/vCcBUxBP4LxPf7aL19fOTm392rRRmx2cSUezcXBiqD4w6/RAgYtRm5A9OV1iLkeo9h
TJOPiDKKT29g56+eyXzyDIlXy1rU2t8IgonZZl5JFIgkckcKne/4LGfTMQXdxdP4HtAOuzJ/u7US
NS/NeI0iOundqnv58Y2p0IhwHDMxOHrme+mJU9wqBXosZGtDapTyIZ6QjqNaYnada1hx0efFbWAe
NDHwcmkXHtA8Ioyrsf9JwqHlgc8CO1L10Gzb9efBOl1fSQvDpWiwvZn/oHIzdolGMmDzYY1APsej
QzhLJYKKTmeML+tpkQysSUGQRPjG8Vn8N0Y2nHHuFy9TEoqbPyc6mGvaGHnjQSorPuZrCQtKdyHz
D/d9grm8XxoDNyfyHM7crXL2Lly//zB86ZqIsQHdl9oA+wgMhqlmvK3vFJxYGNOgZTRffd49nvq2
lq0uSc+oMNg1gKvOIa5ApTt5wAt5bsm7jyYqVGmBavr7NDI09OnWosCp31E5bY7cFAYv7CToKKJL
LkEJWr7FXsZk7Wwc2mZzakQX0aE1MHbX+XI/d9mr7ay2D8Jg3c2uHIJn+FIjT86/yrtNYJTOC029
xlYjbBTUG+KlgBzd1NkntW96dm3W+SbNGWb+GVaNpspV9Ck4AtYD4xAdboMJtLepQcUcdh/OQL02
icxarAN5MxHIuw4UyiWOdBQB4jeZMHmRN0c6wZ2LRmYPKWI3jJFyCdeYy+16dcO2uMSVaDllLN5w
BhQWA/BKtoWS/wCCoxfZHNIpd1gFln1luLIdyQYUfxqvLubEoxYspOeZWh5Yp+9vJ3MGN/DjJkqc
vG+fdKisL74O3er/i2StB58aBcE1RlxYG6iHWHXCe5ONxrxKSgKYqO+jgqk2hwCCLJpXfSyVUMwH
+k6070rmInmK3CVD4WAKdpGKmrt8hLXvuRZWZumnyv9oM4I1ynEVoOE/0R2R6GkuSNvNq5gnmpeL
uX4aq6Vmyd235reubxwHPVXyfi6f+lMoPeALBnVjOQHy3ufTAJpMgucszTdJkdnBn6k7gZZwDW5K
RYlsyIST0XH23wAw5TAOmEiKeLVUZjtXf3355f8EB4PH4mv8DljTVvWHKWBiRxbj/KHxA4UK+0aL
wWOpXKbQBhonoUiByRfWu5xWcfB9pDZ5jmMU8Of7VMEgxXq/aa5TR8G69uX9RM1WaatWwFEhx0KT
8pzdGPuMWWv3G9fYBGJv8OBRAhNRlvAhUKZPDJ8NeMPZmqlrp3+knHfvs2HwnrHbJjAsr98KxhIf
BKDCoXGPTwWipcM17yRXkSuVPAy8N8NoCFIqm0qrHRAwlfYoShhf85zQ5ip3CevabvdbdFADZUNm
KcFTer12kh4WxaW4t265IgdZzOtpMiA95LAak2Y2RMoTOJC4qNrr01dLOEYXI8Hee2YiwmxH/tsY
ywTunfinj4OnUeBT48gfusuqcKxEvEoa8ltPyoMEKgKRNEa5lNwYFXthA/QeZYMKKFEtUMKaPFMP
6w/khUR+Smrm0RSMwP+Ytks04519N78VllQbupa8xHx9lm2GRfqM9wYtUEZwyk2Sp5reQjvtSv+p
crpolt5/ydJcEP60TGmjptuNZpglxlGNrkNjJW1n7uj3L2lhfrClHPh5O06ArK1q6Z6wkfeLl1VP
u8ugn2iLKGX56msx6QzqhtcJnXZXMP3naSwagfNM3d4XHGlyIjFzdRhukQRM9eCsd2/4eDZEknI5
s9qQyDw03lNXhupcULHbdHLtZz4BVIctJR9cZ+p6MNsMIAqPz9Q/lly5sfJALfn6cADm41mQDYtl
/nN3Kdp84v9WCcL00agnFmbh3pBgmMwHfFMhgZD07w84d277mW1VyBEVEjqfLWIANUjKXr3B15YR
RQ5bnLR/xjTP7kpy7agWCDctrE5NrHhIUPA9MMqRc1daXGfpbjwBigyVBlng5Hr/PABu/dm9nP+e
NdQzFTm2tM3ttVQ95Cn7QleHBGZ0qlNibpyQ/tPTuCcCm6dnnbeR4NNh3ytASL7YT2Z19D77MOLi
UuLS2czM3G+4kta0dbqHJmG4T2xoBhx9dghSnEY2Hge/+CBpTdyS6VYpKhaM9ZAOt6p1rb9XV+1T
afITT+S0yDV5ofyIuzpMTYRRSHQQh1FMkTAXphDqH+hxBcOdUFSf13d3pcgJ1SDQ0++fHq19gynW
7PX28giBzWsh2yGlHM3O3DvR2v8VEJPfY9XGmEx3p2xboMLCs+mgEo618ozhZ9Dc6tgb9qQqK/on
02H7pFCcAef1B0eCLaH0hs0TkbrVW/oTYZyrdt95/5YjdoFja1ze3HUH9EJWQ0rCO+Pfq9FRu3jB
M/PAJF+NRlBfm3ALldDT++Avw7q3ICa2dL0hBSqOkCVEfNHhRzIytDJ9p99M5p+UxjM27A6N455a
9yWAp41XdFPIheRA4qfrmrZt1BXbwlhHMvuvMTzeF0SC0L2YdwtkVSJkokZhhQwfc8Dj/B0jDGeJ
/Af6ecRoDjUSctWwJW4SuaTeUwuF/P2gy9g4O5Q7fQ8ibf9peYQ0SUzLZIO2GobMLW1UkJzO+72k
Q2CeZ2BzRN1R86LE8RifF23LVY16BrETDiCQH4gHNZ6UDToS0Cj1sb9QIhP+zR5LFcwRVRzdvky7
dK5n31iiJ+Ciy34kpyvb+QQtfTTAMVxN0lAtnDPqrjbStcHifRcRY/yyJ3VcTvtHl2BQayLrwqQZ
GLYURELLZVIoyLxLUfVgju5SMMIjj/TVX7EGwv6t85tz05hOF0uNcbUMjerTWWbpVNYg6QUX7uHG
8lv829ZTzFs9HED6AGVYnV2oh9VuSR2qHH8O+Vd+kx65FhsLEJsceMSzVw1JAKK3Cn5aRwoJlqKD
0kKb/K8CdbXBZp0By9/3gMN3DeisEuDQ8cT7CP6PYsCSRg7YcHxWf/SIn2v4hHfwdGFyBpmkg6uS
3jglc7zaeaSZw2Og4RSr7yU6ptZ8Q5aGmsQt4poX+IaQDO8rPdx3XYfz6BnSNo5Tc5Gr1nh8OmaK
syAzExB4gGANmuthb24X9jBI1SBThCB1HcQHfYOfaSY0FK65sFb6FPiJ9Yc/X0TCmnC2wJyYMCgt
p9Dm4Z3SCK6k/HGrCOzNrRRQAr3tpDhDX8EWkr9mO3g0EqKuEHW4V5YPEJxm72N7q3pQ80nbCNek
30qp09AwZs0M7OxuJZPMm+Nn/vYYGvUuNx1xpyHGav+Y5UjpmnOUo6QKkiSdvJKO5ehVLCX/vAw0
MPLuMJTXWe3wmYoS4wUghVGzw+9vbyeZ3MODirB7vXHx6pdbWDlS+u3LLToSMqpNMixTBgRi6tfR
97sg1/zAsWRFZJbYzdi/8Bmn5NbkWkEZUFubiBNN2OspAEZxcAIdiWxncX/p4cv32FjgIg//4cp3
edv87F6QDX5kz2aJl0YFGl7+phOv4/PjBGqfGx4FTyEvROhhsFYFMn633s8dGc8SLyfN//zaQNbu
PVdsMiUsM2D6AJ+JKH5UD2B1b4A40/Rn7fLrqSbzHKRD5P981mMLqn7XGtPPMeDzHOiO7X6n7jsE
4xRWf9l3aVXGQjqYtUtZ0JQpT2qStidHsVCqrhaZ42ocDxQygkKLxP0tBjk25UvGWItR7aKT7LnK
KK4W+cokukmEULFhKJmxrGMgiwqq3KQKMpCS5vxr2sfL8ahr+d0/j4JYHv3FW8zh8+Rg/BYFziAn
e3/pRTf4CT+63rWEblVrG8eN0jwSI6DfUXGTRvqwZU4Hn2X1CWAHn+T2+H84IAcB/s4rpYVBCwn7
NTia8Nr6mwtInej2a+e78PPCzMJ7P6N4YvJeM5n2AG2zPf22KiieSw7E2Ny0hOWgjienFCOt+UC6
9UUywTLbvXqQndrkrWu1+CnmlTPj7v+L/iklV1sJ/YNUPcsJy+8IwEiNTWbRwKa+T4bM7UR8Kfwv
h42sYe2KJS4Wgog710Dbyyb93aI/RlRFCiRtNeW778tgyQ4uirHnnJx32GKJnBE+EocBSQKwQpgS
S5hUrpM6xFT2Wk5ALK/wmjg/Z89rUiREVQ9+VHxhfPKYvRs46NAv5OGVVFhcHZKihTpWiEh6UqW7
kSBFlcD5xFZ6OoLPeqoA2VEz7TfrDluWlEMiz2UZg1xSVkHloP/j5rgU67sFvv6e4dc9bV2axPok
PfxOksDIIf3DD2zc3hvlfQ0uScAepDZSScvIJgoDSFaVlnN+tJhGmkvUfqb+xJqifroIFLsCvGLT
/qQiqy4xHiS/Zc4HNLXo7DI9WyMObW5T7iQH8mSf1xcZQqz6agR03NhAyvQCDea2P/X9smjFE72m
5LkM6vf8w60jRzTBnfzNhrBKbDj4fCgjzHL/rDuQQolKBChJkvwH7eHit4Y2bOcuvCxwFcuywcpj
g7jmQksyYa2mMPZANDaT+9+a3T/sNMv5sM7dDLnQkMbSbOkeLB4jR07pPvPztHRnKaqc0/SCY3TO
0LuAst2H2VnXTDQfILxnWwPahvqMKr0urz2OvX+Trk+YmcUvQ1EBKQKsgIEz5G54vMOo32XK/ACR
9X3At1BF8fZyYqFWn8hk6XF8/oagdIFd/O94GzU3imA9io3W6MVtsCweZ1kH799u9aHmkvqDNfB8
RWa+lGmtXC+riB02+2RVm/lss0n38TeIyu2WL5oBqlIjH6ZJDWrwOWqffDk7sb8C7zPQ6W0mohvd
IMLh+qef2EyCqV41Neh6m5+iFXqK+v3zWoAfGvSTb3SzprhifTVPptDBJmB21Zzkvy7tAHfqKljz
3+MjCfGirXH51L7vhKZYpDgwMqInS0SWTSKWebw+cNRCfSxkbN0q+CVka6BJ04Xp7BJ5cbyjsW02
bBTkT8qGY3alV10zSu8zz5qij6Uw7Lz7eObKU2CmxHWTNPgab0TvOtrfPalAQBSEtjGVMBPHzZiH
D95xoVXNnBuZUsIBEsjPdvyW6btmkLYfd/CgGUI9lk/RbEwHjrBzqDFaPc1juRIJuoOTjqmBfJEU
tIl7zSK6afcLDUt9UGn7LDlieyK5uVAsO+/GiUX/nqdsSj6x4lt3vUbzbt50W4WOBze+GcrbjQGB
EfELSp8JdTmJ2+bMOQae1TWmHKWvf5T17D6cX3EJoDHhDEAgtQqEwjIKQgiSRrTo7YN5MVtIL1b6
PL+4jKI8Yd3fZ6B1whcFf4iIEaQ2bPkDtCL7ggoN4+yuCI9WvGkUkzSf0LlZBky5f5eALpMjhvhM
SrBKe9Wb2wYDCibEAn5YfEFBfSvQMFwBI34ueUJrN3jYsDMfMCsjg+CjWeGGc3vWRtvHs2lGqxng
o8eLtMt3w9/bri2KxToFqNGAhfrToucJzt4Q0/DqJ4tGOWGqsUWC4RAZt2rI0NrebjYuaCNGLDFe
xshUgi2ttnhJ6xILalNKiQUpgDj+icrRdI6ijigAJg3R0ZuTgzWIuGD00ZQw8STfwyS9s8CqAiO6
/envrG8dd0917NeJYs7gtS4Ype3wc8DzWVtby2i9NqKI7F6K0M4k24ICm0+YkJkRWJk9VAcA8oN4
qk3jIlFvz1cF2euJi78JoWl1Q99O92xg9dNzIGKPoyjagy7wJdmauB6Roud1X8iPV/5m24NMI4Sa
3+Ls+IEucX6ZBA9PeayHDp+0bYyc5JkpaZHA0sWRJOTmF2u6O9+cAu7G0MAH5A+z4UZVM8yYm1jx
JhWAiaktrmx7vCss8bOTrzkALCI/0W7lpVW1On2i3ng4TiXAN2HphLTmSrDGCgN5949XOJ+Y1M3u
k6tKK9H+aLzYN4gvFG2eM0QALXUWrmnlrooP7YXQ9PnE9KxoQUzQ4YS78U5lemDMqhRalgGUtxF7
2gga8l0OeUgIYAndAsG6oZQckCl6gyaNrZnQm+cFlJh4YQhynT3wX2lpCfqbePRi86BgG0Y7RksQ
NJJ94Ye2vT9kwSjxG8LRMHm55+4r0hJ6A+hG+uDKIhR3T/eeFOwVP1xTEbmwXguQZFEh0jop9jg8
18xIZxLircJMZk/p5OHT8i6p3zgSEffXb+8+613whC7tEMb4BSIVxFAfYPseEUjv5FYLMvIM/xny
uWC8ayzc9zCJeVdiaZp6t9Z5tvYlrVOsGtpembv6+UYldqCaOuHLBVPOPlVRLMuse2lNPdu06IUA
W+en6Ller6zEURqsvVHfnsxMlfIMknKHoWacjZsGPl7AS0F/PasIu6+ldEa4Uxi852tlZHzenvzk
R9KSWBMZ2w6jHZ10h7McC3u0+DXVhWV4/f/gphpaCzj9HcIWviHJWYH99VxOtV8OPv6R9Pkteq4V
SaUH0mVZZjQUySoitdjO7SD26qVDkFz0eB2hBnbv6zDB1fQU5QhfmN6HAMJA9seXe4EQAbS+GapZ
QLS9sYLu/ywl5zLwTZWa3MWb+iB0FiZvKnzqzxN3URyZh9E/sU3qFrSNabHh3c3uyuUsm2YipF4X
Spzvu/l//YqBlX8DpmEnb0k8++Chf2MCqrG6RZn+5ahRN2HXhLyrOjqb4e73uQwSmtzBP7HqWJrP
vDQOSW5vEZlG3gvgKrSRW+SN1+XRFyYX/+vK302xEaKEUU3t7DDefmxR468A6QpKXwkyPDnMTP1G
6wv2xe017IP+12zdjlNc4TuxoI2PzAWt8OTMfID0O1obEboTE9KfPlz5u7wZM5Un7OzlKII9TIbJ
w8DFLiIrurWNHZtB6+O21IjLA95aMzJ6DAPHwvwzKx2g+iEYgAJW6JoBIm8fopTtI3F39/qrZJf4
MUv75quCHXvZhzOXodddnIAFItRpa51CoKCaC1Gx+QkclBFHRXRux69ABkjovsJRniF4jzjj208e
TD/KGVKqjSCunFwJIFwAkPtGSxaII1rguLXnE9mhThPCQAYe43VKNjx3vNkxQIVyTzOG8t29mouc
J8MlpOlOlnI5TXUuzVzs2dy23JvC9its4doE2xbnaL00813PrcrFtl3IcWzG1mxg2aY9+HRiuSYh
r6vI5Gff4L//CIHswWPi/1eq3Uhxy7psR1uXAGmMKrpcgl2guyYJ5q8kqRgVAHzx6r0cnXdjK4I0
gvLDVo9Lxt6nylF88kYdcn/0E9NAZ2HIT9abT4YYn9R2WEEv0HsdgUEQVMrTUf8DtrHtvA1Im6/y
rfYHSCmRFwni6CUDX+OPAcpFhmwtyDKNA7fFln4LfWXOrWi/GbHTHiyN1GC17hhiLHol13DJGOpp
q0upGtAH22gluotn0SRIKf4GIx3h09fqrsUAY+jKqiUyqsZbk0DH498ju1LDPLAzgPoH3NoTT4eQ
OMvDm/n70754unFWZcYmoP6Rax+KwZfBHBjknwXaxe/L7jJ2B9VZTzZhbPoKHKWSqeiWfhOTQrkc
W8eqgytaX6LFXjzfwH5Bv5fsMjQd/Yg04yJQRK+I7KN+jcLvmQFOhujycSn7hXidybCRaDPQEXsY
oWYzlb+eV5GdE5YfOy8oUOcm0P+jR+m0WfPaQD4vZeQk++/CTrFF37rZ10yN0aHpmJWiZ2bbkYqc
ldmsJ6kSOP0BTg8UHVL82zVC2YczVPduuSkU43Kyoc7y6bQ9FYKTf6KgzRnpO+p9r/Hxtpux8Pau
eNonncmZLqibjB67pPFitg5RdWeb4HmqjpCvDNdo/eGFPlJisIy5H8WYf0pX+ekJIjKuTa2y577y
k3Do9uZe1Hiz8VqOSoOyr5bTOcG+jlkMfD91Uhsi/8MawFgdVNeuSd4Qps9dlrcgZ0gZsp/i0zav
ushYbSdJTz83sUayEHSfdpoQG2mUhpbiq6fiH1WJZpg1PtJoHBRuF6bd1PfIPhWvwq2TrKATh9Ha
syJ8lnIgeIPiGR7dZmjneY19x5LJrY4E7njOh82kG9JbbpC2XBPxbWgke0a1qxF9rEk2WeLLVUCu
iwr8dXT1/gkoCt/IDIB05a0Yg2ADSmGTIheKSEiR1ucu4ShM2BVMms4uzbqauQO/B84YwhmwgfJo
4GM0vjxBBo21DB8wLL8LEChJYBjGCtx5uYS06E/N+WxEHfT0H5BbCVwfKa3zf0nX0aQ/VwgWhWId
wPLbVX7Ts7WnVfbLiwzpeeDaRTmUqH4F2RLU4p29g5iJGrT37gJKoMLfX+B5YiSSwe+hwPcjwPOM
zWXZd55rcExJRcutKjmJqJ617fr+5fHyW/R/HMX0HtZ/zG/f+ZT2RZuwM/YpWp2NfeUip0kqXMMe
eODuTSEV6Fl3knE/NzwjJZRUd0IYhKV+3i04R60pTKYtoxCg4uXFwlMmlX24l9StVCGq9ta+7fC8
fNBZVzSJhtFT/qAuagfUYVx4zzlmxd2DiciwXzbB1ICGC8Q5ujB+ksYn32BnJfiWjTLWFQ3ajj8Y
LvuGNSNYkzU8RUU9hlbTdKFOaTkh4ap9jnQ4yA5NsOkO2iRXmeV/sp+/uD9YaTq1ARCL04iaeCat
or7QxAxkRyTjt3o5ODJIP+/rK0c/mWRbOgCyIAruLFawVozP6o5xRmXQS7bkha7vIJSePcwpxYxr
+gnv0hmUpqx3y3+m58Q5LC9s1MM1H7MOjXm6axL2YJrLmcxHuPwQFCOEQNkrzlzDB6dVdRcNQcOB
C1uO5Gt6OuZkt46eVE4dXZyW+T8cgsKixmrJxf/nPGr7UVADwB7kY/3J+wmKlOdS2NnPzj77gNtu
K3GYBN73tkt84Uo+0IOUVwF81gkXBseX2a4nSY6i0lu64GPTk3tVYpBL9D0mlV1yILzthZLi1GeP
B7TJSIjwOp/6dIlz4jwm5bul1gpO+tqv6eygFHBwNvzbbA5AZWylDOCwaVddgwBDZbghgb5c5Ch5
9s95A7Xo2LDm9H3Q/UZMv42oRH1wKY7HO1Prfg1HyCwpy58VxfIotDVqerk9ku/rGd5ni1N59uyg
N27JUSW70Y3uFLZMl5YNgT1PBjq8xIbjAvN2zzeT883juhHB6gANQqNM8kk8Rwe8yQxkI9B/ygQI
lo6DR6x0RzUD6KO8iX64YMMJZyC79rNc9/5N2LW/Hek/FJTIXdxRadi8uU3E059pJBcXCJXSJq9I
YAdzFHj+DgcVRzJC7Gnsl/FM+9A9loo1BEIwk9BuXps2lIWtvEnrBX7uGslWtNUsa515jDprGF2Q
inNP70Sp7d1ATl7hdtPw1XQfnsJREYeFa/qPgmx2+0LccoKZmt66Cy3jdObKTZeblafCWoQq7Egd
rqhAQvheoc2Jt99NG7UZvsfTFsxIGbh1xwR4eN2hCHF0GG15vQNIWLOnKpfWOGx7wQuJX8r5D2Fa
uJsck4VDrmcodtjSsCYoY1gbadGLF02a3m1aDtHB4pfOJ8kHgwjHoTsY8eOQvI06U2rsX5dYTo5B
M+9vqeQB3LOq1ZFPKukQsli/BFoyVyGjFufYp5BbIlHSeRYAeSB9usc/J6zh5pi/vZsuhFklPrBm
eUkXUtk8ZAOerjPf/Wna+fxSMtxvBebhfD7dkttEsKOeD6rL0IaaoKf4jVS319MSjKoNDBh8Ply9
nHwm17WezCXsEz+p5ECpn6QosxiJPzkLoVyP+uKdJLuKXA8zhHADS6g7MgDIFdQDb3OL8km5Ak6J
vI07ava+HO/eVZHueg8rhIyta1eyoavn4yRzOQ78DZd19DBmQDsjlbMot0SB1ZzrFScmB0CkATgS
QmHf7J9gg+PE9R3+XXoJfk9GKRWeTnPbehupi3IwPxMUJIjhRmgadfj2T9z2s4mj83O0ppLbcO9h
Qmc6OgdBpWdkXciAtOXL7/C61v8rgFhs0SsUuey6yyFw2DVx1JySZtwzHeHFrmBYTS7mLqoOoFet
uk6/LiMGlI4/CdcJK57zUydgvy1Et0q7Hfj3JDkadvQrRlD9CB+gdtXpEDPfzv6H3B1Tum8sz15j
a0HVNydOd9dCFL1EJZ8OQUjLIfCTTAAr/gHe49Yx/t/LvAgH/JZ9LtsEoiamQrV+x2998nz2VDmn
UY8sNyOKWa+FNBgH4KdZHW03nnR5mP3GdJVvAvzkzoB/j9mD2RZHda1XXkMRZ9c6wd8JEcQK4jAn
u7Oj9B13ZwZkyeE6W/0GSzdyrOibr8a7pPHN1aswkQpmxpcFzzskPoimkvwAUg+mVNeVdINTVd7S
h7ofATCX5wlCz73w9CfbgwtOJwpDgLifiQrSpgMl/VuI1Nrj2oYFwH4EzUO8ZdLUgYT0nLlbnYWO
q5+9mobv5XgihD3093i5ZmYPlXtVOqBz1UahiV1HHQuaxDqbs3bBCAuRwdtGm4fOa6bJzKQ+RW7v
tOE3as5q/F+VBgP3WLgpvKjAoBI1ezZHTjMhMcAfYRF2UQgN7JxQm4f6RRQ6BGzrQcCNGGCj+DKp
gBWMiA2FmItCJEwzn94XiygjRuJZQqb6o2s+sNMXQ42R/bDNGwSF1aOymvykZR/o9OmeBf+8xxGg
PxXgRX000HHVDnaShIQu9EaxGHC7veknty7Zr5sqLEz/rhGIxlVTfUjzlUrzbn4A+zwReoAv3mHN
pyt4zOCG3XCE5GeUT4MUVieWIsYecAQ8F0pkChNjUY80BUx5A5KVb/XkpVtIX8ZLW6IniVg7jPyl
4bgReDvnSEjQ36nhaXv08ljvgLYNGZvhzKgQwn1677TslW5U7V91UihVp2iM9A/GX8+XNuQTSyll
mz7G2XuSmCLieJrq7zip1o/K+1AiCHicZjz3xLckdGBUGKj3vD0AqdoqKWZZNSTLDvC76e451Vut
AJtzGU5qi9OoQRqocCltFSftivlSGO+9cZe5hqg5rBQF9Gks/ZJdAjUeKaGxJlca7V7fLHFlOBDr
2vXdRkYRrmBnnv8whYjdz+qhHL/8//VfJ/GAyTtAPaJ/iZhVETU5F3ir6h7ps8MrNI2ojLnTW7eA
Z5vWQgp7bgnqCwoE4z+1tHPYdcPb5P8oklCau4zhCirwZWP+C8COFtaFDj+zNAZKAm5GG3FeVZ8c
pIVgRROykl1MW9wNDoAeqtwSB2lDUwtXakvve+h/c7+TOyu+RVfSxCSYNzAc08syTqhCl7dnbU9D
p6D7CEImbGgpSlQVYZ5b+oRfVhLhfdRd2/U5GuGtUxX6KXHW9D50kW2/luGq5sGZRBXQHbp2rTim
wcaHLf5F6AT2xK5AJYVTBxylIZ9vrBIqPuV9b9Dx5At85DJbQI0sLbV29WHB+7Vgwv4KvWZ1Vsg7
bfEjoghFUVXfvoPdJj94v5sGul75TMmMMxTrFVXPiN5qF27eESjCCV32mr0XC7qW7RyXdGem6okS
+a2P9G9bMUpZoKWDTnFrJtxI5Oa8eKOLLeu/8j0WJluVsC+MpvrGl5iUMb175nnT6OFXcozMSvDC
FCvr+fI+pyIwdv19Bt/IikKZoyc8T+rVGxt53WE6le68PvaGJOrEdnb8/yBV20KtO11/Zj2eKLOM
kEZKLIaBllwl65SGYaeokTthNZ7Gcj761LzQxc58k9s4qpQyaq1l0O8P+1DctXpM6JmzDj1FQAnH
O2oMvk42qdIGhsaffI/XGgjIDAgqFf1ZfTbJK83joAGtmiMsW9NNhGEfJ+9lvZgyIbQRjMmiwSYk
A4vlqLLt7z1dZPeEeCIRTvxk1RVKSpUqzt/KULZXob5CNqcENta07HXomeaKqTju+DfCLEu/zlgU
LvS7DstiuBIrUXE16kwknis0UEPR5qYTPWZtJ18GI4hvCt5Qmvn4bO4fM64psrIaDYI1ZXK7T1UC
Ic9oULCGdLoqPdQejIA1GTQRvSNnqVl3w3SFXdxsJi0wFmOO4pqxE+nd2ejWmGTfqCj/kxBCNiwn
1FICdaT6Li+X5U0clpKtAFHKU+6NFfbScl9zYwV1Xm9AtsJgRiPk5GrgY4HId3LyM56C1fYW2kbP
0zZIWdzgUhBr8BJG6f931dKhCPwKq1wFCz6LfSUCUwbyecmsidBSoAxDDSvSxIn9+dsmE48WNAv3
PfBr2hAw+nZQNVchEa1FdOeF0SP3U51UnRi80tBseCUQilIQH8OI3BNijX8AXEbqUwaskoP521W4
meeGD8MjwUgeKZFlglw6I/QQWGFqZFQ/D5h/bG5C+T1W5x6J2V6QQBHYkasMBO5hib0Z7O6wD/2l
3t7tppUbNWhEWXO0c7RDozzrcoBvcD5hf9zmtbdOJtvzX3X3Z7/B3gza9nuwTCehoN4gBbTNyVba
aCa2XKO4G/Q0TSp4oa9Pa2JT5bsG0GxCqvn7z5VvWylnYsnZO/KeY9hkdUyzSCSIYPWCsZxneZYe
xDYeL+BrS2mQV8ezYUaIiYJxMtEFzUCuoHetXtfjViyTRtt028TN9z8vcPt35/x2JCdHhUiiLko6
wVHPwwXEknd62Mv2CtNvzd5Pzb7uXAZZEAm/uk7Ef4h5J8Lrmcq87woNnVTzB2oDrbY75GOB9a46
H/NGy306f0aImeoj4kPCYI9Zoarv/N+i5LTJMNbfvZ9M4m1KIPpBkGrJHeHvQYG5tsiTbanskUAg
1uv2ZfjzvvyRVLRokBVgg5u4ajcy6au4q2MCumqsKi49N4e9Pp4V7cvfvNcQA8TtZL5n1VvaSBNq
QH4Ryll6WEZALUzJJ4DGtgi0zRiBHksQuiquiCTblnebzjJhFozRXjRAXiOskvj2I58Fq3C6m7Ci
OkvcIGX31lzcy53+h3plACLg5kJJBwwE2IxGQ7Oq1Wcq5AG06E+zzJKT5W0TVLA7Tj5zgMi3rYWs
9abhxp1qy+gzbQIjEoZjUQofUlGAH0k/pSj1lenEfpZSuNvg+1TZzxbCmWSdwNkqz2wIBm3CL11x
9LEKkH+SWm5l96O/xxPqOYkoRZAVSvfjFrWAnSBesKIIrYq3Sa9/yOgShx/QloiImuxc13YHik7b
IgTYpqSRV2BDY7ZBNfL7gvIpeMtu5+wcVqPBHURoQE5ZU54GF5sCFFKvbqsSK4fDKQNcDCU9wEpF
E/OK/Lkmpx8mXCHxjQ8ExmMQxQvTSp/t/PCB5nDh3wChBAN8tH85aO2k6D6qKyNNsM2HhT7Qu89C
DR2h4Q9GQERi57TXeuTsZ8v+7Y/Yoftm1qHkRB7JqaW4fXDCZw7wPR0Te9jh3wGOPCiftS9Q8hx7
nJblfF+wO2NoMWiAfobog8f7PHEVtwRuB5Z1nLNxlrtTZYUp45cURAh9Ak6v+/880/gwJJq0iue+
1v8s/PAtiJtn4L3wsLpu30I9ze9imppYTaqsfQyZfo5EL9AMxnp6jnFv3Y282CtA49QaIh8WAXHP
afdX8+ZfTSuOX29Da/vM/WzUSe4Ge3G1tzzpmsHrMFTScMbx+gNwsrPJGJJol4Qw3ReulfQTOiTV
UPKg+5y84s+zrFtpr641ZKKq6WA8B2ZXgOvaZfO92XCWf1JiKAkVo1qxjD4mby58qhA4bQ1LkW48
X9QNcy87AvQiDDURnYh3LGNze5BmWWCBxe0/XrcpaPpdwvLckjrSUFusZmqgsDe9lcl8KxUUGTA5
sTiO899evXOCI37XLBYPuELikWjx63Wkt7KjI/NzXYo4+vLxbtbxjqOKziIKgbpzMLp2s0ptarkN
+lsFCFCAAsDatNhYgvgTqkkohgHT8/7PIzdlYYxtK7465M9PLlzMPSN3d/8zE90lJFnrM7IC2k+P
0rrctiMsXpSobaXX5mOCWRlmK0LR3YOk97Xi3DiiMZFSBZXftT7MLYQFzCuvPuWC8Tv2I4EANObk
XkFiHMztvyAz33lwJ3CH2GlisR7e168xd4eEE8yw6be0ruR8J6laUloZsK9PBhtRYftZVlkLQt3m
HW9MNIJ7fq2eGHUBAatx46v/CTuqSRfwNRK4NxVoouGsOEKELCsGAO8aDaVqSvTANGVU5RF9KCOL
NK+kJKsD6290C3NGFGPn4hNg7Fx8GtYF9GpzE1rdyFcMuUr9OALo5knfja5WupUFqORtvtvmQ3nv
tLxniOVTDr+sUApjmZp8vcK2Mp8kSfMEF/bRHonnQlA0m41ciMcv88miOWUM5cKd5Ehnarj6iBc4
yyyf/s7LtDM+LJCloBj0x/E6OxJXMZs5Cs7asogxGh2O45cFU3rTyi9w0dF0TU/UH8yQw4TKFDW3
LcvowYjm38ytfRUcYJ7mqqsVOzkAkSANTWfyzoCDi0Y9kq6RELwUreC00bDnMb/Cu+Dsp8OjZcsX
THsAwQHaeS6O89oXXqMJ2wpMDMb/SD6DQ9aeajelBTRHzpLodvSfHWWtGxevyQu/3QmTkJSkCE8S
CRCx6KGwK9EUquQj6AojgjLi3QnvTL8los+K194OIbOH853nteQnUulsF7hN55j77puu+XOBvKot
yFOn4hib7hT5NW0C8UBNCiIZYyUomKgtsl2MJaoR60rVVT0W2lGUtNhxjfLrvyQck7XZTivyxXcu
t16+ABjBiuPJ9Kw8bAPTCsvvR2SzXodh92pEO9lHWMfh8FtuVxc+JCAEk/VTeaQdFWCLkYv1RlNh
zcbM7gNSfAhnjCF3Fcq3AV4x5ynIUkUqBbL0OVyAtucYlTlQpdVkcugBndC2ZwcSC1FcAzP/Y+AY
LGxpzhYULFgJKzWf9E2+K/k7dhNt6Qp8p3DRU5bDxojg5G5SoovKslowmY+eda5xmGREvGiKewUi
ZDIC04C960W9bSDTuR2GSArxY4dVpPRusKylhY6ecU79fD0w93kTlhJglRWbWfMkdBt3lE8x2p9a
LI92o4WYvxhmJNUScUg6W/HSxJep0FcGOOdi5VFVdbAYOoOCxqpz5wBHqRiOuteqqz+QqUcJkBuh
lGIYENmtmQME7YrFQ9SEfENe1IHrMkB6GymsJfhSgdwye/Lj1Ttds1Lzkrg3Nl+OzlzUbk7Eztg+
2lZoqyfVIptnTHIEqb9WZ9P0axtedg9Y+w2/gKXe401ySHkq430vvf5j3aCnF1DQqWpMUjte2U7B
mm5Zg2UfwUd9F5jwZ6SnRusNkNNPOki2mozDxgoRDG92KKw/Of9CFygOM83uAWxQp/zKsPOW4U3A
ESDmwAjRDxVlHPdswnZHtyQO1juaKeTlcNB4WEVQN21s5TE/oPwuBFD3QrIMU9bTrd25cIb38fJQ
ewyJHVrSIOWd1POcdNh0ESKE3i37ypDfQiZVnpPVYn90uoNIx2e17zSpnP6uR8PlxwcRabSdTvtc
oiqo3BOTtAstDmlzx2sjUuHU4YeEZiKRoMvmfM1K/Hp9bcXZzvmu3kbwe1goa/DxfGMobpQ0coIR
EwNIE7pbbiXLP6F0T2O+36zLAiAViyz0s8YHbGT4EozLO2M5DDS7Ev9lBa4akW4LMu44yZ797Sk7
PJ07K3FcHhEYl+1NDZXIZWWscBl3mYKtkNesZcbrLnIgD3Ot363BZmkXCbI0szKHrxRCdm2UWjC7
4Er3pn2kxgOoi28Zgx9qjKRWQ/onsL4AXR44gTro2hQOpXgcqBqiQOSCnO66xelUe95KctCEaYcB
Lqhj+3fJYpxImBwpVs5yoOgoklvUFIQupqTFrgA9yAv/uxRnCkPS8hzkaBiGxpk6neMwdlK1mzCD
x2w2dWUGz922u6yDHt2sGHuF8uEMBWXdK7S3DBQ0cehx8nt3GZHYOA7JZcMV/VECNSKwYLqoGKAh
asOj9ucvkQ4NuTcZ3S8ZZdaHVZVw2S+JLplinG+R6MdNav2m74Vex+FXckLxccyCNfz6WJgp9rwI
sbLjKkGBGFYfmM5DOY0BYrVkX0/A7TufC/pmp1h5UDygkpnplU9QmXDjZxLhF4tkBwX04pemqs7h
2ZGEYAELxG2LlXSXUWiTOgMp01bQQgVHmlemcmdlbWafwICH9bbrDH2Mx+ul5s+c8qKlqRMWlJjJ
oWBkB7pPZU1t5oiuS0febEwLGjOTgtPAupzTwrHzC4VdM3qoMcRQ2M44IwKjW8CbuFhDp9I5lcem
LK4OcDdOpVaM6yMlYZe1pfOVD2u5yzVvtL9D7VvtkXXEMjy5GfrMLuwiLh+Yo8KRjEx8Eaht+Vmd
LFOz6JaAx/xr4KBS0xzNBqR1PrS1D3KroKoPtiGI7nk2m1Ta3N/urv8iESn9W3x1GGRRVB/iQpvA
DyJiciGC+48X3xUaYfhFtijz4qFqUF2sC3gMREFzBdvQ3gsdKwpYcvMwsVSeNtqhBaN66KlNblZx
xcU8DQ1me5bSbVFQActyZML7peF5/vh64Vtg3IM9OKjh5mv6PMCgJuRcJ9WA8CjUAriv+RD6dBHK
PYA1to3Fpt8RvM8OWOdL/JWc1X9rx2hell4dIQUeKc8Tvc+Ur94M4iP6NSS+P3o+6mBGUir949JE
kUB12X1fo2COFs8XDqgndI+NV8uYdqyStF82RRRS6FPTLUuOcYUlnTaEb1TX70ZYH9a2cytMZXX4
z3rw7t2tJfrOOPNBnTF1AITRdvAqoe9q6oUyUcsjrM6N1WY6ZAWqLjmTTMgZJyB1GYO7CfIs9Mv4
pF9o57Kzr2GN+549heE67o0wa1SirXV8TGyMu3ReI/hBs0rnrfEfenm45+IeIHKzzp66rxUxvLHs
3IoOSYq19/OC79lfx2F/eO1SYWdneSECqd2whDeRC300PBd6Zc/WcUlNZSrOVsRci0yWsGVgyGEW
y6OsVlL2l6m0NEk9mJp/BoV6XSnUxmODn6Vx/II0AOZF6+hC4crsFCeQ/bQf4NEYKybL4pjxMvdl
v35xNtl9RaY0A7wMs3Q+LAqfsJJ5G91kRtD8A5tHmWjQViZH3xgB6y4z8fXiLNPxBF90Bq6ibai9
8TESWDDr9SjaMXuYkI6s16is/KyYel8b76xfx6b2RwcJCQhKMvqCgmLJsHv6ytCd650kG2yG90rn
MtFAfEhM+jEwD6WaUGjZK8mJjw0FjUghn3VZb40SpDaq1fndF0IusSxwlD8STgs9fIHGoM5LNK5P
e/hmiaQAE/66CYYyf7f7tPQzr+vRzlrQy5fMeKaC4AQeL1m+2NUr5Q9MWC/wlhB2bTO+hgbe1UNs
VB+p20jO+eXyBe9AWIDboIj9Fa89l2bBC0xvjGK3Y5e5kkRgdTAZhiE0Er7xbNaOpaQW/NuOLtzm
lB8EnF2lFMwOr0i/mEveXJySJs7WMPw7Zngl4LjcZok1RsvGY+phaNGD3tzSDjwgn0y1hNfEgp+f
jl5Hsa3sbTgZHVAdC7pNJ3TpiJSGL9zy4pp5tZ4AHckCZY2u1602gp5hxbRoy3ghBk/yzwtJ9bzf
G6J4RWkP9rGReX6luplfxSBrYC8fWVD1Rj63s7Sbgt5Mmxsa9NcGLK7xtP+jOe9AtDZjBEGCpT73
/2nenM7KwLqcYsrVwkV+hBTBY4jlCHyJlnT/AnU7t8yAj9p6sg0cj8VSxjyfCrgDK6yq62iZQpyZ
oka+Q9kFRQM+OCTke/AGh/JOlhf5AVyuhGPCe6mwtEO/XsABKPr357D0dUevhiMubVj8aOfzfuuN
G3WFPZKaOx461P5noqTWvYsElio+k0d7q47I4s+lvHwOJ070m9XYX0DwZlIdjtBnIPsfs1MhOl3q
/qnlrbqG6Wcl9fqCGGIPkV2IDj5YdwHHghhjLste8bObWjV29ql6xlpXcquzwG1F7+gnx5LWoePG
LT8Z6UxAhfIAVfm9oiSkFfXXQAyfqr51dwGptFX9JXe+Cvod8+xQ4xo/x0rcIpop0lPOj0pa9V+j
WanBwzzc8EcabSK8KSZFOjCINvwuOgoIpD85b1poSlpQjz1LX1961PXbhPl+P/j8eP5PC/WoWANh
sb3DaJ4vEbAqhikdWA27+F0oZ+gPJJspxKZlUZ7GRP54sDdA8pp7KV2Ma+RDb2keJrof/J3jUOu2
lf7INQKw4XnHsDYXLLXDef77RR/nKClcqo1GIV5avSD/ZFDleH+sCxM2fbj+Bzm263WcgF2lvtng
TAjJtYzAsC0W6dGX9Oay5RCl8OoaeFK0dfdWMFSbqwOkPkIDEYf5vhqpMOlBafj/owMsfafXUpVz
bHp+8+81POvZugJqNmok75s1DoBgPPUmU7garwsQIuu2HuMQJfjpXoSwK7yuHhQu7pSyBPKrWVeO
XWOaqhfg4s1RhJCHFi/LEzb6x7G9EbjXFU8UQV/cTcsu/gte6pOkCx5KtVy1BUSRkUQwinCTyC6+
OvOcuiOwlrMS4ZP5WRdN7ybNUVpLoZmZeqinjGN4YCaCB6qgIhZagS075GnkNwP8Lg6wzvUhPM3E
jiONI/pOFUIbn55HeOvZRJuDyPUVtd23KeovtDoMCQyLqkgr9BG7mZvYydfZG8m3UbqrJWR6N+GF
hP8bW+Yy1PDUZChH81qX5RVM/NNmhHWJ3weDhADm6e/I1mAomdVdQzq11GbvkcM4dRTnyIhUrs2r
3egKJe3OVmRKapjGwW0fIzyEfI9sBz1IBP4VrJ7bVfaIwdspnGrGGVUPT2BJKilQ4qJlQyaxi3aO
pIqnv76CKQFEfK+7QaNlSi3IJRREpTT0QV3SBUMsCtdwfTUzwiDi5GF6QRoNNHIVcY2+Aj7TAl87
XPIjExIWINX/06LA+RjK7hAPYlFDHDWIoti1+86FZvsnKVnOxYXMZ3/+JP2xOu850Hxvmu66/Uig
Uf4+muG9otQGFGP9+yyoJ+Klz7x6Q2HpcqIQcz7hnatNwJL5YT0bh8blq7Xg+HNBT6d8BphO+Y/i
Htf1CtfD0cxX2h2BM7UEfJheCCgja4Rmb6ADJsMz99IcgMtGjTyvLl2e2tXFY9m3kjgixKg/Q6fL
Vyf3ar7oSYDTNub13WuBAh1/lc8FS86dLPKjFLWjnE/e8EcDGmq8x8ezdi500Dr9z+c2+sFMReBm
fwl+FK9V3GGeSSFx/vh6XJ3sUR6N9fbiIzaG0Jh8QfOvKsKARUI/3Fk5KV1W+cJADDRBKs1YecJG
LQ2KwFp684iZZxKKVZdL/OUgq1s2LExxWPT1qzvos43f4yd2WveRGfAsadT4Y7L7vgYsVEWO1td7
Povzk94Su1OR9IH8gRI34YhOBZ8a6NBjYTFSrNCy6y447G4NuzH4l0PCLh9h8aNSsBvquzkkeUxq
RA58mh3cP9Br9D19XoDOIlw6PdT+Ms8ilqHpi4SjSnof9ynH6HwNA9YbT8OU+hBnsJCxjPdKRiNS
PGzEPCKkaBVnS/qLzw6vcXErODvHsAbCLnE7KjdEIgFD2XFCMmlYg1Y3ytuvEhlRRIRGQnr8ByD2
eaCqhurW0Vsj4904woAZ3LhbhoqpaVxVxZGqDBe9bLvPRLT71yeBu9LpC927V+CPepaTsnPrjrEA
WP7huhzHzzsmFuMATHIUHCxdtAgYWXR2AmlQYcBxKY0isaCBmIj6RbLLAmIr0fiQlhr7Tj5rrCuQ
NJg0pHaDGdNxAC1CJ1xi/qkCN6AaUiL0gdHCdajQIm1kLYnik0MPNoOR+0k8OMAHymH59rWWQ/mv
FDdLSaZDJOWtSREx1gPehNq3T7Yj5t1sNz3JNWbc7yaxY7Kp0SZkDY3IhPDKaxMLpc1L4bH+FcHE
mockqUy58u3dleThdcKF/uNmrU7Y0hptO3rTTv8gLvlVWzLjU2ZvY4k3GLTwJpPdikNwzgx5S24+
KXdwf7h3HS7GWOvydTAKo32WZmmpGCr7T4jGZco/AtMJbAGTaS1ktawBEyOz8unOZmsyJxc9z+LQ
Zg4qjs8oc9fwC1De1xPvUeHXi0nM9Wn0gnrXemsIM4DJ79QCOU1v47ndtRRYeBRtgRyUcdls6gwv
+OrNWQuxWr8dzigTzxWk9AxKjGpjvo97SdmpsBxARutKbcwyI1QVuCaja++Bkcy1WgPgnf1yI51P
xaYxEnvd/6/9UMBkZmWxZ7wve01a5ylq+8aZ1mlBlaP/Z9rRdV/TBPDPsvMSol4gmVL1/5RpXmmM
SDoK1oSw98/d+trtf8QXhI0CTyVhb1/2wKnkxV0/or/udoGbPStLWsIqpakJQ1xTH+kB7Y5u45dS
s61Z56GdvUTm3uq40uC36wbJcmw8BL/lCfzfTkTCvUmey6uI7HlTLPXCxt5VsC04cWgbeqcl9B+q
hBWBlvGpL1NgfF2y30EMgDNwUy6y7NMFuJx6jYD+723ywER5IqfjOb6dwWRe6T6VnOwab9o8GJGI
1tqNVkR3XfTr3LEudgAuA6BHkn2aHOnP7FIfkA8ctTwCs0zwTNP/qdjnGZNurjFTQxAmLA0vy+SF
3l3YzbvPwGqsabYNZVgE335RRKLuqdfg9dWfNj6TEleaV19D5JeZWqK8AipdgNo8UmbaUFuFKKlW
rRa4HKwE2aMH7/uLf3VOLKWjhwi+KJJ+kl4+J+V/nMNOs5gHGZdZLR1conaHg/pSat4P8NLRQaPz
B2XqzejkJfxwOmzNAkVEvGDRK0skiQKHhmnyHC3gRhPoJS7FUwAUfJYIOnycA/Kx+1Cs1efJXWF2
Z5YSa+WEJiLnqHQsTV2g1C2/CHg1CmADVQ3jCFQ6SUS3L4BkFxQEZQvheSO3uzxRBaf8zqqvh1WC
2CbmAp5jq5LQfVO3jNoyWecGQ04tysWvhklCP64L+P7RYpvfjut85/us79wlmpAN9ybAkJSOMSQn
Mm45vkhzP/lw+u5xqAx6LOvUsdY9W5wm3Fr7YPUU4aYrYuf4qe4wZD3m16+8jOz9/pw3btZhDx7i
2h1DFBHszVM+cLyMR730YK0HOlxmN2c1AgiiAovHFdcMECCk5bfArED5diidp04RxJCB3NMtxmS2
0TQsVcSuRG+ORG3kIyBqmfAOu2z+ap6AhYaz0WEqkNmMg2OsvjS2oulXXO/1bMOZQYImNBw+59Ph
ebhPSlxWIPDMZcXA/UAY3IAJOWDQ/NVG6fjlMW5bbcGSnirQmQ1gmYy5gJeZS/euBs5FW9ySvPkL
4UCEAup8ng9YVRhXWCeBOA3KGgwOW4nxg8gG0zmzEvsjaIag/JGzjT0Fse6dbWdrlAp+K1BqfJ3W
BHYRiNbT0/e5Uy2asK7GnXY4z3DQ8k2hT29SFuqtxLT7Du4VMHBT2AuY28Mp3d0wbpbqv/kP8oK/
xDRmlq17dPESMlx1sf9HIx1qMNliGQDb485iZe1ShWb0J8TCeUEUJDvLgoxFPTCFUY069LNzI5Np
pnmw+ZOhSGKHgSkRpLfHdo0zrjZOBKKaYdToKs9lrhn2yCBqaVt7vXsTfVOy1qKtJzie/2pNlcY/
YEuQZHozwyjxiWfsPgzGNDLAvHOWnuMSIRVXEjhqcPoBi8VYbXWygbcxlLhgf6Y2J8bxRdunVhqS
OQjnRHotfapLYCpXMQtX/PFtjZ9Ag7g+3dXtSZu1t0hyzkygAf3+cHf8ej389lpb3agwi9Jyph10
eNn79q1hAAZ/0RG2Drx2bPtyEnQiOtKEmTYNfNeULkTU3NSnGf4WFPYbsqAvpXLbigvql9iWXCj5
YFcTkH/88HsQuGQrzDbp4XtHuIMBiOIPwduGesKKAqiT1H9ymyIU5mbqUA0eDMKgSeT7gNVj7ZUM
OXhnh077kQDWE0aIQ4xtyQhgnQGqxOp0GDxuJciy19kd6ECeHlvoyzC3WD96ZB9wjf1qzb5OvPz7
qt38dKupFJjbJ0fuM0WakzEmNN9o6DuiqGefrRRB3b6u8clGRLTsVhfjZpPR7g8e3aNk6QXSnwsA
VxaJm/csMbleHr1DpnzF/qItjav0VXENpmwBvusgiO6bBz8DVSDo26LjKLsoKlAcJ3wW3ME7tJE5
RmcdSyLqCV6GDJYlJCqLw3zjvHteFdBgdTTGsGGV3B9tCdvJrj2qdP2+TUzbe8+RTsXyBO3n05re
KqEamChri59oDrsMHfYW4Te9V5MuQPmInhax+cEn5+8ZsAqF4YwcQUw6FFtDdH4HKM8VUzTAiDLx
T1klO+Jjuj6j3gn46T0pivzmNt2TZn02TqtWKyY+gXSIUQ2yKcoArKGDZglcdzGWe9H4O6cJ2ltu
8gq1w9ZudsK/q73HXxH81dcvNj7XSc30pYrL5OijroQzBfD6TKwPZn69GXV/+pDhShALCy0+WwbZ
B9zXalEIEXS0yu+Fdj49aeTDTf2YQe5BU+ePeIecR36jpV7Pvkz9A9V6TF0qwOMuAj2pfXeurVgm
YZO7PWya+b/wZku6NXSNi/oqXF9C2IaSV6tA7UHKrYEXY9X6C5GEIy+ZzpVOolF6jwH/qN0wlkod
aGAh3kyxP2AwfiGiCLJenvW9ATGwJankAJ/gnxf3sIzpzZYEpWcxzP89FlKyn/P/gX1cNWlAAhiH
UFLxp8YvWT3ea0TQ+IPZ/+FAHGAmam50doZCBoWa0Xj/SD6Aq/zpKnNeiRfK6lGkmjRSTWhUbwjt
mdAJzF01/5cVDqQqaG3mYvZ+Cxz91vVvWU7yEGW5aP0+wyGxYqnCfyJ+eui5v8P1EZ7ri0jVXJjX
2k0lypJZFkQgP48UjQ/sClhGsTsKrPOkHyTdwlEh9yKdr/Qt4cVeSZ6JgKSMMkSSmCzdmtzLzQrl
kJYAJK1U+reOZrN09GFZu+TqZ+f9/I1lYdSPGml/HGV/XbbDPeUG0sGE/VZ6+7wjnbhZ9TifPfu2
RLe0Bp+iPmg27iUMX9jn+uY5QcjyTx+/8yjZnpUexW8P1M5PVd3FAPfn/KbgrbI6v8FH8aI5ax6H
9NZLFo22Ku6c/WuALbwr3IUq4Tt3Og4+joe+ZF3gutN/Oxi/scawW+SUiZ2UmdDxHv7Ed4qXJzUY
RP+OZmcFzPCpSHxSxupoL1qkIOzJoHjMp9lEKRHIk5urjvnXTMBNzYtBL6tNvGnsD/vHmvg8iC4M
m1xVz4dta29MCb6pHSyV9OFECDQ6s1PvM74bdAB6LTVZbleq2O41aMAWqCNEKnTRFWnld5YpMUqw
INQucM5Qgj6llpKtxWI9jNqDTWaeM1716Ov02RzeKffz8ou0ej1byZntTEjjvNakHgdv5VOGDlrC
D2mYl4EJ2YPXs6rRECUbKInLdQc554rDVtsqZ2gn09IaBIPT8TcRZadVQ7nonnuMf+lhxQuclANU
+avSuQV8uXR3WZJyCylkcE35EEMHaohigruyRUHXgwNKZQIgGVyAGvpzIL+S3S7AvEo8TNf6edsQ
maM2xNBDfe2He/im8SYjM+87DBg8iADSf4DzLSLFfPJ17pS5vN5cISfml0qsUZRZv6qnzyLfJf6n
D6zCJfuLmOK3hhsy/S81U71L6+WP0VaM8ByCeG7TNW1NB/sUHIHe+/+aK3q/fIcNzoqWI73VpMvl
aXljxZ+JEtVxaE+5Hsvh0OS1xk80dpK+p1e6TXIx8x93AqAr160cd7+KtYxDXzazLPUgCm5if+kk
71JQ+5NutwJzEIAX8SWZdUkx0i+nyPXQXf3PYeV4Uf8UDZQe+i5oW52w7CtyZhYICc9FTNQNGz4g
9rhesuyXB5hllPa7FutKdItCb4QJu2WSTxlzy1IUn+s9tFepkkB6dFRQkp1Kdy9OxXaKm1e8Pyvy
tj6jcjqUo/2xGwjjOYqOo5KtHrEtKQXO6YzJlrL6zDf1STNaFJ9JoBkW95RjIe4rXPvtBOiWF1UK
fkN1oh4MFrD3dURKVB+Kiu/4XYVRnOS0qcmOcLh03KqpNF+5h1y9q4ZcCtDbbu6b17PJ2zWnbzGP
gl+QB75eP4/x8HjCBykl7fdo066WyKrthJQW98m1H9EihOBCFhhUz7YkxG/n5RkOHDeyqeWoZizt
y7Yxg2daEN/KMb/1LoxGjpJeVshzrc4tb+XeG1CplZPQBPE6TROazu1G5fhniHcHfcZnMLRU7gc3
K7n7HSxpzMUElmQQhkkJ61leLpPo60geXdVPQW8GoM1x0hSnJELisLoTyMN+hiPMZooApBX73/jp
rYWX6lJ8DozdibzY7b8SNUKG0JPfeEluxIyUeWXJlI2IXJUe/cQ9FO1uq++m7cbiOxQTJng5NVZ8
ez0yNKUDO/DeJocCKzBm3fvod1ETNLzJCca9H3vkZ/ebnYXkT7B9gbJrTXLGFGgZdAuj/oAUlcvq
50FL4Iflbh0AWH2nPbosl3egZL41p0dVd7GiD6lTxI2j4tB/1SzHFUXrXt1QZssL2RsXwoXplZy+
a9rscDbiZi0LN1B6MmI9bmKiLOk335DvZ9uayYVzzyIUROOUVqBb2VXH5hQPj7/gvMCnmuORzXK0
XdAFiqV+UBB0oqdgBD0h0N8FOQzIXaE/f4AB+4+dZVp0bDUsSw+qT5PcCpvnyBtOHJcrdlTXnT+R
QxvGscBiaNvC+8uZaiGXE+W1BsXCIqBN/WVVzNAwWlQ3hUpKEzyKx/tRP/l1u8HAHv3zmPzstF9B
9D4WPR4tSIwPZA+YTOtKyyRxtaBVsaVHH/bDo3VSt8CuChCXpqumjbE6vUqkI3zK96xg51uLzqor
47Boal+9eYRZRTu1eD+Y1wZWxOX6qjfirXf1DPgDCgLI3FTenf2QHAp577rt8zPq9AUqdwGd/RTK
fmDl6aD2zkb07KMTuz8NC+UkwM85Xdqfg2rS3tT2EaZBKbOzFLDE3V4ia4YZFzxvxL4S6Yb+nX1U
xrEmFVu5kILho2qyEXdc3gABLCw2rocHdeFc1le3WH7djaEWKpYJL1wQuWnZ63A6qxkdrieM9uOW
DHjmYYw+fJwDkIVRlYevmYi64CnIUREjIJgauQfYdOghiB09DPzTDD8dFT6xpuhUPzcpQC8sm+u1
daqms+Omq98o3H/JJmQl+rZnHyQjTagga0bQDPk4AGxkJn9p6hvgJ/BA21LrfdpIAN8nrCw/5nHs
PELk+d8ZeE9yWMA0RSYCA6hrfgl2kABmZ5CNDqnr4nguHpx4V0CARZxb3Z+PRsevHycvmRAm1YrF
JhEH5u6s8uq/DIzkLjo9tEwxlkyA4tbJbx1ITaxcDiKukyl+p+L6pg3ti+iJymGRqsOn6zhjSbNR
S+LCJrxudKgpA+sC0AgRRNmdBOCM0ynskz8bG8rT1Kwv7goJxhhBg+IBX5n37uTPuYhOsnszUQZp
2GAA0QhTVmOnjYyhzxxNqH4fSJYv7C1618i4tdJSz/lnfLAhMWpLW/qwd7csai0wkpY8XxIAN0gO
/T1Ko4mhl9zT76a66kRRwW/q2AKDhGNLxCi7LBTOK+s5RQH5AqLQVYR2xFIg07v6Rzwk92ApwnwT
jxwIewd9S+cmF6lQaNu+5twJvQB4UP+jBWXxg/QTxNs8vAWZVCvjjDa/AZ7Tmfc/Xs5pzUJ+7501
9PhANRMGKcKFavCfOoTAgPpJr38hq7gsU0yK+Q5CHNnHRUoVux/EKR87jajN5zpNzrJwfgEpykwg
K1m1HGVlwE0p9ZS12rqzbo/o9zWSlMVH52GcLy3meg5KDNZBZEkeKemPPcozU0tyPnM4HnrMN699
BchAe40zqIcy24QIfIE8+MEutNv/519OHG36oUzov+3dW+vanUw5F7ix+kTsJzmfkdrVxdTNRXee
vHtgFgLuPGMjESloRVq4l2mTUybT18w+7qP7IWuvPKyeGlzCwSchHSuMw0AQ7caFdxwpahYDBAkO
nkXSd5WmqQx0YtlO5PWVjZLv2nTqY6lSZxjLqmGwRoWXPrg/Rl9w1/8eCfArn7BdFyHHl+eIxs/s
RmDO59kKvR6f3kk3XaNK8I4MO/HEJpQDzOycqOArbE450MZBw7pcx7jSG8jGRdesO1DzBZXEsOF4
hz46vW7EKimMOP08SNQL+Ex2Zk6vrTDaKPkjlFoot19IUexb6KpHAxWnFuhU9Tao9Smoi82cX6bq
qoLFDc0JwvwNsvNQU6rp3D67xCtqdxZphjb1JV1CMnFfH5fjmTQbc3W6MKld2ik0pqeQ9t+2M3mx
aajHvKCiV4kKMEZn06bJJe94dpZDl+54NCbO2CNmNFaF8zZqHfbj5KupF53Y0t5SRXcfWL3kxPiK
KZEORAz66H64hfubsqFlB3owNRW5k5cMo338l5ayGAQ2btYnhYcb+9diUy98pnCkCNyCLeVeHHrT
iFFbMrQzdfoKUK3Z5R5L9LH7z9ZjhONRZcysVCx8+4ZHKc+6Cs46NC7b/RlWKvtCRr5a3xpX2pPF
mklilJ9ij/I+yv4nWyTi6Kho0z85rNxsP+cm9aYh1EKRphhmejKt4RdZDAE1K7jPXr6V8YjDR32k
O/p5EdjRrpDbZujEpAkEOqiTYIPNPqv7Whnd0pWW9XTiV584+eFOR20q7OpgUVxD2FDbi4c0s2y+
U/f6CGXojqAiottC9ggJT0tvM0SL8uInEevY5tMIC/hvigVf3KdnDLRHefXh22olDt7pDYXSrBsI
PO7vYgfBy+V+JjjWsGzJLzaTLl2pNiEgAPmIPQk1uR12AXKVjmy7MSYLlBy+lEY6waBlBvRNCz8+
lVr8IWDcVdLPSiOWjFDH3nGi35F9cXacbWvKaU4nE+gXqiDLM+c/L449t5ob8LPA3Ka2a7PJSNmk
5sZCJ+SWMBQW2Oh3zIjRukwPEaHpLn00yd/4wRdfgQM5tgnnqjjwrUZFQ2Wzmmkh8WaW/3+hG2nV
nL7Kv0hc8Fwg0H2SoPMyI4c3YB+3fGgwf88SAO9Jt6RvKlNMhlMy+jsM+dFdxolo+VgCVZ3PTwrT
TYwvTzDIPpAGfYIsMtppPivzHwmTIb8+R3Wfgwd1g3Xb5M8nC67gCaEii2U9KXZULg5j4nlrhIrF
doZlD+6gkkDC2fZHfxBFTKrv1tjJdw9o7ZN9GIBG9GF2ySQkZMQfpIjPnvxQuFXq4ps5HZJvLPzQ
oP5dkvy44cr5ITVWsVIaTcRnBIxvS64OguJRrYp2xd4qcaTLeuvkBxnvzmpzzcleTTXylmMkKFQT
7/LNRYoP3QswvgFHeyOB5OwJNSgMwc/tH0XcHGNIheqDBZIcqprj43CI1w8pKCJX4EzJDzHHki0M
kIXKL5w1YEGCuB0vwnTOBJGya3L9EqlahbV3GIVHYY3VNko1+ApGmjdJQtz62mm/tpVsYEdrR+3g
+0fR938Y7baiKAf5wnxoMXNefY6HQChJL8pHt4+x3K1IlWpLdvXsAsqtv7fwNu6FDTX6zoFOJayA
YB1IjVMq233o43pMH1XsBhWWZZAL1fYa9+il4TtHF5hAK7z7ZFAzO+kxVspMpJOEmMnPN8H3IFzv
fgMV3kQQXcyDUeCVGvi5SZXcQTVArNWMGwwgPYWk5CE2FNxvkI/SRoLB10I15PNgWl1K/BJHaWWn
Om9AW+P5y9durps/AEOZC8B5Mvmtphl0fVbpFyJGK+x3i2EI4a+n2CYBRbTa/HxPe/veL+1QPV6y
/5rYIfUPYr/7pruVkVsEckdsNmn53uUk3LS1X6x6HdV272HrOnAWqYxZg6nzNszuU7leiI09BkIc
+QzDyNJaTFYqkil7UkzGCqo/nNBuiIwfeuPDljXwWQ+F1p4CKfD8pfrTSWytu7bOqLhyei/D9iZL
z/gvFEuaSSNyUcUpleGXEQKHyx8Z+NU/vGbaWJ2WiJP44gPevB+2hqd3zp+oN7NgXs090jtmo/EO
sF+XkovXmUtDswGNXKqN0LdZKfBiJWeCD2E5VhN30GSU+ACXHSQRE+gTclFwBl6132+bUNRHp50W
72FxPz3ZA8KjN1z1PdD8FLke/Wnq2yZtwtlXucMx4u8v11Ixbha5D26iyKo+MMUoWza8WBPfoDK8
VY+iFWC7Nz11RuvO46T1fLgDCdivpaGb1ccbyW04a8Gs3ZuL0DsVpsuCCFFDOmtyehAD4LIx8f5D
XHRYmaGh4/TDhPiTQZnZoAt/5LHGe2jKBaifRkS9tvFnzYt3OS1Pc7ZONa1+Y4mybdY1Ggkw3b9C
cbyFupMlrUshEvwWF+Q5hDcLB7qxMAvdMl3ZdZB6fhIH4yQRibeT04PeFwoxp2uSj4c9uDH+hk5W
IeWl/gtzwX5kc15AEXYrtF/O4m9WyFb5ro4UlYbbYmytcTbu123OPrlYepPGAxXVPjju7IgPESMf
p4fvDaxqnVMEctwSo2DJDBDArZivwLBf0TiUAdVOOxEzNBYezO2sv7iZ6ilDXgqRhcQukmIVc+Be
l1JSFK+5UAh+d2nJGbIWxM4KAcJA1wigANA1aa1kEoY3DhipeAkovv8j0cCatdRzqg1fIVmcK59/
84NjFTerAdAY7QapJ9zs+z3cEh0t4+NM8iuEUtIM3+Iu/oEHfxX5W4J01bwndmzSYVCFO6qk811j
BPBOlpC+0KuzCwcofUEMMXBZeUo5LvL855tINUQn2Fg9zf7zy8VECnCJ2ZneRHH2VHmY5Urtz5un
4t1Cq0KKOP7X/YUSbPHlUIWAjzX9M4+drQHIGm/UoQBm3HtFD8XkT0U3s+Bs/ZVhHddiFC3OxJgu
dwRdnt8aMybKnZbNVoktzA2sA+MXnpce+J5I8SQQyRbVYXYawIUZUHFdXgzVlTF7JASHmMXW5RHQ
Fp1mYVmnU+FcYvV/yuWK7RL4mvGacn8Bm2Ny/ql6RbcQfcxHv9/BXWxa4uBKDe1cW2izupCnldlf
784ASoK1sP/HkyWDXSGe1p9CRZX2KoO8We1GbqnyydIIv4Z9wnlwXELuJX53yDxFW3dm94JDwRZ3
IiKVFTTAxtljDqUeWHylyNhW9WR6c0FttorawQ4pujreS8AmXymQiFJaiDp+PXgEgVZVDgH6XFPD
JoIqzeYjJu+huw0+dAsA6Y153QYJuArSDzf6BWbWwM9nln3x3+MD97OBZ8ne1ov6JNL8i83eSjzj
Y6Q8EAe6bFz3q8FNRreeobqdYsj2j7fnHLjTPldWx8rQvQGd+i3qAiFO5HRFQOgy5guqvfe05C1v
rt2GKFNyQ1ahKmFnxo3DD8E698wyM+dwlKbdHwoGt3xIxe0ivDph5O7euc0ahghn7WE6Xcf4LbfJ
Wkd9yieRQDSEuWxVt20cAo/FVlIQ07dd+xmA/xefRZUoaas2x3D0v1u+9Yx9iqpxFhw0ansrO1ni
mfA563df07LlFwkjUlTkdtUrGpOw40b3UvovrhrCgSS789LFpbowBomtHSKYxlzgA3bRhT4dUQ3+
0Z/agzukj3u7m6SHYchfD4m0KIT4frXGpCOKcf2Ch+0e0Wr3Se6yoYQoaXgSercIH+Mk5Wb666Kz
PBwTqs5Hj+2PWyomvkV2cTb+/FB0SOaSED6FrtLK6ypg3IgAsEtZcVRlaVPk7zrbf7NLREzKFFlZ
al1hAAKFvN1EkAYpPHKK+ficPTF8FEvtaU53oO0hFfp4+531cxpLWx0sqCGSU99UO25U4vSV6ErH
1a9oNPnSAxRuWzzQvSHC0pXH85ZfEbMTM5DTtc1GCc7Hlab5UKPVlRsG48X2F5+4qQ+2OgofN9I8
YjBnkOhBjVXsn28bUCcZRhtmOxP2bX8SaGfIL5X1m9HHHmtoj9nSuC6eqoCDi+wlh5Yn1514ORdO
IaTg3CNfiuD5wXUveGymjzNBgV6Pu8A4tO+2+xJ4TxYBA8vHMQEBHtDGNRFlUon7+HyGi5AG3rWO
FqgJSPfZTIwRCQgslht424LLrZGMM5QpJiZUCL/T5Uk23AFBgbI/Ec863Utz3WeuDStkfv/6mVYl
uu66A6DtJhZ4D7Pj84m1IKczwKEpm3Ogs7BFy0xmIlLiqlmcEoek/jZvT43vEL4KmMc1RCr3/LoC
pcyyTdvZwaFFDQGfKm8BDYXniyX6RKayeQZ9biBZHqJfclWQ3sko3YsrrhpCB3pW6cgcZILhyVdg
fUxXEsio4yf/d6JTRakFswS2imW2ooTMUZIN7HkooSENP2GWNUUlHNVBt134Y0TYfkIcU2OecZxx
V8IYbvj0HCebe/QCWdtLzxxrj82443lYpr+8LHjClqldsy0dvMeBZ/y/ZOK9400fFYBdpZ5vacZr
aeoZM0iEwpfECjjfTpW1ON5YeG1ah0o8n2MciVhkrZ+K7jPKXGPHL11dtKnfQ6eKaKtpN1jXHfVb
VsjI2+bzyV38Z12yKsLTTVBmW50KQK5iLi8ikveIaYE6Ds2AEs3YzApqD6ioWIV+SWX6TSgyMupZ
SrA0lUJYVzRPdV15x+Fo7R8SjK2Sh56gZ+QRjyhNWn4rwZ2ElGG/1muTlnFm4EC5U0PEZ5nmW2UL
gaqbpzJyen8cbJYMTU0GJhSHz46mA6HyIB4cyeUWeAwC0FdI1bxLWyu09d4Uk0+5Ewv31U7bep7a
nbA6s7gTXL8GY3p+vheIAWGTy7e3a41XUQrstsRKD5eanYgdMMR5o8kPa7u2kF4fk+d1/br5dzxb
9cp7ixAFWxxXzJvuGYHH8O5lT+xR4iTQYSXRObdbDQbEYCT6P8QyRJyZEG0ZPrIUGJM+JtmKPOT3
UXxlRZcXYItz8Kc2+GH55DAoQAr8A7y4UwNvgt3Q/SHoYX2elpBHnU5tlJ8n6bD9Fzbxw+0YW+Rg
fyR9vX8wnj8iCLA2V5T3DZlyE8u6v3Sy2RfQjfA4+uXoKExBfyyQ2unNuCu2vC3bGkDP5pB572QI
WyV9e81KQKLuse+kok+YVzUaklacaDWnWmOwv9Iw+dtUHaEETyYtNZCIbpho1zYJI13x639VRWYM
AT9oCkiyKLdgoPI3g4zLKfMomqxY6Gnau8/g8RJqLIOiohLlUF4dsQOkKZr4k7rBfTX1SMFnhdsv
8ukb0XdLMTNw7ipDHgJVAB5BQ6/OMGhphxXlHOwoczIsQWTdfDlj1eGZJrqyp0uba1BG0vE7FXnh
n9DGP51NeMuxhAq56e8Ym9zsnGz8pQXBfNOo8/wQxFrUI5mzl8eMqgp+XVnvLGdt5qBQ9wbtfUQ/
U+Y+hEpESLfdNP65qZq/DB/ezHFS3/8I9qOjOzjQSCSgCMVSwGvi8D8wTrGa7X0T77ATi8TpNpVe
YYrU8QlnM/MWcQy0aGfObRJnlJxWnDKx/s01arz4q8ySzpYg/BdahZVD97sFkOhBktvqQ6VXljkk
xOETYsBMnegwBUb8jtC2Y3+QQYGXxj9tE4IduBoXf5Cb5ckPuvzZMT1XUzTSmmOgnQ5JnJMNysiH
hhHxSc2xx/LuZfglh1Or/T/8E0lkfvv68oDERR6Rf7m95lz4rpjWiTJ7qUy62GDuLH7kaZgXi7/W
08Y09ztXLej9t4CtHYxMWvtoiHE/hRoNUyBVFmIstUk1VxaCx/6v3zx3qmd0flx8sC8D1+LZ6Tb1
E+FrLuCOvgWvE+TY+DcYbhX2jfjTxonQz6WpDj3dvZizBA128PoMYoGqe5YM9b/1faf84eKhrwR+
fkOFDjCliLBDqFdsg3Os+qjm/obFkCKbwS3ZZkxQBujrN4dXE9uPfmW3YUlK4jllzNRnTE7FWscZ
xw2Oo/B1AG0Rx90xzrig4odZVJYisGpaLPjVCEMgD8StKph/Ii/Hlvmi0MLZMJ18WdDtzZjX4vnf
0KeAvJ0aeEQyjGP8Z4ZxddtdZyJsVNtCajnYEbSVWqi+JTbbzmE3SRwlMZdbi8JmMZybPSYPHgoK
uWV/ei5IYXh9EKvCnP3zp6kFa/agiXbEhroVw77rJCkbNRSA8sErM0ru2jhaYQrO88H+/cPaJ+5L
Tlu+bbBtGaLLGP4TNaxdXfxqK5abYyHWaJI9ebyvjosBcU201BYi0lQ4uVf2lN6fwJpn/cc7Kv0S
Gz3ToW6CFPL233H8wtoxfRHWsV3RZN9GKXeZVnxnZpyAhadKZlRyBz4Qf66n2BAXgJNs1fcWORKU
hcBYmszMXwvU+Shh7EVXpN1HAE6psZHwbThNbmN7a/4A1XDSsDITnm5TnpVl/fc6eQmYInRiyJEB
LbcmoLY22VOIBqHXr+T09YS22+3k/LeGPc7TrW6oPEGtmQM7rJTP4ZPDbB4JfOAmtC3gLo20aC6F
JBIhPHY1M1S/sy77U6sDjTxZfmkIQSACfswVgDwOIA24jwncpcTBTSaqc5bns9Oy8CFHWj5SHjKa
1wvR6rJIxNH3bgT+cW0+sbcfHftSafb4H4JiFR96Kgs/DqNnCd8CFWZ1tMk30DpjXFUxL+H062RL
mKfvo4toigBZiV6aKCuAH8wQ+badwYtwseha/lNQMY4ntMApcATAxtr8BuaMjsOdh9X3svTeYYzb
14IU3g4kZhCd8rh75byyVifMsZihY+5htA/AuMxFQt7ZXSOtKlYaqnHzMl2+nG8bt6Xeb6LRYPjM
KeL3drc8VRqS7C9ZA1rD/4dpZwG7tt/04N9MYNoY5sotlhze8ISmaMTGevZxOY30RoSa30XYFyVh
fN+BBYxn068DHq54Vi2YG6Onz269qRnJDPj7D6nE1rrZ8pgc2h9HsSonCd/ygpg0a5ZO+ld1JK3K
HLgjknEwpMoikqEHa4SqOVUaNfXZpwIBuFX5bTVzGj7rl3N65SjDU+kyzR37zttS9ZTFlC1B7v2d
gfObdJ5k474NOmb4U5nBZTw4/H9waRB/qTPqgs5J03OUhVqoMjB23UK4imrev+vIAmr0JQYaEdoH
3/JN8VYzMkyTTmlJeVoLE3sVwCIVynAxvSuAECH6ZFDPt+3eDluhAgz1Es89ZcJWfwTQE0gvqQyq
oxAFHqT0R4SCY16+ekEueUx/Yf2sLYl2TmCZUt5RQjq1F7PWAsaZjmSBx6krpf7SMTGDiZ/eoiRI
GyAja1HnyAtq5wgHPTHspD8E/+dUTcOnlkQlqdPsGtqw3UJeVs9O/HXqfFPl3OeXIl/dcNPy+CqT
AkXjx0920ck56aW2+IdAVQj5GXjpzCbBS9QBYzMQxBScdAe/2pwsxo6JKn0inXDGqQWpcy+GFfMQ
KfZ7boCebld2UXuMNCFd9bDhx485P7xM1OCHxLP1uuU4558arBKH52Ig9XKPmLdqpo2AGdbJeRXy
t1ZRM5BfCxULouB9nUk+duwHUHwnN510epMzOegi5WrAuvZ/zfdurie/bbWZWdNmITrJSLd5KNFq
093ZLU/202om/3HI8pdOc3fkyikshE/rY2HX8h4kzO1R30HEHiC/iTBoLzgL+VtMfNAV2SoYCELE
0viySARtD3MzKgwuizBbwhPFVP5P/1LjDnUFtsTkBSgTnjdzrB4+wb/javhgx8F2Ht01OzSXO9tk
6VZWDwFL3W1sbR5PnTfmj7U4urAbgqxyap6DXWtuSlOFqggrTiu9YLXL8QhVTSHvpjKwajcRwA0c
hZAy+yinZycOiAt7FqhnzcSb9t6Za/GtfpOHOgkV0yTEvAVs05Jq3/BGTib9qJtM36vRyiRe4R9m
8L62oiGGySI3tYoBwczTndvsAoEPxXgqcH14LpLdGk4648rNqrbD1XTtLbygW6QQgXKmFUfnLXVT
Rfjhe0u43r/8yscOxY7GWFiDrhMQ/ntoVsXMTIcncmpYiAEyNCJoAu2nIseIp3zczhSLf6A8YaV7
oRwJlKsfeA/ihoPud64WjGNt+MHX9zUqRB/ilbF+bDQwA7ifWr9v161y7xPLk8bwlpZXlkMEZBPc
8PxwZgYgPwvhngBQeMjR7Fn5DSLuQwH8xP1mpdP/CA+KaFByceGkm+Ip8S3AzPRoh5Cnr0Qd2pc7
umWljHpBxgi0+lNE+t5wsyq3qlkwSPtcRcxDJ2p1MDAAHiz9Egs+XuFYdwa8QbltgH1NeCJeNLB8
Pd4IFSXcexqi+mSwV8mjTtU7xrla/IiB3lpQTTWe9Sa9CYa9vIOO6Q6BqIiQgBP0Jfp/Yi5QwmBg
qzycjVLdWNf6zATPP5uS13HMekMM68ZTdAY/NZF/OQYyuedWqjNAbrn4+5SC7AwJYrYmB7KHBDFg
oKbOuMMty/ClwfGzAfpcBrzDuDzgb1IjLy5SEFv542cAvFfcehxCmeD9LY8FWuF5g8qEH+fp52xO
t0+fh4h8MDVJ++yPYZQT9g4f9sCKRLF/5vdamaGBot4Iw9GvNloDY2N2QAtWkLuACRhHEASZ1aBF
rASUVz5OWIwzEz13YPJZ0FM6QEdV+Bz4yvMfRu43A6vauV3Xe0t+N/0tcKwhUMvhwElTmnEwQT5S
5NMyx/GuDoUpaStisbESz+MV5OJhLSnMoSbrggLHywjcpuJsNgsKMk48ZSFeiRR4gURmND+08PRf
dWPe+QcJ9XLhqQ0Bf0UOQFJZFD1BvfDdbnt89PZLY/YztOYFrtloCWfnjcpsvTnlCikWsR1W9kLd
ulsIALUHcUWc1DfO2QaFr5qC8IrwM8d5omENPLmdk3SJmVGX+ZfBr/tm3lF4ta0iav6mu4kdk+Qd
Irl2z60wC+MB7ev5YJh+2DWcbeqkX7WedlWFXXqRuz+UjuLa+f0iQDH1QTYIQaFyKHQ/rD2XXmbf
SwFzCf7ce0f5GBqQJ/MBqrGL8a24Lv6NLc+E0PQAAjLn6OCUQkgDQiEvwCGcYW+Xm2MEf7bfX11S
CzBpPhr7KN+lMvvN/4LTHbvVf1UFXIXjXy3d8w9JQiPJmUU4eNWluOdqxelUqARwtfuRNBhR3EdS
X43guirXAx8srpdeYl3LBa9FqO+t4LQzFkbPrJNl22PYMhzN/IXN30hk0okaLgl9FWf9kG8X5pyB
bww7ja7APuJLCUEWTOmBCeCsU8xnxale7ewG2uPbwmdAdiWxIc620dqCnBsuiA2YmPC+YZF72584
wPo/6GipUz6liryNIOsUmjRIa4QB0JFZeVIQK4wM5c5G463H135bxzdbLtFAs2YDnxll4/5veU/h
dsLWCO4hIWhW1j5AA+y2nZMIvFjd2Albn9PUHvCD7q20sLFo+Fa3lVzkeydC35HnEAvzMUwRLmii
JldcvjpbDTl7AZtPWtnoTpk9A34TLm1bjUq4bB62Cjf3l5Kv7kt824Y7M7Jb/uHIumNrYOr4yCD8
KWSQ8PBMIvwZa0ORwE/DA1Tj0J+gYq5Vhto1WVwbRgg0IKwUaTB/BuNd6P8kXSIs+LfjMDJI6Fhu
vuzS/+sFys7MNV3VY4UG+SO0kFPVMSmjoytA68HGmcoJLK+/c8rJXgBHfN2JIVgHNHZPW5t7Qn97
IU3DKLCauGLkK1XbNczt3OKg5NzZ4DZLnxW9n3q+O2Ex/PvbMTnjJKgRtmBVRJnajaRMGFsRmTGc
2J5nJTkyQfxeJ3iiWCcV8QvAp7Yfydgq0QPzS0xC37OeeTSJ1WZDKJhIj9Oei2oVrjys7Wm2cmUx
Yy7m8NSrXpNvGVqGDK8qv64ikroaEfJERkMRabp3cN1nkaSDtSFAbtNhTLcJPUsU9fvTMsYu9jmf
iAENBC3lrxcIINY2NkWZw3lY0axa7u/Y9WhNks27hE9ec1u150JLfiy/Pf/UuffcwZoe5upmOX/X
0qPVEdtMw0i6He0PhwWvPwuGivyw0aJhbBAen9ohEYS2R0x6NdocMtxo0LY+f2RWsARJCgPTh/Jz
XAqwunOmXsx3UXtFvV8ot6rMs+8zCAv+F7LkotAEv631/sdmzEhOrD3aw79M5MMHWaSLO/+CJqqK
gsCuIJa92rfqhOSdRrdmA5kvKfrleQXCyUdM5gVPjAtGI2Sky1dDPBe0EFzpqu5wGXAktNSfyieQ
+vKO+hbgdkVFWwwJZCuMjq1OGGknTcAxnOCNziDSy8J6RLp+fNnykg/cnxZh0v8BijKG4F70UcRn
mI+o2WmxHW7FMXwqBeBZP8M/+DWAfmVKodpVrs11xVr3hvAr4CuOO84q5Ved+0Bo7IUZWmYSZipd
SlvIQD1wZyavYuFhtrlQObRsOTSajjlXYw8bq9APsfZFtfQG/tn03DS00E3xJOCbfOLbderMM9cW
29lC7w2XsWzuYBw5pA0Qrw3eGOntmtEA5LvoJoIgmC+cAWR12Mugzp0WjiQiIa/cx//2NkfV/ayj
r/WMJndMLaOVz6NrG1WvwlDiPvXlKUsshH79TrFh9bM7+d3tuvB7Sl9gISXI7YIrKpRVDCEyTLOR
ZG8WWQnSqMEl/BC+FgdleC3Ai5uFMbfUL5mLMIQI2zN6oDl/QBZk7x6Lx9bmbadonzb7hNtTGZti
R+5Seraxxf8xXZQqT2dx2YI7ygkcJAtd1+03Uiq/bDszIJWzLnEMx75XBTeZ12+tSJScYqINB/kp
gKIdXx7sl66YdEL2xC5JqdIL5C+Ly8tIwf6Or5lIKuMOAxo06PnTNXk26cD5cQxPtMGkQA+Zi/gI
FzrtBkWZEo9tpe35BbgdF+D4RJasLTVNMV5Wd6HD+q9NNAZozLFhKzjq8gGqIQcJ0ZRWgmlGnvme
vSBUPBYNSSod117f5ld34+q7l4uxQmmfZfdttf9qTxgOXyUUspdmLnWTWEo4QAyZLYakh+FL6dQA
YbZmgENWordCX40eKM4aRanenwfBl5GXD0KiJ6x/Da6e9tITxh4V+XZmLbHspEp9Eab3TylnL4Tm
XkoGDo2D42w82JfZvuFdF9/CY2/436H6LnsF3Qu6DwJoCP1nBYZ4ymURnilDG85NM5vAjzQePqob
4nM8r9NwhvlbNJthfDh0OBQPT0J9oe1u9fYst9NA8nFXbhVMqq/z608fK/NMd9eEp7n7fMe69F6A
hD3SXdz5PxsjTZOzpMqJsiAJxE/KFVTwsQTVHARftCyy5LXsvCcFO12aMIRy9DfdzS8A4mHeFExS
aQdiimYtSfEcFmgq+v5AMN+HvFXIWL58gAvDz9VFVe2Y03/f3YhdVRJi9HqzAbYwSOu+60FVPEqQ
bs4QR8pmXASbDrqTtSIfyaLD6LG2KyawJWFd3DZvzcsuVz6PaucULpVBZmSjq02+hu3unQbutyLM
ZmCM3OgN+brxn1wRaBRVW/IMjBP8FUKFt3m9Tr09Btk1B0Ex0MsEmL8DSNaL7sxrQKiuABVhpWFJ
RdsiOb672FNwiWaD0Z2+X4lqqe2E3op708iWlKJEFInWYUfrxXeAH2AIWTRN1B/Ydy77P9MR7Co/
pjUOiPhlR1jkXmK602GltHDYWw2PesCKoD/hk9cxAwWDU0f3XMrKdSvKHljqBsGpnsErPi2IyFSa
ekzJ0f0ZUMgVZByz/vq4JerFGqUKGCnfp+eMJ9xOziHjyGaGhlzFh8i7yyn0ZwSxz8xBjLKiJig2
46j9dT32He6xrNGnu2JWxABo0J+xPmu72x5S3VI+tFHOy31q1yNHJMfIwKOCcshW2q+AbUm1wHWQ
wQ2EQRJjnq8G2AI0z7Sq2Lbw7qTafxWqyyLae5xpeAiO2P0I6D/A+Y7XqHIjbN3iJ2mSPLxkjWwN
uBW6dDhU3HrKo1PfTkgptRr0zF8ur8pm+SVH6sFSS1aTBNcGSkuhgnLhUE+JD/pVzKEjCMzIuNdO
qtfd+DYi3by0pFbNUQ6h4OLTJEeYXQmvIBSRITkcXrusNoMVEJeLPLAuaMVB0KkkU6tkvBLlUgWF
BMI/7GlV2rtxq8AFMJs9pDMU61X92SogWdfDOZCNBd9LITnmFp5d0ylDHRcIMPN3CAOxDGRGXGm8
ekELUekb5eBVpM0oA3oscbk3hL6c9yw8ol87UnlwCzutIIpF2sUaklbcOELN2Bs2hGLno3bvKQvF
PW0ns/Dox6uwbBhH7qR4FNh7dvKkMK6/fuc7+dj9HMJAWy2K1v+Z7H41vyazOf4XmBilA29UqfcF
B5z/AHQ6vX7cVLfCuiXlcUvi/nVhpIq7awgAnkWf4+aO9Wd9lm0KhPklzKANHY5ClqVeuvxSBFNf
fRI2z4P4KJgquCMn+gF7mXjyK4imx3ESxy937cD4mLq1Wqj1U3/1oTaCvE4fcmMpPxB2j7KnpIiO
OXeQ/6nPad2OkVx7wqv4/NKRz9Kl0I3/mxISlvLQukQ0aq75gK8fAQjfXgjoJ51MrSDdY1pC9Dss
LsJhDknRy2T1amVRhR+8E8JrP1ptLF9dUzruNWZIfE+lm2brdfb0j1Ihd+FpFsUp20yGvoHyrQel
Qxvxkuyj9aXDqkgwjbIHWatQyuy2TtTffxKco1N/y13wBKtFbt5wJO3TeEc8yMd9KpaxmXu7YitM
bD6RH8nZ535xlWymZjiCpHjQ4bI00v8culIkK2jv/E2zHhPvfTd7Mk+EjQHyJUsMHTgOUYCHfxEJ
b5V6ULp+CENWttYGLRjWx9QKLQFowch8vtkUU+0fB0bmgsoklWtv+Y+VDyUDJlTqS2UBze/H4YPa
mzqvYUp3FfP6qHXdEbEdDyo7pm6WvFcJKrXhHOOqGDnbIp5AhcUzvFsbuUr+aEOM1I30ak5w6g95
SypPjECqb09o9uhHHv/NWq0htJsKSANSIqepKCVJPX5RiCHYi3HXl2X+eHfBTq23J18vjEVhbdes
GwmbTrqGXj1Tx3T6UyX+fPxD3OHFnLtwQd9WdMwngumSlMoROQF6c6+V3knxd4PXr60ycOPinku9
G+6RxXP7ETETrHbmbJVKTxjiFVTBZ1hOn5W7wrDZstX6VFe4F+0PFfgxHKrCJwZ1myPTOjsUPDwF
dHu4yZCjR+MlY13fN58N0m0o5MokgcECcq4saJsyc/WHePUYuCbDUGVIDHgiK6pnp55T22npGBvB
oFI5cYUNHGLR5MV1Cevs4cTTmUSvDncG4hQ43ycs4sFcSVBuBVwDlB5WVYUPrG4ZChcML6et3vG3
getLrMeIXws6OoX7dY3k7Mr6LZI6g4WSgt9jj98+3elD/VzatxuEDDYi5s6v7zb6zIwQ8zGbmVUS
gBaMQC3JcQP0p7HUrVNZCpdhKbjuxMhOmwO09oKydGehQ7NtQomom4ZNrbugz4kwucOubsPf+NWy
wDsyXIeS2KOo2P2i/93sYW8njFV4Kew3VwIkP1er5RQwb6REtI/inZmusWU6oakHKYYJ/B0LTUqu
x28jp+PWTDNUY9+IDq/7SOpT64vm/Et1IOUtZv7DoH6sBPmOp+NGrufhjv2lWmqHdQ820VkkiOdp
Ij64FOk1v7OC3SdOTWgUWUcb5kd+M2TuK3CCx4Len7zJc2iTdIB3Th0fs3pTFuf1tiaDLdyFYorC
mSdGvr7N8c5aNPzPcKwdJiv9ZLOpJfx5t/ZxBgitZlcIlM10Ae9KDW9zrezUUViROTxLIfiaw/Qs
sqwBdkQ+yt56xkYJKekoadkFijpfoDroI4h4pvJEXFxcKc/KcsK5oxkvQYIk1vpIsxdZpjw6eleh
bL4YqbsyOYs9ljVTchrKd7CVSGkkxJI7GkP3qq1FUVAIew289qWOjcIu4qJEdLgSOAzy76pb4dbt
+XHSNWmNClPQmTwY/PcsoZmgx8rPpgSOnvS4l57B4I3DU9Ol27L4nD9vU6s5OQ3JAOO+oQ+9C0NS
4L+Tg+tzr3F6bkoLIHNJKQhQExke/kGgMpcgz8/+fZNg5TI8VNMNZahhPhD1tLeOf9oaHAcTOM2D
5E9rkZ8DVAC3Gq+zzu+qTOQd2hqijRbz0K2dC3//cJxibUwAFefBuzKvSw2kzhQ9/DTgRy0BiUmZ
OqWO1Z1aFDxz/0g+IcxCFITWPQ/gf49bP7hDsTu4hmEhAWRYAt402lzBM5Ndpm61SAN9leg3mGZr
FwagOC0etZo55HqAJ/DRj744RNmopE7NtCYQ2bvKxKapqkGrI6X0ZG++JIuwuaQg1hUwVPyyaRPj
CEZLi33Xm0+ZTHAmUO8UW0mIzihVe6/Hhfpy41EqyDEw/howLq6jjUSixrYwvnO8pshiZc6R3qTT
3y8MmT4oKL1x2ZR2nNdnqOIyEjwcBEaZStexLw2fw9aGh3H+mjjVo8XJWLdgqt/9P5jDe9mjVTuK
7Z64AGqc1pq0nQnhhVgoXzt9oqIx79OGU0C+r54BvvqMfMgSQ+ejqbg8hQekH/5FO+TunfbnZyNb
KuGdaSoG7L33OeVdLhhFiRka+MFPiJv1vlBQ9Vcbc9yC6RBONEzaj9VH0PfrTgPI4hmae4Ptv/I6
svH+ajq0zlvihEcZO8zrHSV5To5LfyE+TeADlyeTLmO7t5n1sxFsBv8PpVVcbD5aRkUPpn0e9cRR
eabt4yzdsRu8nreMPkmZETweuvgSYIWVhn+3KW/tvIjoi5z97VkZcjO4GVPVa1h3Hxu1nMrG+HFH
22n3SOFFf4LW+ZVRpUF9TLqaWDUkFsYKe5WlrH8ql7TnK6UL/uKWs7fW2QjicsCD/tObGtgyMtHU
6DLyPlWTOXMgM+37YfmQvp4Ml0KXh3BtwbFBzYq07oh0hJxAXKBckSDTLDQNmaC387XRfQUu48Oq
eSt7QcjEht16IHK19zX8sgiiuc+1jIIAqvgvnw4Yo0rehIimsmqoO1cuYTbOz0QDyDsSHCORkb3Z
4QaidkHOwGdr4vJQ1KGgWA9DA+34xZl3/KQv/0sWDLTanMPgYv7ZlO7wRLyRNksfBYz6I9Z8/Zh2
Amifdl7zt6+u40eKNfT0i+UBlasTvMG/cihLGypjLSgrHkYfJsVjjs++8yAt6DiMgQgpcaPgv7aK
j1OfiDeEqxVdEjgK9+WO9z1ZwH4sHikBvax1pM3z2yVxTRDdVAFyGgCcWfIe9gMiYSaHNyJ6s5Pe
D3ijyaFEISrN1ufEoFsG06FxvghrPZxgIdzVNgiufCA8MiMM8qnuzIonYtgS/xbBrOmvief26JmL
bwwXHwsoK5Pct8AJ+0EszuXsesMXKsf1BBEh3ye4xhIRJEte7OIUeHn+nWk4QckTLjV3/KAU99qt
crysyRau8W2+H3nIpMeUvwS5Cdw/KNA67BCI6yYsFekvlZQttpHZnzS1dRpHE93tEd5kiaWsvZ6t
xfUgUPW9HquH4HFdL1WS4Ebwb98Q1dtQJEQEJ0acKgb65vtavRz2XBpLXdAiNl9lDL+9rHianx+F
Y5bLGw6b3V5mEuR9rfio79pEdV5kCRB4erBAwJuf7NlIl0X56+SZzCqhwSeoW3hRh4d2LUPa1VZb
Hk1Q5t+FL3tB1yeWm6hrbkqHaVzq2vN6AgHZU/DjsUyUGM0NiNW5r9YDrAdma4lkhaFD+jUJU6zV
f9M9WslyYf8QOLMl21fY0ftfA6xYFHmcUPPnrs9jPOM0Vk7HYoPeo0STKC7MRBOtHp3bJuVYiUXF
P+LiuLRxw76pyq0pLemc2M6kQPkSu8jFDXIIjtwCRVlk18J1wJLb0420FJgPQKnljGV5wUmAAKuc
JKnPcri5hPXI405T8lNPsE/P6z2LbASeCvQsF5K1N9v+j5JnSqskcAI4w9IjVXDGhoMM9tP4KM9r
ZTJIrl2EoIPjhr16pCRyHka42o6fjctQhn5EPV7EOuljKUQcL2WF/dbDqkyk7vEHSMpw4MUm9qw5
7fhpGtrL+PKNThQVUHPfCEl7bCtfQrel+d+6NBGXBmqeU9/6wkrPqADBGbxhE0bFN9naOK7iI3g3
Cu5P0LutZsSDTNE6EMOPdBFdh8syRdfXuwyCOLp6+8EXw4GRXUl6iL0fgSSJIYLaKhpsys1cqJ0B
GUqTxSVoi7TpVmncPfeSg5OkhTEHBrZ/FqGg/6SLykW66S04g4UfsuQ7ZR269Zt1XUALYFqX/tm5
fr1bgROfJEInYZmXDZ+X24N2zt/gLUDNsFsJCN3lLrLU6suV0Ph4NloIGVxcPsqbQEyeV1wA38BE
rSvZQhd/6ArEmTZ/fiRqGuCS1H8C0R6eF5CYwsIUQu5ouLZKLMdDvpZ4WQLO6Bx/vF3iBGI4zo8w
cL341DB7LAzwrZAHtERhvLMsuUgi/6DJl8OsX4Om+/WtgXUMUVbWuiuzAowP8Zq3zmLYolPGniQn
/GrxIONO0qqvLLeuz3q8/3LL3LUGgbb59Pi8g0kbkit+rGWJtn68QA5ML6YxlNA3vZlHOYFr+G+b
FczsNkoVSz0UsEffJewVitRGhzamQnjzzzNhjzp90xIwnrxvO1Skn5SK49zsoFa0HQEwFff8Jxf9
P2ap38kaLbEbmC4n0CJRNI7+NA1DOnKB1TFf1itB9nRTCW+AgtNzBBvJiZ3filwCXKLMj+gQfPI/
nyArdTeoDPC78kdmtxeMR6Vuo/rDkUBqKLTzoHt86YbDRG+dU6JSq54wVjBVWChPM1MI/JbyVmRQ
pdfjaad2DEqNvPkpXcaBP0UCk++uQU2VIOftP/w93FUwRTHtJyc5FO7lcuXKT7MnPgHTk8rXn606
nDjdYB7eviFT1zd+/hg97lAFR8SKj7IRftdGqYKkLs93zGQ8KHw3vyOFUY5IDlireL4R7IPEwuXp
vbarZ7b/2UNFR59Aur3NeYFs+i2KO04OGwKz4yBSZHLs4nDcyFhkLNTruq5ul0v7b/MGjVRGsNC9
HDajO2BHQrWGoDb5yvLMFySb95/8dfTx4/lzoZlZOJJ7U1D+TxCV9hVmBK0LEFMBKzHZHLvN3+UI
J1PnYaCePy0SIuXU6G46fB3vTGNVlAdFcEjtb2kTef+1hqJZIdV4MK9Hd7DGHpeETXdV3G4+uLle
9xiKprGXlUjQKfulEvMaesSf6l3cdhOZSbeSTbYTJ9/YN+TOT+V7oz6voiGqp4N5s3f66U7ps4UG
DZxvNEDaHKY32NyQ2JBdIxlze2wZM/Q+Nxa00nk32iOGINOO72B8klas9w5oaRG8Wena/8NAWVJp
aKxIQxh9kW8CSWyhzHlXxGBJyS7cXk38VJrGOLGoOWA5J9PHDLzhGrZE/IOvEXHahIAvRfKNS7Sy
Ng9H7OTz+8R0mHIdMODwelpbUEtEZG8pBhbYkcmaizTUxD+bfFDCBZ2c3/BLXrug0p6F3sgV55UJ
cDSQHn5g8EbK2Mr2v/TSPb3WnafDNutptehQo3DFfj7jopdniSebV+3egmztMm/9KcMc5CzdVCvl
a2RSBLzOIM+/hHUkdHasInxs3tOiRNDS/6Qn5e/3F/Fn9uFOOFrJKHJtKQBmbAwJu388NPPH8gCG
NTNSrl4mRkCpBdRGPvMnAnsD93yUegldHPcTA4IFJo0w10i+VjWnxwX0fWDB7PH57jJVfdnHXRAF
q/eR29wuhsoRgCn7FIlh5izwHct3zqLLv0zie5nwn8xUxulpP2pbTJmqNeJGES6E3i7YE0C9V7I6
/9HMyqhsv5YRUXRPrCImJN6TJpcnlOxQDT3lkr2roeiL1B0v76p8H99ca1wpFeoKJVpi7vf0/7py
1uf2QMJt3vi8JFFr9lG2PKawiJf+IqxTdI6xQrIiVyyl8SWRN+DCdoFyN/AMlLXlkmU6oatvfCu0
puRfqmn5mELMRadxgV0WcrQdceH5namE3V/VpmlC/bIHaBnwcmHmifOy665JiiFhgeuspaSoMOcn
KAAyp1IbiACTrh5m0odVMp8k2Xj8wPHf290zuEas2g49PNP2pZQWzb3yFU6qGf2wN72Qwq7L3e6A
CPBqFipMnKWkZxCOIlZJWK7paJpiHgpqcuvZUpYjjOi4Ncz+OSclZRDCKAYf9EPyaSJZQAkfoLaF
bn2eTfLJPdU22qzz9ERCDeeSk7NWsgv4d4nLdq7HFMbkqZFl1pZAFVbNnrWEr/brN4HWV2Dinq5/
kD+5P4TFX70UkNaRSzjKe2Rfmx1YqedKc95E5nikxSWmia+VlAxHVEoJ4YKYoODprvNe/sj9R2qj
Lds2+c4RflTZ8WMy4b3maICll9sTWl/E3TpX/8S51EOB3a19dLTBTP7b14b4PqLsynsv0No2Gdus
oSJgygP26IXmljAoY9a9qRfCeNhPGqo7GQAS2PA0pewB4zAd5WqCHD0b5JXKk99hSppYC7r96/tK
7YqfSsYKleexB1nryQUSRDGa2eXBHlJcuW8DX5e2SNSJ10KJvI4x7KCvrrLJXEbr9SIb4LeiyQuk
drQGom1c7Z3wYI5rhphxMCVdMKnnkJ3nMJACiP/OlR4FajD9opQNW0yYUStu6mdB+VH6JU5+23Wp
gPQy0lJlw5SVvEWdf71HWeeIOkBaodY2YhQg6fgNFEVCuoPIwrelbAgPXou/jIik+PIGfop5fBMk
gHRuC2qkh3Km9ToU7iNx9rdMP24XK0wVCpnQ2jEk5uGOxaaABbBlbnLampELYTEyGluVFRf2NkeS
ab7pkYJ74+ALDKKY1BNIvTJszItJGFmoRsRR+az2ZGC4zlgKpLkZ95/QOLCYDPfi8NlTg9w+tTcs
QXq4gykRT+Upfa0VEmwrU+48Nshr3x1GE46VtXKVccyryK0bMqlBPDskOBTpKjBKAN0OE6UD8yw/
jKRgwgDIDxcfotgCGr+qv8D+PdAwVsKJpI7KYFREswVZJ3JekwLxd1FNqZL3Bj5Jhzybatq7biun
IgfVTOH7/mZPy88NpBjGQP1JLbMLGSk1Dv/zHrQz5U6GO6cdOzIeYCliHve8j3kP8fg9gUqkOe7i
zs9a95F4Yam+Tyn+JkHmHPGuX+wZa8X8oAwEM1djU/UFKEDjaMbTO3c1skrfcg/DjE+EGL4c4bXV
FEGKUs8/sxB2FOA+H5MCjlaGurODLycqymXzkMKNcI9XsQgwk26H3mOjeGvHoijpuqUknidcupZC
KoO5PI1h8X3QyTT+27XmnM6BkJ1u/T1nwR9LMVbEfoeJujjnnT1bnzABYQ6sFo66gElB1lGpNLh9
3lw5FJIN4EQainTgWHmJBgysvgXWtdJGSUpvd3mGH2+07n3p+r7dbM/Ajs9Prsvtop4gNTnipVBs
s7mO5G1cdlgAlb9iWn5EdMc7nrW+mVdOGVaNn6pP5n4ICaHn/IjJOdRzbyZcEMMR8KerPQ+ZWD8d
/1SI708jLRwSRg2ecuFKWDh9VChipXiuz0FHFfQPlEuPiJXMZCD5Cn7VAzqw/i3bRQfPFxg1DzQj
zH4sEjhuq/8cBbw90NSSXISa3ZTDva/Fd2MfmM/16fZ1Vbc1TXkEJIyJEuBmwui/8DLNeecOIRqK
h25ndwdNqJqeUeR9GG22szn3TUkO/JcRecFfUBBXQPHbti8h80oeWWZTJPI2A/CBr47g+ihTortG
eHYfL59e+gBvJ1DgX053kMmAJLelCG2GZ21YrAK6vjPa+cX8v8jsvXFeu4q57FX4sDjw41ZYe17f
oBqQS8RaQN2fxOQzL40tI8wkFBI7+98NhFUEEJ/D09UD7z9b+YK6W9QlJdto0Qh28niRixmNQhrT
XRMLCdFwRnpk/d9HdSwoIHagrEPBhvQNQYyQ/k0vMXOhuKfaa9MSDDQw0nx27ODuC4AppUY74Ybg
uzCx7LHNJ+YxUsYB6/ZYpAhYXX+gDOxHyeQIGobMuAg9KbUFdiY28Z7KZBczA1U18chFwRuVpj3f
KqgVayBZgkJNqd3Vj04Tcw6ijmnROu6Cc3d5yo+NEetGcxZYKfpmFTdwh5WgRmw0d171TVyDuAAJ
Gnc9Ti8LKNNMsVPfBCyyH0X/8AGnVke739xDv0GWYzawX8tE+7oDTVK6OYMDM38V/MSwXE+b9l/X
llz9fRYjZv5RO1wDtWDPlX9UVR0+3n0KPorSU7WejKcEJ2KQQ/oZ4RoiJjlEXWfCmMzW1cTds4L3
1fFgWxkewxUQDQvnfCaO7Lj0v447yx70WrZ8RhXsL4/gokHZYFUUuy1JV9MTOXwTy1mfT+qn9iDt
/B/9HFTPWibl9MdHrycw08cDFJjrslcyXUoGoNcG/dFt9Bv39ckUnLGRWPhCPbGThHi/y+H38Ku8
m2MfRylMhq4FfzBB3Gv279xk/cikwCjaPyj6EgHeKgtA3hWpPRyK2jCnOoXq5a1t72IEYSU1ocwr
N+DK5hJFHQdikBgzlyQAggA5NDoBjgXVKTKiXUCrefFWxIditUBjUOeEFo0CnZoCtFIc3wTY8GR1
q9xpAXXVM/2MEHcjqJx5rzXMZIZWzo+s68RX/3FhqvPl/lr327h+V1mUtepXwnTPgDYxnXn4Faje
oEZdl7eZl5aSrL7DYYG1G0IxYCsFQYZKmIdPA1RMIJvFW3seAPbohnuyCkGMADCtur4lO+8d8gF9
zxv6nMamUXXZixOfi0W6Xc/8Lbs7OyHCBklAgCUrt8GvDJCEQyMTRL+PYhDiefJsPapYFVfr1Ipf
tvGm3kqcEHdCC9loY713mtKxluiyydT7eExCktxAzkrWSLcbfXi6vqRYw+KBAYvbz7dilztxrhmV
ORzvvyZQrCGOCyHs1U1Rr6SnAh31KXW1eGrkF6a9Gv/u88V5ZQQcFZ5eOPMTG9Tcd1DC8d7u86C6
xMHxlcgoKPmWA4t/C5Sigj/UjFdrvZ6Xxwe4QGTIT4pdV3SG9EdHK4Ss5eFrj0tyl9B0yDvSx/0e
+4EzWC2SN/trFICJ0t40KV4/Z7vBxvTH0gu/RNaOgRpim8W01Hw/Ow+Um9XP46KEwQ+rhDQpeG+H
KW0VF19VZ8O2yUgfekb8nckzhQ1jTGdJdgGg1vl0izruvqkSyOem6B9FwimF8WxUnoQyzvrVKWnr
pj67mvzM4qYJ41/4ZiQs85yvW6DZxZc7v0gg/d1aBR20zRvNsZ9Yw8kTe6ers/jToXsoixGM2SqJ
Z2BhPHdKH32tS5hc9OjYAOtAXSBkjaB28opZ0RpK/hDGdf2uLHDztwALwc6SXMNAKbtZku0X9Jh8
3D2Mt6xNLLXdkTyw2w96xUVz8wbTRRINXtmQRAgML7aA5hBb2Z1a4r+OCqxeFD77PRpznTDRiAVc
WVmtHaX7q8wlY0llk4141zeQWWOI2+8nYGfltP5SFfyJu+qiwYv7gZIcuRkrhqHK4y0YvymePLd/
uIumaHkdLVlkxJJugAlJRXjn4PRLLFDWAxqclVbosfHWXg9Mm3rdUje+GXHq6Yphq5oJ6iGJwgEb
4pPBEQ567diI2/1mhuMtiZOBVdV5r1WBus2U5XmFkwfvI2jRdsctXxmLtOHtysXWH7sAji4Evo0J
OpJ0Frof+aE63QtctPx8p245GwK895OX8S5mGM8G0I5HwOZ43O/N1QeNTQWRaq2ZW7O+XoNvsz38
F7mDdo4v7jXDV8aeWT0nWLYMPbH94s23+4RNti+lIj1Ho4b4KlBh+671fABzzb+B9AKeJuhLzvPi
UHa40lZIa6Z+FZ5DhNPKMOd0jFj0GIEnJM/opcPVG03QhS9Nqek/XyJJhPJZuNafrP7zil++m82y
3AoQIaXLXMhZSx/aZVm729kQ+DItQj/qCUSJZCYLGkU21r3T+xTVa/4dHuKIRU+PZqvsI65YM5Xv
6ZNhBck18EX3EwGzaK8s5LuPzcKb+pp+H8pBZyCre4EpEwcW2xMnFkbUKlmVayHb+QhbmpKx7YNh
Nr5IenB86vzbctvxKHA5p+HDZiifWJgmiPWcIl76gMWGtM8yor0C4PTR4/M7d1gpwhuneolfM3uc
v0cTaTB693Iyie93YCIBYQpcWWzeqvfBrDAAh0d3Ni1gv7uV2u0Jrq9Vnt+HXa9t5jyuIoTN6IUT
y08DKzpiVRuw2p+HmGXZz9gHPc7P/AxDaITRxbD8UdDS4ONYRbOJMlMK798KRZzYblsI/YE/MAmW
t/XQIATxvR3ztDNlX4netUQMaxxfj8yAoURS13UKqdLrG17abRWCnxiuna/xVM8zbTwt4EpSHgUu
sZ9DFAHVl1Iv+/40A0Mu7awwWM4TnJg61f/qVm3eRQH+2zxSz2TEepCYxsCwKs7AA7KfP90bZ3K/
Eit5xQrn8PQb0+r9/NPcVeV3mBNrl2iLWrWaaCUIg3/pFyY3RzxlMm6UCAmoOUeX0mfaYt5oDe/R
JMRuSEVvv5En3UzKZAQr1kH00OuND2KLIhSQOa6+mPyrIkITVkTT0vKec3K7I0vI3K98bPBhveGi
4iYGqealKwrWLgg6Ty7DZlUtrnUdKiY18ZSTt8A3EkZokkAcgSUBup3qj4m6JCb8XHtc3mFhC2ys
oQjD604QZhtxlEb67scXr7b+082U0V2/jcsdTiu7N+RF17Fq8aOfZcG5/fAmRdaAtxfGUSExK3Hl
6LYM1/yLLvjl6EPuWJEROfTvcW2IcSiT8hvR6cZlt254WVvOXYbINzJcJMq77RRZBgjCvwe9Rqqo
00KK6mUmjar/4RT5fWMGspBbwq60+E0Eb2vNNMLADgEyHl+/s+6pvj3g5a5w/NRoLs1OpyeD3Sl/
PAHKmGC+wa3kgMO6waT6xHf5guc6OTmKdHDx2ZzlRJ6Pg4k5EM/pN1yQ97jq3dAEffpKoBB27RIY
ZhBCY7EQU5aYJqqrWhkb5LwBfa3rVcz2c7Nbp49EuqHg4hstnGFJffXjuotGHsUSFT4D81QIkBLq
wrcq5fW1q0w6E++K58SpZ82nh3sCeqvTe3FvE9q92KKkPucuHanXWuxuKA4r9ryNUPfGI2SFWimW
wFgKVD0Io+uTRWklPlb+Z+q1mdMPCh+hWdwUdL/qHERw7fzM682Xuq9cOem7i5FcxQF+qgNNK6tU
Qm6W22nHvDgZ0Ig3kVpJXwOH7Yx/sYJ7ikRpqeIp+gywzkoJ8VydEUIF6x92wr5R9QiQQNAj1hg3
njJjtDOdmBQnP+Xpuueifky40Pr2fsMJrB+M0qL2TGA1QfHsqo7Fw2Lp4cbFbtJTPAya4kFfOo0c
rbpySGfVMtahXyyAZHyAb42oQFgIFBlTuAF+o054vk6UoiIsDyM3gXmm8iu7hdDN6TpiDar94o/z
rP72Fk5ygMMpi9lFHK/F9b9wfcdaPQyAxGptC26+IlMWq+OX+/HgpToBcI3hh7nbuW6VQCK+nfiZ
zNmILRIoA1tgfB3X7kUxQvW6BiCdWHPSfXfh346kepVO7d+fCHXGDF0CB5cy2KWY2DHQG2iLb7FH
J1j0uxHWSFhcZpln2VC5e/VRDYJBOgX92DfWNrLapvTAd1TLoOYTmywqOG87Dgz/g8HZzD9+4dpi
ejkerLvM4qYS5FpVxk9DiNZFcfEAonDuwP/JryPDWrsLpyAmp/ZN3wsU7elF9OyItd99FZ1GzNSe
oNX2GDOhSeQxoSfVenBiJR2b2CEVZ99o1SVsGqSmljxj9B7fLX7Bd5sh2h4gI5QpEZ8szDQNKhhP
umJekrxisRVnrimg+xHzaLMBtyw/Rej/PsC23odg7J0PkL/Ov8W2smI17NdLjGdrTOmY/zYLnK+0
u1P+JY0fXBIzH4OVEfVk5gUagkMTV6xSrFmRt35gN+No347Crg0gR+pP0YL9T5sN1kIl0zZJoYtz
QBtAq6aez5I8KY6FSMqjKMvQT6eWHuENzLDQwomzZ2O2eEZVgtwa7Sv7B2xd8w/y1vq8sFyGbdMj
PHX93nXP0FJJhPQv++fAH0bxOQD4sIu1d+I/5Djl+Z0IJGFOf6cW+S3uQGOapldPM5oWQL2SRFk9
9Dqafv50Zjwp03wqeC47P4XyQ5yKdsDADACh8mM8uNwLDF2D3Uv6+WYcM0BDsEKQC9TFaCZdj6oQ
0es8pHomggw1kqZCizZ/W1AOCKYtI1Wa23xJ78QgziqIjS/Qy4/TJcE7jdld9AzrEeuhKDuFAHpO
SbKDr/k3s6phQX/JfdSd0oDbdD1QnavnB0n1F4hUixVo79oeD4TbRhcEFXLEjmJMzVJVkUjcs1Bl
3L1CJEPp49gLKvP7vYAFA1skILCMsAQGTS9Xp7lOuwMbaVtCKbWrFLRGrxZjo3h7tHv4OZS+xLxf
c4nfOcTDk1cAuJbAjziUawpKPbocCFT2UpSHOneH4DkiODr/Qh9cPLDXZT5kWOPyVEFOCckLbUv3
3kChQcfD8Pbz60G8IPTAsomyz9ufx3F57s5RxxprpLWyiDiNb+sloHd5VASEhGAh2LSYIzFg3zqI
3zePRuMKVSVPYKsqJTHOzkToF3zz9hVok6MtAVP0c2q9dmSsD8UzEWEma2OTqtTmlVa2ZlicIveX
0w/Cibt0SIX+o3Wl1KyKx6MMe1QM0ZKeYMHtWKjyocgXM0PW/xBknZqMYiFNFsylVJ5fGWMCEZzn
F+6DOT6W0OD2rliAZwHv0Mk5Tn2XdGZYgdP1ADZLSL+/syg8ViT1oYcS8BM1PQ1P4zQNcIsu86WD
9nLGod6EcSsKVCs4wJvs9/ZKvh5xGcXTkVz8axKHJY/m2loEsVQW6Ps+F+qchV1ARRKdm4iuPRK6
x8IlbP/7ar46mi7AvKa/2dkyhLSJjYu1apBaQmfc7coYy7z06KxGvJJVTqYqos8esPIyyu2x3GA+
DWWMhyyOH1HTBjnZj1BDvwr0eRXJ2ujbvuxY62ucD4VhWCjui7ZZ2WsirzhDLTVwMOM9mY5a8iRh
0EenmKX3/QMhGeWNj5EG8D7i021/0BpBC1lqVLcffwoIyWm9sKEb6Eq29U3l8iP1vN+am3/8qHXN
AQjwIzVas2DkRQ/c+yd/+x0YnCV+8SLVIBUjGfTfOWLdc4z0c7XNLTXrOXr30O0JSSRXENWVMcn/
pX9711qtl+TMikWkuE75x3vcbs8VSpOV9/oG0Ix/eib3vScRRPoVSLn8TvyMJVhfL9i5JjtCA2i0
bYksw/vHGF339CNdKzuE/zP/gP1uS6/sYIaCl1O2wZmSEwllqyKs7whvfZWygTNFvUFAXriV7ajl
42DuhuuqLx2WpRFC2E4o3BQ7WifMAWZqLMgdrHSdnmQ8kXfw5fyvDEmxec+JSA1HcWFQVp0T2bPY
yofWdjKh2jvYU8FMs4s/qes6xtLHH3oEoshX+wccfEWvneqqhDlgr9/6kER4b5abMrqxOixQIRhx
qvmkhyiUhrs8K8Q4g1/CpXkWdA9KIRDmyQRQfdjEjSykrGiHwZsEueFDYdzM+mBA3jvQIWpyZOgq
OuJqQjzEuA+ytHP8jgGQp+yJh8PlvAVltEgPqp6B1HvuyYvNk4qFTYDzNZyMbd9JdX0SWiyKdY4q
K7nqOqfyh8CfS6D3SDd/C3P1yeICOyTU0dHR4BHvr6WVZXcCA1lTdooXTizNVULd6To6N/Bi0Cbu
qxHhwlCJ+XB5FhBn5LBUFnO+2RbJppeP/FHTcxh9KZCk7yvOHSLkHTH9NlBCFt6U6lOXntufYpgP
UU5W7V9BbfZjPfDRIGpe/5QcYVxfoh4xZy+dwHwpS8f9C4sqpkrpQUS/FxYTara3bYjcd2T9eXaR
qd97lDw378ZxxuSxPwmsh+r+eN80kgrnXIIUChze+3xneZz6d1yWqFwRvF0nZqZsrvLrgcHvoViV
YEUJio+AAoPENiLA54s5r81FNBdG1MxiNWeIHc/1qPV/r7beejG7oDDW931ft22Y2LuZMsliCLkC
JTwsGBiG/Q8jqPS3l8FYU4qr+xN15Inag+Tu306F+wT2ANt1MRAObPt+kV5lFHxg7OoMFyLIY1GV
H31O7JBvm74PEqH8qQ0/DEn+kb4wCPhR8YNIVkxdFFiRMolq6I1vkQTL7+hxMauhKRnQ0+0xWY5m
Hj7fh7bA3NdSTs0jVx9Nau3DpgkYj5jirWNhXoa1J+Hs9Df5O3PRcJVoqmfV3HObYzdlGWAgfGSd
vNnIa37uaStjkwHc+TjylbKJ+zbpura+XqrHrkL3Y9JOSl+JoPNrDrv/Dr7TRGnV4zbqRS9bVpen
rdwKnebJEHXxAcL6G3kM273vDN4YgCm3lmQQd9yFPWAeg9dVAG8avS9X7vBliVtf15jWOwXpMqkI
BADxIoO29KzfAMaIvOoPyJwOD7OqCcB/u+gLZyalu7NZw4hDzvuls/GQHNHl3qPKUZBmfZTjR1ph
UnexoeeDjalPrBhfhtSj1Refl4h5qUa2gghmLXnaneDyT4nI5xP50rIJqEwLAq892AYBrys1EeqK
nVITPAV4rOLhWkmOFNrHCJ076hoTcvr1fGcli/DDNEBZnwMObFo+B8pW9hwVT22nwYcyfz7WVhNL
hW78iUl3o5+Ok1zh2+z3CSU/sjE7Z765RL6mR2P/hUEOhlSULhe3fpwC2iHuwd/4VN9o6qxENbqq
SJbzYzEq0t0AHcTVYtwG8KS7oMpNU7ScYIyGh4X18OrJtOd7qkAa8gVlputQhKziuU35EfV5BU3g
P207EA2Z1EUtt0BaVdl0Sku0xft3lEMnQZqnyAWgMNIebR1JoOIJo4/rdokgZdPDiaCHvfmWatdz
JCR0AB4WLdydJPLt+xUc3rDYQCibA3uRNJqP0e/zoWyaPytgM4MCds3iAvU3OD5yGQmNzk+QzhH9
xMxJlhEmuywE6Ku0asUhGwDrrH9linI3KejvSZOCK1kWXN/jI3aPRYZ1Lx9qPvcQfH0pshy7cIHP
wnCYTD7Wh1H8sLj+Ncg438Gh89EU287+gqQh0fdmnGAvkX2uZPtH/3pziFCxoCUMdx5olgA6c6S7
Vyo6uTuSwHmRjmcK0seNO6TQXfdP38dkY78RiQxazjliEtwU0qSU2rrdrf5wKLOAnKRkbAZWXZpN
6C7YRGrj1H2MS23bj9jZaRkvNw+zOVJWCtkbpNT/2b9nSNow5kOMiU1kaGtljnRlxFOgjhHhlKXa
R5KfG2S1WptBMedPaMQ5ChcY63O1zqI7xAr3xRS7cdcpbWAXj8bPyhV+W/Pv1j4GBG4ZhgTuqZs1
GDYDEGfny9M2ZpXNn9//eqInxPvg14KE+M2bOWr/6RvrRwrG6ljWDVa25rqcBNCNYbQ2sAUNChVt
RPm/RvNPRpUbXCbnbDjR2ZyZdWXiadpSHZ5/29Rraomfv/74luJwa4aa/RBj3IpESBIVEUElArKZ
v8K5LJgzxhuofbjyc2RJoXlZzxVdWzUjH6vUDBpODeAcScNuLvOEjDXeDSiurORK2/1rGTU+STI8
ClzybCJq71ELXHUA2gEpk9nZcSnXuu/EZ2XsayBfadj1Yw5Sl4wImqY6VDoCUziBSOekUp0/glPY
NLuzy33NNhO/9FGCofDKgpgBJ0WMUj0TVOK0LVhG9Z/WiaxpbFG2Gt1myp/ntXwnelW7V5tPgUAw
NRcIPel9KJP3XfuPHSBcwbvaZ09SWMuTnL0mEcDcpel9mZH7StvYPuHG6Qy2qQq/vZDnKRZkzcYC
yM6vIv+6p7fEDJ1bneiK3PN/7oxXWkX87uU4bv0pRGs+DaircTRiK5x1avTQrOq7S3GmXSJJM38v
9udVv4I/hXa6Gj5/KaZ3nkTS7DxWBePWmKzwXNOWooLX3SiKZV+RklZQaQkYl/YyeMzz/GzMJfV0
1xqZ8shMTKVRvpIzucvu85GjYHUzRl5Y8ar1qvkwdXiguaAIJdY3vV09088uxurq56gyj12vE5Bo
rITU+qNMRym9ZKs7QskvhhyZOfFaXnh5RW1OTiuLdqI0S9KCPltupaIDCxcoDklsYupMEKuCYRz6
MBFBzAhiYhkfIWfEujAtvxxfIqXL9z5Z6zT3IcZ9oSftskJZntfcx5b6aeE7RwHMsShzGGcMnyY9
adGnbKNXxxKBJMDBb2BL+ZTizIQluYUhQHBMjpuCdnSBITGQDQwns0LlprbflZc6btvvKADMm7iP
nayqTrXAO8uQxVeTIK4eotpN7BbZyAuzwvmfemgzh+TSpfqGgm337XzA2aMYRE15Icv4VilaNEz1
KMsDW4Wor9xwEQWOi2CAxLMHkvJWmnYenJoqiFRQYwejT4jDMnZDY4Htr7PFjFJ2sVtg9CHFFUxC
uMdizfeT9liRZBY/RJ+I5CiAVtBJS7qbehXOqltKEfjFWUnSveyiNkoxe22DAiHAAHdWlmyVSLBp
pqW3mNwO7vi1cW6tRJGd+wtAiTbr4ZS5pnsG2Jso5oXCZSjQzNxhcE1jN9PPPp/5HoeUoPlZ0G0C
Xj5NjDJW7WcCeCDmydWmkCCbi/7DiHqnH/SUb4x77VYT5MjNqQjvm4S+b8MI1Hi6xVhXgQlLc95x
BZfUN4Bf82ZUeUsfeDTbhB8bnImV48P0f5MBf+d0CGtHxr8zPwkD4re2zvh4RCKjKkwKDB/vIAoD
8EKBZ8Rm2CEGpFbChnwfMd1BCRohP0C85kyNKYYYjKWWTtL25x0OjrAXNNsbpsLZ2OS2EgPK8R23
cf75xKe1ZHSS6qEyi2iwqNR81dgCVb7mVnMvz0q/NSww7kkBB0gRImfCv/ZKnLJNCA83/+Fb1s9R
vuPjGTXLd9u9oDMEVVOAHOlfyCL2g5zzSR7V1FSQy6oytxfrOYDnipZoHyWDz9+Er4yWdo2tPYp/
2szZYw1CMkXtz+uJv0pkSs4MVctcw4IY0KJdvMRYCezVWs0K9dWTyox+V3Vy3p1KuASq2smKmCLa
BbjzlYgJpz8MoC9Dqh8JzH1wmUqRI5IriIDHf84Vr1O0u2bbNwdj3xQKPnwR5dSvqsOgjgtPnLQR
3AVA6pEe6tJ2ZhUVznlJT24ytbCRyXifmNzVp1KWgM4yQay8oXcPxgkjccxcLA8Y2NZ+w7GnZ4sF
A++RIe+ORzkoNpxhj9ZvM14kwPG2TFJpmSyqm7gIo7ZV8znuWQa6B92o5oDbNCF/aQGRjoSIwbVS
yRg+l7Hyd3LulU6K3E8EidpOYN4LjXW1uXz6j/zEsmNUZ0tOyM4EldX1JKA3eFpU1rwn+sJ0dhbr
NntR2F8E4siPQBhrOG0kjivUigzHzZCKrTaqD1Ab1qQ3APau0N7Jfw0SH9qnMdS94sKhtDPXot+n
a1zwuQAqCXsCZS8uJkTag0mCP6c59kCZURDz+NcnL/89ReOA2E/L3Id0PiEb7q+sYCM7ynuIHDyF
JZKauxyWd0S/KzMc8zzpL+Lr6rc7EchqfQ2s3ELfy0EtuuoKb9+/sZydHvemhac59vnyho8c100k
S/QMUaJeKeSN8EDURDYgn06yxXv10g5Kub3ILKW7Brb/LrVjlySu82mq8yic3dquKGQStwdrf9BL
z4nY0snw/huzif6VieW6QyFdKq/3JNxyGX38P+CE00esJ9L9kNtS/FIoFWtJOoxXr+Ih83AlT8sm
+OfG7XtKNZNfCXyHvg848R7c9yxvGYbSFBiEEjcqZU0ktUCOQ2U78IWhJyQAhVFe+P/QeJNkj+DY
0ZMDzzmAsFvjoI5R80LAAxwQ4fw7RHfKEjeDTJvQVGgqkzATF165byLGiSkTc29DwZOPEB41nwwB
ymlSuLbgsiobhleh7X18Fu7ji786OcVEw9A9LhjEwP5hwJsmnRNuhPZY/5CyrsdSzUz8E/YF+C3f
eFjWP7WkNyFTy+5yE7iLAfU6kfW1g3tM9syymHxoo7fbKsR+Pc35nVaD40mieUe3SfMsbleAiahX
S8o7bZQMgg/tPkRFGHtU3AtBLs5OrttrV+6U/STu/YlnnPGMfS1zfDWcWgQMDNPHTIPnp0A2kO9o
VTRhjNT1mHNVu2rUhldW9aauYnl1kxwhL6JmqCSKilPyuF66D7r8XnpmLbChZ6RJCVpiISkyUO0h
tadfLmyiZwk9/6wiqIDRXB5PEWO++KE6ZYkXeSfDvdPXppwdvDH2UgeWJDheO3Gb7cMJAZSN7Aa3
hpARA1ciVzaC+B/r4nUZM1gYBRtIxoiQ+NqFg/U9FrXSCDdzlpWzP5FHRJCByGLBRSnj7JqLiHUc
Kr/KgZ+gzCYlXPlCKRxm9VdZDizCNadabX54QzhJ8eFbK6pmbEdKZ/g2vxJAxrJTWRIdIIvUd0t5
l5RIsAWL/qKjvoI806xbA1KWp3xFN2a+hTaBnMWVlNUAgOLqvlNHaWlBFVG+g9iAq/SH8G/ZQpI2
tG5H4sYzUlfQyP+EYaUbPtqDF6FcgG9tgJGUa1J7br3PHHrfwpt2fGLRYTcUfnRDSwOr1v3m8Mbq
KhirUbbnoNDGLeU8ROkNBCi6uT2zI7aw1dnhwck7SjQb/rLSVnAMpsXoSW36BmAzw10+nl8CPN0e
YqY9xn+886NuLPqoKUa3Db9eXrw7bIL6J1AFQBOfmWpGim4UeWhdddEuxVWZ1Fyv6B+AjzRNterp
Wd+AJLYNtTR4cpY0XJKrwCWcEORpDTeVF5cnwMgRxIR27ljDh+Pgg14UrnExIyQWmOOQhRjHir2q
1rcB59HnxjaK64jlwOBZ3WNLD38JuRvre5ee2ds2rQDLv5IrG0zlGFsMJ3p/6i6pivLjTpf87sFa
YGlSP8pLNVph2+JO6Y8E02tIMeewAdTiOEmISXGgwYOFQ4KfGwxGFT4S7UzvDZFHZ/8/jMq6vK7z
ht/DQuuMTeZJZQp382zAqwwyA0FFAVFzr1kbIE2kfMGi9PlalkwJPxRlvhGM8OnyD/1w8bbI/lw2
qCSkrkCeB1QJcYO3lhDHb/gbvvvGYfdxIb87p6LahhjPOcN314B78Sw1e0ggBIZAsQhg6G/T6G7y
LEHh1cE2L3JfyDsFZ1mwNUQqq/vkHUwaOINPpuvOimdlyBvHJVM06ZGi4ShNc8yk5nJQu84M6meM
zZSwue1mfRYJCllGv1wabxjsq0XrULuY8tUoVeoBUHxa0Vp5Y0QEAU62jyNaCZERevClTRXfO2en
kMpfnsCZAGHy6KHlbBr3PPmXSmBSbLO5Cv7jsaj81h5vxCl/IzVT6WkvrL9wGKxudMLyV1nRrjLy
B7LIITs1bDKfKZvpNDbUgPzUFhTq62E20hXds+iCA+BDIsoOni09d7HOMrjteUPD3cjwDlUuRa0e
DZ+gB6mHXDEiAP/lBSkEcrqoYEqmcOCeK8bgNXx78kKCfllWTiaC6WAJproEL6x1f2f/cb4FwLtv
0Ueid5w7/qvh/e1ku87mhdvNP8X6P96oqX3+p6PU2ZVM7cH2P5obHZjy6UbAIQuZgwev6Y0lg2TO
xWtwzLhlwxB9fEC8n68XFsocfGTB0SUa4ssj6YLgSpfA65tteeAZp27kQkFIvHq1M0v+C1S1DGLk
NcdJp3eqqc4N9QyGX6piJHcc+386mpb/4gUq6Qsf5N1NA1m7o2xO27ds2I1cigr9dsS5ZrSZT8Kh
uxW7iuhApmv08H6FqFpl2irC4Tz3ZjARAzSVzj3S3LOQZNgY6e3Mnnx1tYxtiXiH/jI7aRM5agtJ
0bGQhdF/Gta4hB71nzo/yWsZvtY6sHXupNOMJJBk6VPR3AOaegnP24JqpD7w+AORo+3+WR0vLjWa
CvrjtDg2Bd2rjCaRj3/0wKuWXW4GYqBos8JpuRztMWOOGaC33sBq56YebyKlrhSwFTlYIUxBXtbi
Mj6Dn2cAyktp61qmFfT0Nk5NRjOcGVLD5x0XJufBj4DJEio5qcnthMPhlTtNW/pgH0qDAkZvUw93
1Y5LTIH3a8OsjVSpswqIv6guBc9qw5KvNBIQEPQsjFL6bkzSu4jxuZZYaQwwix6hMjICmTxhZOfY
/8agzzHF6go39BuhSPmJyUlYeoL1vlYaCyEK7goB+Qt+m4pPBkLlcjGVwHDUl3F2EfsUPKy+iKp8
zCVG3Y89pDKKJkwy9i8pQnrqZgu1tTt9E+BMRsCPzLzBpZUu81TRPA2ZTSYBc0UI9qW6vV073Zhx
uQz9xyvYSYyVoeEgZpX4/bazkBXn1q82trG24++qR5550qPFfszYpQv0dExwG4h6QPqrBRLk5X6F
nrjy6ylMt52owHzwaPbL3fwqz9dGut3vp4w6ZB+v+cLopTD3LBcJbfZtzG/ctxolP5u8XJCEgGQB
3dwljXaimJxuMdyUXYX31z5bgD6cuitVZYfPqkEAImXrlzylkWAGpYY92mFwvCL7Sy/9x9u4orrR
EUVtNkSNtq2B8cGzbADlvNQFGcyw0cKCCmf3oYUuWQcKbas6LJVd8WMccQexaTDnxcm/WsQMXJam
XnFQD7mhrKdMFr9OxlGViQeqJdSjl8PZDgrYBUa5a5294pj9D+xE1vjbHByC2i1INm89OhqJGBPa
3r9P/h4Lo1g7j3acUxrL2oRyB8JbMRt3upFibTFjQMgX14DPS5gdGRXHPwkc1RJxYI2IcSePavIK
EezewMNuGRbpHaqvkergzVUxc2vYXetaHkOq2+E+ylyoDtAeG+kYen9Kn80kloEmpVfBnNjDR5mv
HdWi1VNsmNjM5kUWIeQW+tLoVunFnntLmQDSixlCSBFrI/x1bugjtLxqpU6wdQXIZkeo/7QFc/RY
M/FQK/Dkc3ceu+NXhfto3+G9D9qGJC/IgrF2/aAelExd0RuH3bTHJsvuv+IIn+R58pYEhM9Mk3RX
D7cbBkLgzdAKH8HEtvWRempDe5fQCjLTv0T8tfPiPGAfttoTd1oWp/8eDx1clq0mRr09b8RAxWEK
6d7DZvrUc8+TeEaIHIKU357UiRdlo5wU2/W0+HS+u2/oPriUWSGJjEQRrhSWNDmQei48PPq0zrEu
FOkNpmu+pMCsa/GP3H9oWU0KPIRhgqEXOMacpeKAuht2J0P1OOFX3Mq/cgDl7kcOeClLWjVe5wJ4
Lv2GY+g65D80dNNce45kXZ3MiBkpEypirUq2O1I4h50S/W9YXraTz6hlT1sFZeACxOrP9GK6EFiV
7F7NAMhlHzrC/+S/9YLjqtnjRjowGBuzM3h9La826jFzYH1v75Ouy5by9mdwUGLxiPP71mj8dI7w
natI61x1sQfQD5KzsRAWuUZMck+dC05n9H8ehykV0sfPxFjC/jRZRBz4S4jQzhyp1OLcACebxM4Y
8iasfC426HC5Q5K+F8rFBAb8KskpTQYX33lNwKJWQAlCAY4QNZrUQ4hi2o0/JuDkarzfSgXEqox4
qDRBKwDpskoDzlB0wLmivby/gzNvwiVfygiSU+cMqTTjI5F1V01a5awBCQZr/Mm+D93papyXestm
ijJYc4rH4Z4SCg287il62/ppgU3WZbi2n6h/8tecFwqd3HlbBWqET4L7qHP+b1kAawbBF0/r2TT1
4ESJXUcHkiOuPSRQrLIJxApIX6cQi5qQzNwd7svTuXMqzxB6rI9PYDHlOMyJ0HpLZkM7L5PTh+pK
x8OQU64tgbhaCB3GVGxKa7f9jyUZVB4g4sFrG0ls4690ZmxxZZmupBVdyQe+9dlVeoLkEAT7LTx0
2Hb3QtSQ2YCjd7h6P47PGR2bMGpOPsACCFARlSvt/Ih3EtsUVVWC1+4sTDhZYyo0+DU1jFQryyd2
ZOFZLfoOMPP3N80MwWJdfv9qNHMVaEpDiqVRGmTjXdeY6O0yU+ZYcr5KA34t/17WQVZFKqYxoxF/
TLgwYNHhG/iVAASnzltCkZi7/qOCJ2gm7qutofhlkfC6yxAyVKaRgXF+UkTH86PlpW4LCxc9syvO
na8XOd99+z5ghPuE4KxTc6OqQZwJWLRhUvTNx0pz6CQmRJbfS6d7a0qMdLq9OkALdo6XgLAom9WY
IzzofkESZeQtl+4dVjI8DTrh6GCd1w/9bArGSVtHhZ67TcpRj3kM4cOZsO3KctHUCE3B83F2x8uU
046CEVL5EA6J3hjs97ZqleVJOKvAqQ0KVOZz2wfUsrhTA/ssUWvW6SdNpJMeQuVEbExkA5iux2HN
TQJ+6OETSqFHmYHM+04WxTOVI+AT0X5YCGTO2bpODMWiimeScL/m+TvocdQoJyPnn8nva2D7S8sF
6aHkIbjVjGDYYglBhcUuvDOs4jvadrJbCBgZarHtlba1SbtafyFNIAOLeFxTOtPo3PiJUPMuVdPR
0vhT8bY2dBDd5LtBTn8Y/Q3ddaXVECVGlf0zOynoh2jrms3VzwUZ72tMNpMVUAM1fACIN8s5/c2v
p4DSmfNWzncd1YWHU3EwbU3kb7ntwPIMizPdwjVLZ4Fxq6DK064a+CuiC3DZQJYB4EhDnu+jGeWW
l+v5UcKcHK994uIV3m8pIhJI+R8a55Yx8nhwxOgzlsCo8CF3mG58aCUDsn2iQT13mO5Kg4mfgmpN
SAaBh1DbsQ/P4rd648S5y1XuKUxBXMW23ppIYRMampDY3fMwzwZBDaWUYMWues/pJ2+xyMG/9CKH
OzldWttB8tPORtHruJfM4eTZnrh+zHXChnLiKpXtbiZIboGSuWfVo0GzLQe+5n2/xv0hmpejGqb+
m8mNuKETRrWhKivX5QLT+Syvyvrists/xRKgvn7WqjxMSNjXAFdK/OeA+0PLcX9u5DrscBstY0jU
utG0QBOowzb8/FiouJ5Y86mjN1HqowQspOZHSyBTeKDBalHcxlFql8LNFFesye2H8A3zrH3ZhEW/
dRnk+EnmPgifZ0adP1y9YdcpkrG2Sjrr2MKVQbpjxSXiaIhtTb92TMhK4bJ80WsgFBIY7TnGD0MG
+EHzOm+9DD4mgBJqvVbbCPVN4Ewk1gVbtX6IL2qzWF4lsNHXhvAKLOXeTH8DmtyxePeyP5mKDPy0
lmZxV3uAeB/frwjq4g3VSURFHNfvr2OO4XqoFIqxthe+bfTXdSnVyqiiJ1eWYuwCS8c08p0hRtjB
tuKW6mqLlEID9chMKXS3J9PLrm2MvytCboM+QuTmNi8ZiTqH2NbpvXNokLlqQgQt/fFDL6E8lfLw
qv47dIxEdoBDMc7I55r9OuF11h8GjZBJBs8WPgajrQ76aG4w3o6mBVks+08AWNT8GEggdTH2rdoP
HGvnT8sfLNzuQHNOlho6ixzkidJGyx5oNCdkE0GsD8HKvaRGo2T6rdL9hOl40hoeq5+xaWUNFqoD
Xig6XwXOTgOLGuyxxg66aq+qhrsGzkyg5vEFQVTvHwC896IXl5FuG6/uLJeYOtwvOCYJ73nexSk2
fYwhL2ev40FGGsWBe1zJ2jW0KIFfpgkextCTSeYNNcShpcS54aY/XUk0q2of2p9MZ0NIzTK5LsF+
8aU/gnL0bIlzYtuEZXSxa5d4Ovtm8EnqooHfPpFw87fhNwxIZ1tP3n5xtnfafSNwgTc8Y9KS+ZMi
dmvIarW4DU2J74bAL08w/omvdvehcBjfXY+hVsv6Ouc7se0wqZ/wzoT4C374obaAdQns9yveZAbf
RyoyMHwK8Ccbfjz3+50g6vtpodoKBGvbN6dpHtG4+YocVFhucMbG6qFTRHOepwPoszXZaFI6bA4C
IKCwmmuCzti5tYLZC3CN2c4f/jvU7QsWHsg76a7ko+yHBHQamrrPThMUS6pvSrEpobgiSIRismkA
kpywC8FTEPBL6E//bSzN2cct/zI++sj/UNkFH0IB/P+TpEnGUcPod91SwCqatSNqkm88gJ5bt8mM
CYIJGsH2usacpBKZkzN8dtIufzDLX+Mq/TfzCImvhFwrSqMExj4TvZL2na71kcWoXWqGkV9RL3LJ
JMbHrIJgTbheOTX5DRO3ldieU0nN6Hlc79//ZLVDOcImJ4+sG7mjMgX0Z1qCsALFvgn/NukilNc2
oOfQ/ByUXRjr3gtCpg+iZxLU57uCUxdjus2hTC4I2SbiqRJpW/rP5SNZYgZ4OsR8WEcN/JEv4y9R
quzbUSPpRY9yMWfsWn1cOT6O2e7wBjrjDpTfgUEzfg48F4Lw75uz9GF/hPbmZNuLnMG5lZ/rh0/z
t8SN1P5FjZ6MS+R8JNL/MhicFgevxHcTxmmdTOtLsKXt4WEMW0k4abKNl8oFbc6+pG/TwYd5aQOI
XOCYlNyYswNVvEkku3R+CyybogRRGXGxQXehJxQhZBSzK8Lp77ULvOiQ3//NwesPeX/WkXMtBPAD
PNKgaxaLbaO3lQ8opbswkrtoqri3hfxnSj0MnGVqOV6VrpO95lkRb+BOEiUEjvlKO2rBhQWE69Jt
TWUc5nMy3b5E+uvigzJ6XWS8b34hC7iMBHvbNgltwwrsvVXMXT7j01wph2vEyWkiIabljF0Ers/R
mh87a+iCemcp3vvEi07k9r9MjcvzCwfPCyeNSnuh5j3YW3WqpHwmfXRfoOUQeTr/LtdACpw0PM1T
wuL3wtPDAe3NGpD5Ti8BiYldGFewYJ3JwK9ddah1AOguddGXlhqCkDlGzDcJruWvpRQtbj2mJoNz
vFJOL33GRRYnAiEB6p7JSodyXUhQCAhhRi7VB1Wid2Rb4dduE4lD24RhQ5VpGqoQmQniIUt532jh
EUJd8av9cgfmP1dbkleAhidzqCBW5MwcfAwS6E1Pz00KUJEWbNDm13TIPGafcRdBtc8NNxPvFl7j
biZGXhDi1VRLwEOjfuv9B0T4Di1BmTBNudy4z+ZncU8yPJCSFdYN1GtZQ+ZoeLu5s3sck/a6hy+e
jwNJ9F5ZftOHugfXz4JHB1lDMoegTa4CutOrsUeLoIitP4PAFQIyaEotRKzUivHtNX02ZISA7CMP
QZpxt1v66QDtBgqIar6eG6vb1kC6AnK0iS1Cd5XrlQ81bopH3dV8zItMUC6HkfMQdjXnq4DV4XM7
23+PmnfM2RRhdbkAWhnB4SW750mYO/gefQ/LktCcLgL9flpqRaQjv+Z3VCJhrvSt+wFhLKl/jqGG
7VYfWAHjva2koOg+4Q4kd+C89acNZYt/dR+fkHEaVIEUC9hGQ/nJE2ICSDY4SZC+pKE8wocfV95Y
HFp8Sz4isVGdV4zNvh9f3187QiXXuz0lDvT1/Y/iIrOVLfTUseFWYqvlSyi8wpEQPnKwC3WQX7Lf
aDW2kmbnYH7sYx/2KmP/RlDmaB7zMzmf0FrOAar41G/2ZRgKwla/a4iKLByBDMWpniHGKyykghK1
j0jvbS3C/PUEQ7NoaYTyFhy5cRoVDxjH5llR1P7OYNTYpLaU0yetXyoksdOWRA6Uxa3yBxd730Qs
K9awKNI6n2png07CCfN5cGurt1gGB8UxnTKX7oJ1PiJVEXjb81F7o4F6PAyl+nD8dy9A+jfUutim
D+JNOKVbcT8yGrrcJ2NiUCPRVTL1T5WYzRNqL7/s0SbXNGmZPCE+TMe1/8jc/1ajuxDqglF+EBqZ
QsyQXEASYHKX3049oosGGTQb9skomN6/Ba7KAq9YrmuL7PQbDS2DCbCUFY0FBJ4AoWk2a2bGU7fm
RoO7ozykkRttu/ThI/7Dlmso7kW2tzIoGXRqxOJ6GuTn294IqVHJE5GdrUBNgTvREaZCu4LkrDui
kr9hiGzXlY7MCR7iABJz6yKDlx4zn79dyCO0X7Ggwb4sXPi+q6DDx3K3/MpMWFzFGmG0a09vbKOj
MaeQLRpJZHNk7RAIDkAIxpIoS8nZgKkHHpS05oE91V6xLcAUN5ce6f0qDg7zYntWXucCGvLCGHOm
vDvkkB/hI0Anngs3JK6XaEAcHq1LAeUElo4bEKnzEou1Z59bbKI3yfthqRJ17etsIrd02whoEQwz
T+VvwX0EDePMtRBzmV3KSMEV+IwIfSoQ0bUh9b5QcY02ieOIgcAMLl5PiiZlNu4zSnigCvY56eTU
IASM4A62QykkmogKofvdDZbw0PsoRY4YOPjC0nzFVMWG3BTgSordzjj+B2D9PO2+Nd8RRCSaHaLN
Kmqdd+E3kJ/Fg1SRyouDta4kgYCDIYVeYNSeLggyW1y+AkrYZIPFmrKGNPSaSDpdzi/J+rnO3Oo4
NiSpkvulbQUP5u43c7cUxdLlIGT59EEtjRUjmvrK0d/zxxJq/p1XSEJ1iTFPx7Ye2Ig+CYkClbr/
PDdpx3ppiHRWsh5Dv0BAUjlbgodcZqqo3KaTvR51+DFYf7broD6SEYWfSl4UjSiDTCR66JcFFHrr
dQVb5oUbXKPZDDKeCWrDQoXU8rBxRcd+KSKv1G+hdSRmC2JxewsJ8cX8+yqp6zEFx6oljHgSiFZI
SwdzZ6uSCSaPVRoWVTHObD3/QNwLWNZug/8XmfUyqj19RyB3vbHmJ8mQtTAh1SpC7Aokuw2vW/pb
2myY+BMl7Ss3PZpdsJmk9EdfNY/uEDUBsR9+K4Koj4jOTSGwIbPzCFVjkdjhGrxKTUb18FapEAY4
R0qKR7yoG4Jt3Dgjdc0CSVWK+Ito/4KWxQIYbxS3A+cdN/OsZyADlaEicNxOxD5in45MOSHySlj8
tnLQRAgvMtYg6lR4pccLUM9MNs6WGdMPc8hNa+JvrsEOg6ELtTaQhRFql7X2xcyzYogkmqXKRnMu
iKxImX7asqMlTMTRGWGNRmRUoiZ9iDx8CJE7sh+2sZ0Zs6D1FGl7GJktWJn1FS7z1ZVMYgE9nyVC
cMawSqb4OFoEaA5LUTP3YUli1AtcCltinUOsO4D5ZpZJgAqAwbyucOXIrkn8+B39ikZGNwm+y5ZG
ZdtZhhIaDIR7TqnLaveH/sJYm+279rewBYswKqNuPnsoCvwxVUxNiINtLzoTtJfq3JdWv97ggEgO
Vb/wPfqbEzgjQNZ+eAatA3hProKUasnJ7/hMCpWFpiu/37E9NZaEF9f3dzd+HSO2mgaQBWspKrCT
8Q6hQFLuVYKk/jVIkiHCZCnsO555lu03qJVp3MycT7KoqKMd/rqTZFdTBXTxEeEHoogPuzutiP0s
sd15QDNv8Dlx+Oy85VE/aqz/eEIJegzkScHdp5Hu/CrHKlemVWmCrS0hDE3JCXEgvr2DzBzEj1wN
SWwFV5pdq7MNUjsCN1wNBC7tVoaJaL/t4EyAAz0yg5T63WD2a/K/H3q+CpeveFirVqWI8tbma1zR
41qfooFLfPzQVWj8REyd+vUpJM7mNqYR0bYkEr4ed2iPZ2rRke6U1piVq6DLfEmRoFCJT/rzX+//
jVLVBpT2b+8V5OS15H9hP8uGvT+WcbTaBqlOBApdQCtZq8vhDLYfNMsVpJ9ybfXeMZxKq9zPezvu
CKR6dS3HXRP/b8j5MwA22qYXTQWduG74lQ+9hGOmZXaSUwopMNjzueH46bNAKRKoiZNl7gHXQecT
5kZv6J578Ph+mJ+P9cCmW+/niEfEUn955Qh4TsyRzHj99O/MTurmy686nlQcHyujfKnIV2flaBYY
6nCpTOZ4p3ykDKyPrPyVN0gbXKAvyh8Fu1yHphjiRLJL3rJybSu7pkQttaD8JaD/N1ky5UC/o0lX
wZXOJ3BPAZAyntYEMoEiv8QCT1VJw696nm6CbxCF9191lRVM+IRouCFvvmWWsIdo7O29Pq733VUh
p1a8pAWd9cJbs5BYuz5DMu8wCflLszkCI5bv5+VWy7UK8P+WKDjAwSEQiJ2RYacJOMF0HfKclg7Z
xNSZ9Mra5XLP3A1TE5/n+MwWIcdYD3E1Cz2choUsAsIm1kFZrJ30XULdpJp6B+m9o68lHmDWm1aJ
btyj4MFiGHKK7u4UWEKh9Th4KPtuZKCxLKBQ2J/twh2mY8ki49t7H25PacdeQRzqL7PuQumKc4fx
PTdEWP34sc6IzEoWedXqJVQ8RYnZL7qrvSRfBk2UQo81PFRdgSLAQHSd7rug1BGZnQgUryzvEtBH
9V+7IE6+S8SjZKxG8D613yTfqv8HvZeNC1COJ0bL9MUCUeMlNymAs2IKHCzmORhYTw9KUMV3QKJS
sagGqAMusxZKZfcXVBg+d36F0vP4GGp8IilAlG6w193O175dDJfJOG3sU9iabq2eQLNa/jX7s/A3
IAdI6/o+KB7z961fX5E+144N/Hl5Ul0OpCMe+BkRmct4e9GnQS3Gz4pt4qlhsHmiWQhH1pnR1jhe
g0+V5riSPG0w12H4X0RnYNb3Q2XxzVa3ErZxQw9RIrIkYRnHPtUJxJGjMxq9wzFGtPaEQ0KZT12B
SosWnSIwM3dqGofSJK4zGJGbURfJ4TnYEUILn7n+b1u11eNATQnKvLJPYRVk9wC416sN2rXgJsS/
ZjCuCL5WSRWuFvJTiZiAuJnUQ/ZMwF9TmrtEkUWKnIfSVwuUwa8c+KkjcrX4/pLnH1JV0lSEG0KY
LSMiFoZ2jv82zxYOfgqYaOdkke7Yxbwa6x/jd18LFM/WZexhulvrEXbn7jQrX5F70EVkJqISQB55
fqy3Sh5iTq9+PIQF6JjZU40rW9PsYwhEPrxagqLNnTcACsDk2LysfGEIa6CeIoZOJwwoqKgRcC10
gHZ/QGuzKSkE8m+yixaKOUPlGE6BkjNNaS4V7QvnDjaWunH0yWXV7cKsq1WxsTaLrNbi6wo9X4zo
NZSJgxQDG8Nf+1d3GlLx2Hc2j+79bc4O5FQyxMwdl6WHE7vjQ5KAQbdRFTXfplC88FJvCb/0hxhf
RuUIVraPSWsKDTiDCqN0/DkVtZFv1IBHZ1gx24fNmBD3ZjH1SLBtqd8ona1rXV9z/dm+J7JkBKyf
IK68oTpr/mV6MHoQwZ5zTdcNjZYORXygaMcbSsmkzQUIe+eYp8E6oKKBfhIEZqcmsEDdDeoUWnfg
hA/4DDsvA5oE+7NnTuqBeSKtE+SEElY2jm5fSprnIA2S10VEH4Gg02OWfU1mb6W09VVhr/W7Tc+q
EcjXr4VheeW/Q/Y44z+RxznmWjr7T4VZ9gPJ+L3FFMDZYxwDwdkIOhDjbZ/jVjw7blXAsCJtuqCK
QskTL7LqLHQ9sUrI3VvUsIbyfZjNaXRTD9jrvpV5y5LvIrFio9H6LOUo8sCNAmrvMaEAYfjpunI1
oWm2VIV+UDBAhgTSgZdDiP2ieFuWKie0QKBQvMABHi8djbCIG0gmdpvByVe7aXRYynXRF/tuN1sI
mzBSoGD1UlgyAaDZ3JOahcwETtfv1b6a0uaDxqTSFdsL+x0PKWRj1bXxXj389Pmlto4ZaPPcr8zK
W9gLcce3caAhB0gWQN56cAY3WP7eWepzGTJdVC294btFB8jFAF5Bx04kaoJiKH0eLyLelCvG9e+R
48x2MmVVdZ/czTt4mTCfYYZbm1jFX7XGaQWjHBzA53fXgLGs+F12o9zgj+W/VLkJZ+XKPcqXT6Jn
Tikwc9c+4jBm7yOdXzNEfHv2LBoCSB/CtVrbCoH9UH/0MbN9mBjDimEbAfvyFlHCOKgoNwK3BdXS
EpGmv0bS5OaaScoHKC4evjxBg5JnVyQL3JqVgoqDdb0kk05gG9dc4kmzgWgItzEsZPeD06Pa0bhb
Ykgf32wny3KNX5n17vazBwU5shYwH0t9mWxbeTkf9i51/AZUBUhCWGD//9m/GTB8WPfOXwWNE//S
z4OsZ5aQ3bGSzNFN9IXAW9o0eGpySIgvvGDMGePBhMw5N82tWxzTxnFz1rA7cGCtnBKcpHMQVZvi
/89pMAjan7XwSB52hbqqRyQcrWy8GYjGb3PCKMfofNI/2KFtWYSZT/WWbZmS+PNaJ0ppgZ/agOii
5mjt6N9OWEv1St7Xv4GeAo4iB6CwRvFDiYbKObLTKHuBAfjAkOKFruOCFJ7NaneVIe1UsFHdBOOl
etHmbiVE9cbkebgerqDMDh81vukUGD8J9IaFdjh6o60fnbZ4lwTUZD7nmy19Ce1B4xy6fG2VZnUU
/6xX8iHL8unh9r4EIlNQ14UYcmVHiMHBTiGvvFOvGwijX1B6Ot4VgJJ22w0mKcQ7IaCKbUnyCo0Q
fUQdJY0Tm96fK9XenQUIr3BrU3Z8aTbd3zjiUHyJgutNixmK5QlwtiiqvYHs3lFQP2ukmUGei0iT
QZu/kxi3s5s7OmyD0XYFM0En2qeyB60ROr1R3kSWd69kwZpCsCWag052uAAA+0pQ98+bRJNWVbbR
5azwzWYKdAZA1DLcGnYvwc3wlYA9SX+CTor2asnosBocGfOkL9YjZsanZYtEZzr2Q2PlfjsTJ4DB
+wT6x+h070zCoVuPHgaBNrUQjq8cnevU6p0xiUmJPM91zgjxSWKBvtbmDiMPTzS5dZ2ZU6ogeAgh
gMHHukC+RPk+I3x/inReHUuE8FZvcUZz67hCfNbVLKzUcWqkAzFs1JFywvS69JjyDkhzGHtFIS4V
9AQss7fbnmez13kwzEwy6TPLRqskRJhD38s747tbbaOHpqOMMfi/MRKcVQepRGxP9Ztd18ICCmRY
f0YIYFWIpBraG96ajWAN+evW6EaPPQm1NSNy6lt2ZY6ARKZt36IsPZ4NgdVe4irMk1kp6GRNtsgR
oQ+K2AdRCkeVDQMYbonr4XBlOpoUsRgvfcGxnZVZjELfyJbBBgEUihB8OgxKwjEgo0TnzKRC+tGe
GhmaauiHDiW9Wl2vsXmbFfpYzUknhuYdQuZmu2TX8PNm+4wU7oBqXg9tFI87phj/AH1U/70U6hEK
T5whVcmX6yYMwXGGez7acv55AijGIXySmJpxL3APF8HtW8gSudtuZtWPaZAPWqdGOhIbwBr0XFdD
OIyhVuH+g6rGU2suCw58FvuZjHUNACazrd3tM82DNxylDxQIYCTHz4ThKInAGRiVxpOB1xnICdan
XIX5QJhas3/b1sU84cLBZHVYQSpEsa5iuElQktZgJj77QoVAwLprbwiXQxn3+xnXVtzpJNFTNmWB
Qq08D2HwdjxQVGimN/TA3s9NSPF3tDghzxxF7UeCNr/+TUKIYaRCmAqjbth75X95DHn1En6EZfxG
eoP/G3T3Xo4hf6fu9Oj8q+qvTpK09MKMK80Uz+3MbyNbwvmqsjz/4MNEALk73dGHbEEA9E/WKGoT
bp6xbrU6wACzCF+clV++G9CASLZ+iHSaYgJY3nsSTolqh2KWa2mTFdkna+sxOZyJduYGjDL8dbIi
qeP79rTkuLNiOWQOQuocHwfaPB4nZvUxrlwDwdxauSqdL4i47lUvvOBxAqLM0PNXctATAkGdALDh
517PGNfDvmnFWp6QVRkVedSsWfl/WCvUoZ8q5OGIDegUKZ633kUQFpuG+pVUYszz/Exa4H5crN9y
sVbyd8tiW/AiztQRzhDUzn4u/jcXCmdxR29QkjCfhmcageqG08rA2st3sgyB03Mi5rwQhYdISaX9
MogUgoRMkh63OrUKMDo3GO7nSP35UF5x2/fgDTVElSJIEqtRcFcvWEqEufCRDHBMce1Axqw0AXbL
MiClcbZsQH/V1XU/ebr/OKdcIcYbJD7DKuZE+1PpeBzaHMzm+3ez6+lzWRDhOvgXvMgqsNUXUIY5
qdRK6o7acBNglGpFOa+2JDpyUDG/oDAxIzrP5IID4kWZHP1IrSXw+IgJxh15uWI4/Xj70Mi4mblU
iEB2jCeiybn8qN4seI7T8c4Psvme/1OQtIyMDJ65vn61tBD5d7hoA1UW79SdHgizST5TMkWbolA6
iO5cQclx0GAoIe1lPQs71Hxv9Ami52lSnLmowwIwaW9Q2/oeRlW9EYRB6l4gbMlGaAZSP1Msz+8Y
WUuz2/fWqjtOmh9qzI1JRYnIeS+1kK/EFECW7GsgiWDnLjrbEq55uET7G1qICNDIymUx0XlCPguc
eGakYGZyQQ5WJsLM5TGi+7Wp7+V64qfTaQiUVxKBW4JxmD/XJzuLRAAyQqXqtJhAxn9q5uTzL262
553O4sIZUxzac2ouTY5m6TqROcXbfHRCaU9asEjMQJe77dcfAkPOA3J1Y1Q+dAx5UKomu4/+ogrJ
HiScqR589Q1ZRyakxNtxoFQL5dephvaeYI//kh6Nkci9CO4Mz8Ptm1IjE4JTv12wDH8rxEIHCyfX
HL/vMYkc6rsPpqbaCCLeb/t4TxZt2U+56mQuFFahX+SrvmTONf8flfXlKdPUfMuyz7rzUGqk/mwl
penAryNwZBTSx70FhpEGESWwaK9cSMw4XaTuphxf/irIAQw3u6O7ZDKrqzPu5oIDuFBUmCb/TotF
IY8E9UQRbVS46HPD2vWF90b8GL8hmnjmVpJReiRBR3Cko03GGoPN+Qz+xZb3XqXP3s4G34JrRtqs
x4k0woAyLfhonUGcWROrwB0DbOBOOecnH4AcegYr0M/28MKYEdhq4Mi2cKvIb7i6UBkPkVMCULnt
VbSTpiQ9vr/y9W0MAan0ObJRH80KMEr/vPDlpraFzbC+k8HuwvqMj2P/M6TmO3/f+Cd73UxumDpg
c8acpZVIF7Dewa7FmdLJ3LqZP07mCjzaYUGNpqrAa3t2fVy8N30a1JXPRK89RvJiEAI9ToP7QXAb
lTLRXCeih83xZdm01zQU/IiSz+FLINNsmf3fi7mHcLnPm9DljY7mD/G/G4eMYEiZXXhXQ1q3Mvvc
YxIvMvop/m5bqh4hzYZuHzgBbyugJJWAkq1zua4Wt9/dCE6zqq+XnDGaWGTh/ihkQgBI9tVszpJM
wmzKCTCwfBQsoOHL0sihcKpvqY+r5dOZJJ4Ajicl1kLinq9rSofWo3R9iShKkE6OqjWcfvcQ/X65
ygBHaVz8vyTqi2ZyCBqDAAw6z6sxf4Y6mL/vUz6R37NAEgQx2pKlYF3HxzHotNFb/ADZ7Ld61kl8
YyJ/36xbmCrSNMiOBaoc9h/MA4FOk/E8j4GogcitMn0cUExEG2bnpD204WZum3fvVVoqOrX9oc2I
jYzXY86MbS51ZT4Un98c9pbxDn/0OrIpemYhkWIjko6+p/gp4EYmjT+RU92aVyv9DAZR7o17eZX3
BesLmnEvxCTOulAzYEKU0efS9f+bozyUhiNJdnXrxYHP6dA2V5G3tbM48MBuOh6pgsOBOpPDo+Rj
hAQ7lqEByA7URyPRiI6qmsGUvMwWZTA959gkDIF5DcJCyjERZtvwKc3ldbHSSwj9B+hfeAGvOscG
wel1S6Qsavnzk/uigZSnq7WiJgNTHt+kZaqx5V361yU+Ud3nFYkQ8h3USVC88J8Nga7xeKWoWSQ+
Y1iCXJlnTbf6SCbY/x3M0Fm6TcAQcnmBBRrjPfXpHe9FAmseteJ/86YKXZouQepRdmetR4v1taMX
rMBmvj9tjoFiep3bUQFkbUR73kJI1mSnGe/ZQ2f2aBvGMUaaqakXwd1NpMyP+/oLoPnFk6gQBK4D
zPPmDXAo0yEr3TcTw9i3meQaZqVp8ruHBTTWV87ttw9DSC9rI/1K1g1HvN0m30I6GDckIt/xrBHx
QZVAQk5Zad0KpmBlJSeZw0qwqDvCzcCkWYw4CqbTYh4VWTYtgE8U6R1HQMKxgpwx8XXceAsTDeiH
CLqsxNDGu/kpuaY7a0XzzMAr9UV8SDRu10zlX4WdCcYMVAgffeLHiXwMowQNpQpFxAvPoQnh194d
0mcCaBruC30TQKc/NeotRMehVhX21dazhoyQlSpAPHg8JMtxXNYWl8HxScuaDEvc7KHUXbMHyzB6
IUkeg20wmpndXD5Slhxxs0+iXo5xZImFFNmEAYbzuRtN52pbs89u2YgCKUSK/sujUV1et6qnYom/
QrS2WsUgPNYCeA1Jgxc7buairMqra8aSI74HpUtEY6H05i4zZZsxA7agtemPP7p5X4CW5BRzpZ+g
Ur48rGjYhE4M5FduKBjYkANNKeOH0Y1d13Q+GexkRwCzZH+6Eea4TZiiCYMkjRsPwWkP5irZSXlk
2cfpQ2hmZIWJwSH+xm086m0Pa+igKEg4mymIqfW/LjRC7TzzeIV2jN4ew3RtKL50zertNkHCNj7J
rCQDOzywven3xc4/V86BSEGc0SCpeuNGeuHUEEPE/hpsNA+eOybjgVTmFriKs1O8j33iPzovSjgd
owSqteSBPS/4g2ykrL5nh5sxieltocZis+4xexHgDv78NbSmubX7uD5duskXCQzuO/O5q/gr2fdG
q7ek8FPlyJ3+2EukTfSRD23l/1UxRGgbFI8SlILOaFcGLpcOiIplRAMSnHoRDQ6gCSz/vPWmjOKw
2+0BGGQMuS70BkWflxq5mR9w8AAyoKcU9luQJ1F26uJJdYUNzu6i5b1XNH7t9uPD4DG1dbhpwGnm
8VnW8ubJP/k67xwcjroy9bjYCt7rPSlX+yQBkY6iT6xH4mZLvlpESCJEnwoEAtJPTzrGHiSOIBSx
KjbRIbkXTdGZ5M3OzKAR0stPgtcHu/98kcbF6wJkBXdNQWdcg62fQfUWHtEA6wVAvaGC7GW7EP4S
iD/TS8fqL9nERLK793HI1V9SPhIb4o9FOFnCHJUpsOpw5jd05D+Vk7bhCzptsxOo8VfdUWPS9ibu
wWIf6gzqOlOLovPPj9h+9498L4tU5gHWLm0s7UOyIhLQPM0ZGdHEzRZetbWX4fOGGbIvXv+41Lns
p4rO/UXL1FHoqfwGcbu9XIjkS90mx2L0Ly97PxsCeUlg5Apz7LwWHFODNwoWR/OTslBxcfWzbITk
0zbcg/g2IaiMvQHhQAioWeZBk4jv91TsPIPUeJE3KpHdLzDzi8Vd+jcDWvJeRwj8gX4h/tXMWHVr
G01lx2CxxqQaZCadUy54aap7jdjE1pGnPKWnku8zJjA8y4oUxS3H/0UA+fAuCU9eAsQTr/l0/7kM
2C+4VVlqSXBWkDeyKSM6hLAVfesp8LTASu7s0vBrZAwk2QjRnIhk5kIGRCc0Mn2X/UBh36WDwbRH
cPLRur7aWGIWE29shWjtaX3ogK0LLhaj/NgRlOTCgu/FlOAfeQFF5w3FUWQStb7ZUhHS85VNrz8m
IpH1pmNd/4XXjgj7hNN9vhuJINRiH06n5fBq8eC7o9ewodXejqcN9MnUYxYCyRz911DgF0sKfVYe
QDi8wj/+0VE4X9fdXGB6y4Yo2/2ov50n9c0ymOKHUOKAKVxKonXU/i1yV7GXQQSnNUgdpW51S/rS
mTTCOxtBl+f39BrPgD3MVp3OYxjskI7epQeSw6L+lcwqyaq2vUZXcYaGSiwcHW71SzMMsrIMc0nT
z3qYHC5qmrt74d2mLLugtJaRbdGHMPSfMfBhv1FjzQjdDP9tkhJllIfWhtAIPG1mG0JiEc+5Dm07
MTROBQkK+hwQYhqhZT+UxTiWgAnj7WdMxxWUWdzJoYx+9ea2K8i/ij/b7U48Q6QW745IQn58d1+A
8GUbBjaUoceQwdO6lZxggrMRHqWJLwc34+zHjltzxtVKFASo+NlzBs4IWfF9ZwtMJT0QSSZ4tfbj
Etv6XgpECjiRdwlotmPJI7HtDLSjLOClFv8+58jz+93srhaAF/AjQ7pIfI8hwTy5A9LnYYpO/Ufh
7MhkFoyVSAhfmCrDPlP2fECrOIjqDoHhGOp3d4baCSTGJdxo6iUGL2WihfOFvPR5d+emhseoOFrA
FgCjuekpX83VIydzBLT8+wni01wpM8R/5oy6NTmLKLmg7qLgBVmSZoaenbqqfxvcVYfdgPTCa2r/
Abh+ogSEkNlniNtosa58BCeC/fH0b7smLiwcwp/MJUKMk2GCsyIvjqcMf/66HAPsrDhnPp+E4v7u
8x6Yki+eMMR34++XJXejH6EbiWvPF/pfiAllQi5620mo2l5Y8d+7TYqYxt0BSR6Y1fraiFzbmS44
BAEYQzS5y2FvPpxJRa/ULv49oCHXQHJRDI0+QyXPzViZKhkm3RbbAlKMsQKHUcq623Izgx7NUqB/
nLBAcTRl41FHyXGsHqZNiF4Q26g7n22Z8Lr0GfVcgnCP3LrPXUmWQKIwXcu3+0tS1sOalENO3BLP
JjT8iNq+QrZoCwhw7rGDh+YxQm0sX/D0vyUaxcuMclKGuyXoSNDlajOpbZM0S7wFjwrTJeqBM9sd
wUQE/t5X+1ReEOKXuKEC/+DqTUl3qadMK4BGqd4MzTFM/bs5SDJVcBjJlSFnx38jd6a4ORdYjM3z
a6Qhiz9hR5Czz6tvsWsl2NodClLiqMuGFtE0bQFMhvdw9JdJnZQ8dQS86I7seBJHDUxunCc9g4Jg
wBZdNm8/1wjSrcWKoJMr50e2WW6Mq40vp53s8rH8HITo/iHT8gjXSPZh3Z8zBAB2JAr/KiYXc1Hs
7NLO4+rVyb3apEWARm2Ds0LY3A5w2/DTuW7OfQx8UvebLWlyrwg1uy+IXbVrkL6RwstLdcbe4/01
QQ3BGp4jrR8p49/a4m3M2BePwj7rEzl6vteHyRIldnSOjSPDgdO71ioJodNKyKFbUlSfB1+WSzBI
fh2zAmQNRIRj2o6vf9yA9mt4UDABylpTU7N69JnD295ruvtsMIp8HkitEHqPyv+nqyybYv94p8rX
NDjUtGQBXuHrtCURyUSheGhx0DuS4SkGra01hVLlP6JMkDClZ1yxfcl076vToaoN43xDOFMTUknJ
/LXP5zxf7p1MiGXMMvs9VwoeRNBvT6m+a8N2/xs6cfQDBZjU9IO2T1TT9vlM+MCf3YRPOUqTiBTQ
puJIgEYjOQfVpxpj7N4MW/MkrrHZgVEiQ6KuFG8tcW09ao+HqV9Zvb0TN8VQuwBsUMD1cC7clwqZ
nLGvh/16bRFnkKC7NV5I3EhIMNnJteSkr6Pp4TNniLe6/0xWg29z38pAYm5vM6aRbT68O1Klv0tI
c06S/raYRqjEUrVxhWWuZU0kaZhaMWIensdwFbNo4yfvsifBPhpz2mJDW20ZGjtesIDcZ2RLGeHZ
JYuUPN+oaBhvPpU+CjZtBOpBUGtvCf2BYzzH97CdUX+6j9cKs3yOaskIncoDbgjpbOELDSImbuQv
NgWJAQVcSLnC0sUj6KjBWnyqeaSI3CmivI/blNTPKo0hBpkIIelwtOs+l+clYSjTzYPDkVd6lzcp
5BaapPf+JZfe0YdqqcmP3I1StB2LF6UPxJ6/7lSIzomPAhLnAjoCXDPh/7athDDwgDlGHaxLi9Oe
8+MftF/sUOPoh5Kux9tIkkkJIlmVUG4q+VapjlKldNBPMkUUiewU0b1dFNLvJ+cW2k8kk8Oc4G+J
372LdJ1dHK/2aEv4y5N0lk0jwQO4qUDvgTjzyP8X83wafPBUJi2PGp6rqKpOim6FEvKj8ffWI/WA
5LPActFg0WHtoip77iWDcNPaVB8k2P0DszOac8X86JFBaHjZuZhq9pCn3eUvoxoX3oeUXz909pL2
lJb746tYBVooHvyVGucXUz3ob3ngmbK0e4lPsIq5xDOZsulBy9u7uSLx3zde5W0BEtDj3URw9N8B
mgku9k+e26/VaylMMEhxhdE2AD01MJLTOX804ACV39goK2WV+l5Zw2so5S0864FyHN3LX7Mmjss7
55v1dbLgi1sI278sZFMX1V5HMjPbz8jxYDByPsfXFLcPM1ZJL3vIQe4YbusfQfjPQBC1YKEUPZbp
1ifa6Vk2T0DcgdkIwyVUzYZjR9oFs+IRPhFU2UzYo7qPaw/Osea9Aq8ITSSQWYojIwULQA+j5PGd
AIbjkmVBIfzS4X1T8eF5/U+JbPDjBBI/oO8SAap9+eS+bs3Ihhhe4UBkJfY4DRzfYmVzZv0kIDoA
8auswvkHkkP2Xqe1aP0a86H0JzH2je4vNPtOB54VqnegoUz7Rnp0JP5Kd/C8MQcaNJTrZQ0UWWPA
HgY0ZkumSsWZbKyyRnx6B5chX2Gzbh1RfXjG+2PsEVrLssmyXTevhV5CjqbbpIukCInAFTrWCW1J
oEnzWFT0dVS2cZLJ22IfVvxsGpJnkSdY3g7hWFEi5VBqXa13njYRemlI5asySYzZpY0NKLpwu8k8
5Vcr0PjRttCBQY/tEZxRke5h0z0xXWgEfHXIsg9uSgAsUtAQirXxw0VSD4GVLBeE+A8aglzLzWDa
mcZJwgNz8+3QCSuV4AqGrceGJWAPHXkMiv2E9BKDHhaqbm4SlOzaCO/3Bhvim9A71csx8xzNJPGJ
8qxqFDwH9IuDgDV7cTk6JX5LpGXJFCE4ldC7zyNftCZrS34KgFibu4dQxMgvvfkAlcGh2SAduL1d
sel48VOJZXAIkusPM3S3TbVw0uRfHdk17nqY5MEZnxy4Rm4QMR6VXRm3zgdVAFA2xbcxpXqRSBKn
0xjDMDSyLf2QCqD+ci9LSKrxK9Gq3OL2N6VVv0x4utlPzA7UaWnoJzLeZz9F7iRk/SdMH8hf0E0R
tDTZIMwZDbAO3pFu/Ha8SebJjJzJbv/+adzY5ieBlaJLjfByhJu0a3ukVlI2jU/id43kM3FdZL/j
LJxTOgOBDyji6RBXl28lONuqNVMipbnJ/2GzZAnB4AoUw6P3IlhYyEjglZFhAx2BkXAxoTKu82J0
8/iGXsdSc/EtGCFATzaOifuuRF+uTubgHWrk/0xPdguylU+qsQ2UrQhihwQ+kZCLNAk2Q/L6U4iJ
AEKsjFtkQ4cjosEmAv6t8hZOJQ2XA7uv5RRkWr7LwkK4mW8h7uUkNMyBcCEX4oZKW2yUM8u0nqhJ
sa4FNyDqvNXjeo+UE1vtXLzWK7nly+OzTDjJ/+s3OL0EIUZZCLUD/j5mwME6OfxVyOLVuw4DJaUd
8u1+ASvymHXnjLKo+ym8PjlbdYpVK2eUx4KI4nvL/mRZQ3W5qEAEFtg5N+KFqCukGdkGJyahTpXJ
SWOM3TE79hN/dOWRtygRkZ1tXxvGQ52SFtH+Vby8e0jJxvkT2YyGLgNj34eGndxzrSrBv+aEcVyd
AhFP1uFXpyeiQxsUrVwubXFhzl6+gZ9FDiOIf2ry0NXiodPCWJq6/wd1pjLpr3atA8fSPIcEDnaf
99FVhgzImcDJrmSoD11TGA3wWtrHzjrPuUrSWWJomuPGDWL2RF1K9Xwp9OQEj7tHZKjjCb/pwa7p
8wglGihKcXeMk/490wGFRsOQowvd6VTj/lnh0j/kBqUOnLaBGcfe02CQSTrYctEdv+g4skpsW3H2
mWJOIjCeP0oLAHdlCJkN2y1umSbMpVqNoC6IwgrKo6t24fjh/BbeVoWB5oHJLBmwHzIX4c9vrUhN
/wq2wsb8zb2ZdYgyEwJHSINSkZ5EJ4dq2HkhFSJuXmtZNUQq9OI2NhWZLRi5soWpYkhBFNuqdJA6
zI5o3LOYwn8Pk5ylhfRMaANASHzJjYDkGZioeZ1tcdrM30f1nMSmdnV1uOh2n9vzeLB88h1UbpZh
5N2URwHQoMilhynOCzplLQOg5NXkIfCsGtCHdQdKLLfHi9U5C+Y4ITQ4E1DnlnXE3oRKqkPeQ0Cn
fH/CPkzTRv33gSTGhfDH1NLi1EqdmfWcDVRG2fJYO98Fw03rS6tprorfD6CbipUV3djwyCIEBMxq
raq7uaXb1D0BRaKzXe0G+0DAKag8ZgtZY/CVWd+8NbCJNUdVCIeaTQVuxO4ajAU4jlcqsNccvfUu
ucOcLVRYRtcoa8OaahZsR2NyxhkXPoDem05NAs5JgEDWtHxshIkm5FNcbdjTYplGwPA0oKBKbaM4
m5JnsEf/+3nGKK5yj2P5LDBBKKA3WdCFCKPu8yAhltZ/yXL2uWzFYv4Rp6c3PSjTaAcbqyEfG+uH
tCuL2eDDJMPSbTcS2ab/8zlD/FDfspTkF4l7gleCWjrmLeWk21N0Pe5c1JQSDixepo2CbXKIh1Ep
ngdDZdlVp77bl9k6NyY61yNspNCkBJK77MPkQehXpvQNOrfKfOkAfpWnTi1JmlPgOwxw3SFXq3wd
ZVmtetYh4QmNx3U0QeJx9ITDgmAq8uLqVlu/Z+YBzSHFZVDP2qw57Y6+3LzMnsJ5CfB6QbpokCj8
jDqSzKDjnuNVPPMKIOQAg/zZ0CIPPal8j3pAekxRzb9A+JvsHNjeuvDZiRkNZVBqfAkQGyYAVFBY
G0hRN/wLpvxsOBixHgM4yrpsBbw1idLrc7pvCdTUFb3IDx+4kUmf9VU9smdlxrzzhFiuZyOvbmZv
zf39mXX/sEMxSJnybXAgiyRemPUhjM6hn8UTpVZtZ45cH8q6v1mIgrLknWu9v8K1ItkP73URvKJZ
qgUbEl6INiRixDkAIc2l2zeKs+84u94N57FcleDMeh25rmF5/YR5UFc4JPg+2WiKHatg7qaf9y3q
bkW+sU8o/O/HjY2ULIAoM4OVzLY9njVQuizQIKaAkmY1vMClTC2BznneKQcLUyS6200cP+c9VCUO
mVqqnlgAQXncn2XHbSDhp9HhobbFehN1/ihXRVp+3GlGQwSBUvkEfOSaAnxkfetEviZA1Ivwk51a
LOEdHeBr20LTl6RzdOEW7eiXb5GNOTNDIzyxbtBordsvze040s5bh7c9rSM0EZN6Q5PAsbfAqQaJ
CsqEV1xdb/bqX2ciQMBgLSBEnYrVXSTSisRgN3ItUkb5gofV4FwCb6l/c7n/YEirlOdqBVbODN0V
VJMR/xATHvD1zJdNhtTAQTtv42oltt4XqSqxF+LRY6fHKLFsfSk6PkAM45rqlkSAu3X4IF0R7UHC
U7AEYUdqYM+7G2k+Q6oh6mOqDVjAqHHD932Ze4DUTTYXk+Se2GmBN6hNVUHxxqmbAIbT9YFxfcMa
3bvl9168jUX+o0seUvf85dRO4X2l4aEsGlLCIXHzOgK/sr/s4vdr48VtB7Z3HLZ3gt5+t+uLfPJ3
F+Y/Iv50A6yvXwaW+qKy74uFY+yNJbyHt0iLshuJGDyCtOeqFNgsqG+p0ILorT6c9vsiAfKwwslP
XgHPmhtt5sqHxhuUPurcIKZOkEdcS8AauMmeUTqkI+8vbn8BuKrVZ/+GBpmuqD4/2XwYmE3spJaC
xLp2Gw7663QSNpJ9HjDgdhW5AeGoMlVUoLCCkIobbMFJEIwFEBzs04R5j0UdAw2LiV/axLC6cfQf
CFaciDV5x/N2JNxwcIc0kfxXyu28qRUi8DuVL290avCsVD7DZRR4vUgq0gBkvWrJ69ER7duZSIrs
+cxWjYb5cOrXH7s5/3gqu0WyJobLCkbFE4/icGDw8c/tp59Zuzu5TYgCP6b9HtonpVj44I/e661c
EHxkGpKraSPHZYbPQ6sLVa5VAFx11UU96XwTGYOYD9MBQb1FhH7CfbcaBnHDfWAhc6KuMD95rkCI
SSz9WJxmkuzQZEa/SQjFpq1OLYnfMRtdj6zhvDY+znzHSTh1cjUXIyvXRK0eawRDJWAE5rCAzxoV
kIOKPNGiIIQa2JZQYyR6jKdBophnhdNHQo3klIx3YHb0igrLYFYlUXU9JiG6ElfwztgTSJjNF+uQ
m1mUs0vU6/EST4wnQGbxScJ2n1kzWFOSsxIx6sIaw4Lg9o2tW4vA9kxRTLTc9kbVqWC/I3eXn/Y8
3xAKaHfoMKRx0LToKw8Z0bzYaHitmeNzaDcn9Gi+3JaqI8YeNfxHOLuVRVQJ7roke0/rvQ/qOxCm
ag2PoUgTW5ssXNTaANu0gVFgR36rorbjlAECSh/Sfl4wU2C2Nq1NmR09gxIDsGMMUerUTPg7V9Ar
o4QzIg/Q0ZiznvJ0HqO2oERV/kBNFdPwGRORYHBr0t1tPiY8armM+N5gwI41KTv54J4tkAs6iq5F
ZISoW/cu7RNI00S8wobaYuwLzSMtzwTMF86N8DgN2ZviUEkIj3IzVbE9/72gSccMZy+6PqWgVtXo
W/aT7ROtwQn/Pa9OG9W601wKUyNQ6nWzo90sTDgu4fp40K4NsRFHPB7z1+0DWOeKeZPOQi7EahFF
ST3mypmzrcfo/rTD1HhMZUARpXMey4f+9NiBtpPPR5gLoQ810qHAL2CfB0xPIPXa98UjPH2OxnSR
u4gNe0rT/cvRUgpzBLWy5Crz7o6WAkzctXHD8WteVrgWg7EGeXMTO7O3y0jtaJ8u8mevhfyKbNK/
3Ztt4yyJIB3eDbCU4EZpK+emZ73zyzpeRuTTAjsXyMChg1puxBD80uiOZLHh6Qd5dAKHW8ntqmT6
k+OOo5ZbqM1hqqwRFP7wvYxDWlIon9Kg6juLeo6rBn86ueoMaGhYPlkjFgKsKd7uUkLYvw7pwD0w
YlOjJWc8/OMd6ipM+zAEYNXaVF2/WM8E3NJBOKyre2tyIHPVkmzJYHFdyX2illCmylPZ40zc5vKh
waw8Kvn3VJoTK7/6XKD7l9g9cz9S+cQSr5hLzsXIgQ8QsbpEahzXPvn1mr9D9UYoaZh9lU4k3WVW
uAICliKCyKZzanF/4DXS3BA+J0WyAgt/ThUbeX5773SJweMwTxj36WZCx82WXOsQntVyhb1cTVMw
oJ2S/1FqM97fL3GTCnowJc9erZWJonUvAlei5DJ4FvBf/uMzpDlLlFU5OBqAcul58YVXhX1OXCND
Db8lS4aYjNxpeHddp6CaX2YUQLBmlth6Rhmc8I5mAMpoc3q7Yrg7rA0yVIIHciRBpSd9TSMkky9R
lGy9wmJwJs8+7mKoaVJiqXu6Wvj0iHL9lFscLtHnduzKf1zVqUlhHN82LDeRD9R1AnhwR8gHT6A0
nhZ4rR8CwnBLaD9cseZ2yjij9UMsSDEU82ylEF6GunJCZJS2qcy7eEC2QznXEDK1NcgNt9If8gCL
6Z87+ExA+cCeZu6KuIVfhdCCAUMXdT+XOhp0HKEPqAyuWab04Y5HJVip1ct0wgo/fexOhFdk3bwU
dgV38ATju5rqijwTgn2ppFlyh506LTSTUy2+oRe9JClz4yWkUa5T4A79+xTWoLdwxApAFeO0+fc5
T9IlIf4hBFeedVhfPJpjMJCA/66NCwkX+iku/H6seTqxsOdM0pma+f3qHfjgEqb/cxyAXzLyfWLs
wEvel8T746TXOYWI2bjkFiL5B41Sm8VAiPfLduAswomIdJ5WlLtp+esJEjgYwR0UkVsVJq7NuJ9/
5ONk4yb9+fa2Zneu3lFE9F7mM+LeGfMonFPvPBRXlWsop7Eh6CuuweyOZiV8tTH6FdtX2Ji+EJAk
PrK4QEOoHyGdCMK4/y45LfFu3So+ZUS7nRPsXMdz8btZwU/p6KZtCx2hcuQtvsFefC3W6d2yvpec
Rive1p3wcjdL+a3A4KMnmfEsWnr66Y2ZE2+KE6E9dW7pwnDM+BKH78nGfsNbRNINHKvKMMZUaoUa
cKa+4xoZzd1qTAxYdfRUX4cBxedm050pq8eEckTz3RWM9DI/L7d+/5BSfqeMQTn+jxlAc1+kFZ4L
f+2BDNQ4Kp1a0Nnjr9Nx7lXPmen4ZzKt+t//WLyx45FIpBYKejsNfwUDW3O2HOoZzY7Vnxy8C/aU
EBfYttcm/XWsN7KI6WFOafzm2dYZPGZyOd7pnwbcCIEFuK/4VO0Eho1IH89sBe8wBGafT0Aq2GCw
obav0ipE+DKaJliuZ1bPiTKPYoCrBfKcNX7anK1EwkKdAijCfGBxf+pOxxG5Uy72I3Bb5/AXW3CA
LjY519kENc9FMkvikfV9LLuPr8Qx9x9UBwNGhZtxld0y9u0Nf0ts2kCnM6D+/BGrF7vPfcBGCfQK
qxqJ9vzWGajBJQrmMia3v/QmORv6hOeYuAb/YKttpSddB3YbflztijwO6dJA9DaJ7Fp+HiMgi7JT
JmC94dww/RNLt4WOp7z7WfXdkqciJYJ5IVMOEtiiXOGAVmO8S97TWqAu0cZlPwoZPNK9T1r0vrhf
cRcSNVAz7YqyfwBOdh1Lb3IU9P7Kjs+4+lK7BGavOmPQgNv9CL4FmwwKJHOM7MTJLasd+lJnbuVc
/PsZcfdffl9aTcsOGXbSVzLgelWyri6+0XEc7Vbe6Df47QVaOY9oJgFctRUTt3bzpWxUU8OfM0NX
1nyYdXJQiSovScAsK61psD+tN8UoNad5Hb6NNEKZVO6b4cP/erugkr+uTdqXSLKOw+P51j7OOEnv
dLrzyk4PPYjVIFxZFr202MFJxnu+xzyFhf70Zuu8CZfUpP+7sI6Bd718BB+3KIJKX5py1UN6inOW
DiTWwuEex/fbiUfSWQJ4mJDozNCL/C+uHIjzlSbaPBrBOJ1RVG7+9MuJLA7RA/yZUHzZRUxIP0ny
+3upFiqKHPnFOP6J1P8LgJpkjy22igY0d5vqK9Y0cOuRdP3ZroolvW+N20h2Yh7yvtxe/chz+XAi
AItfN978yNJYCyX7FfF8iHe1krkUKsROJhpnDRWke5tNDq1sKyFs5/11QTOxWsNNq1+NlRHocE42
lSSxn+vnKM0OkaW5fETD/N1htl1+cJFNO1ZM77oQIu5L0j4O1BKryAHHIKCBlir5cWUFWKm1P9nO
oHSGMR041rgX/KYaF7vPF568gWEjpge/4NZl2k2DoGmcWLuYT/5GaJG7NXV1e5FqoqAba87/dxor
F0Ru/QXZ3kpvjdfIx5EUUmhEON8P73stMjEzYJXN4iSlFBa9I8+Rm3Pe1kpD74TQzUFt1VSn21IN
AiOLK3myKjnkZBLy+cjoYS2BNr5TyLV7AFiBNFe2CXBqiQHNyQuymDSNqfpCys6KmTNMQoemijto
TB7NKq5dQoI5wgjhhdU7u/Gqpkejz9xmGEuSv2R6L5KxHIIy7V+vl9YT9DwBkkZNhYbwNw+BRUZO
L60NAYaVfeyLxQIkgJEvYEfa7wgSoyFx2F0jfVIGUJHF7uq1Vj0YlZPdLVawrkSOCqK05yarZSrQ
FMpFN1n1kfuI/QgVqtcBkXH/gS6DR3PPAhHs/YR/M1nwad9oNPsiKpgftixj4Tv+l78D1+Tkvk0u
KTTLML01v7zu/W5/FFzziYXazYconNCYNKfwuZ5RnWqiPVNQAaozZg1F/QFYXKiJf4k3U0tq5GT1
rleZ/eSt4rFAU4JysPJvzUDBF67Y2w+0yosIabOT7RYeuhgCjCF7OucFshkfkLRPu++tTZ1Z6GiE
31X/xOdAnRSkGQq6MLlcaN0jeQlLcJ1aHhf1Z29YkD7/OntEzmnl/wlv+1lIw9WhmXxhRko5HQ0V
10lRpAxo0AGki/w982R0KEC4tEHExAzPvsUvDjr5+8le4fJgLEBgWDqciCQo5jYAq3/Y7oqZT2R4
2uWiMrwjbiXq2R9MVpKWoFDmYOPxWP4MvY0TTdZPJ0r08DvyUXm8w5ZVlJfn3KalgQS9zZY4aRdv
YKDMzIuEYxw47d9/VjcVmGeVUzcL+sDypjCUByiBAPpQqpiR/bKQffMQkpUv0axCUodeYfdsr+mA
FKOwNC//CK++nPtzDuAP9Wf4iq6NAOjZCCOKooNb8mdBHhRK+gH6whNK1qEgHkh6zi+gecwy1v4J
dpaNa0dpB3wRJePleybxdGAKbFC2gVTAS50EMnku7igueJeeEzvdBA4nRUuPQRgIwt2FzpWK18dP
YX/9lA8eKXf2iukrCbX//ydMiVhH7d/TmfC9W99a1qmPIc7vMwqDlf5TOky8DktrhuY6WPUgBxnT
gVN0DTtPFMCc4n3Kwjp8umuSqGSSDUEIp5WBZha0kp5ds6he8bu/gZQm2a8bODu2NMxYo+MG4VUl
ioX/nA2bN6OYh0Qo8YhlI+6wCKOi/Xw5/1yWb7uNUZNsk2nK5cqQTakY5dJYfYK57X5XsO+nLNII
tbcCzohgukQ/LKSQ6wg5AsMu7uIu6F3IZSZi5Oq8HRqEx1z98pmk65X0n+t3XIeC2sejqUBKlbvS
UhaYousSDAQKG7QXAoQXwYWT0dl08aQJbHTOTQVHRf8s60RmxOetAh180JcT1z4BGiGox5tWLWeb
IduBEbAfn6VyWqzg0mqmbCNN+c6vPrPqAlxZqhIDQoyxtPXuoaL2UmZ4kyMqddieBvUQpp7Zlgf1
TzaNT/l0/XTQeWrE9VhniP9wN+hsbRN6QUvlOtsnOdqnbL9R/bKEu10BlPzFkN0HwwcZx4C8mgCK
o2rt6UCJWLdKbjffg8A91Kttgfm6tr1MOhE7AL+0rl3bi3MUqz8VH5mdR2Ra4uDwvQhE8L+F6Sm9
FVgcunV4OyB2EuE2I+U9fOtib+EVFkdev5RD+1OKL7SsG0GI3YR6C8DgqhojCj/7Rxs7Rnivo+LM
+hiURazmJ2cOLCt0y0Vn0139dmVs7iRDAYzuA5ERd+mFmc2mIXfUbJfJ2dOjGqyxFvmgZj0VxjeG
6L5LnyjpGU1VukPIUyZkdE/QA9TbTCrHBp98FH9CA0Us4PYHs5uYwAnDE/Ed8wy4MS2njwI9ZlS7
rnrAWaSjQKSfdLvH7JXNaZQCbAjNaizVhYP9EI9waDIwUBJEDAI3eQAH5Hrkwupa+y/9i19cq402
QIg1VX+YczX3o1MOYHKi4CXWe9HYS2VjzaySpImpMBCDw0jD0xVo55ERIq2g2k7q5U1HbReYlTnn
XIIsRgKpNAvHMLIDAVOtm7Vnarz+ipxmLCuNpulP4bPKAIAF/5aBqI/iJ/6XujrOeYrPIRYYU5Ps
khmy6FaEALEJ3EpsgOWquvxr2wyGm7bWDWl2DWhr0c2+GbzQVrIt45iSYZXOwEnBWVR2sYROrtdW
pOuudzrXC8b1YMR6pW/OPQsQHJ1wZgFMhWizEioCZZ4IakRyWpI5mFonZKWyOeSCk1tsbfJmwgVc
PmT/Dx0YRNmUkoJ5dORifm8MFk7JOgXVlbVHYGkqcuC5055kezdRQNwiePAfX6GerZIsdB/AIOui
E1woeLq7y8BTb2xzELNsfCHcq1IlfZV7mEEPt1RNxgskMxb0jj6wjXXDxVKeCDHSKw33LQz0w0Pr
tNaF3i8ZekbOuJttXzB7Yqp8hNCdg4srR+TLTEpI0rL6wtPOaigxkW1/giuioJYpf4rGywXnJrzQ
DfeN/YbEk/gFhxtd4GkTkbN3Qjp6HvC43jLjiHEZvhucSetmrR/9LnbcbxgWlqCoc8V56I8OH4Os
89CHPq393pOfYgaxmfeqWsTiWjfPAVKM6PnE6JzIcmjhkXDzLXTSaqyJnXEgumBknipTGUy7pjt4
WeH/vWfO+U1CcGo6ZDGLGlkEl3EtBUM5YAsJ3YlV4Ptwm/d5PzaPYZyLGQyMiDGPaJ0DyQ7Pwpp8
9u1WCYPKIutVbgbj3bZ905BWL8YNGBL3qct91d/Z5TRlkJ5enWKqXXxXqioEgMETlh9SrZQwHt5K
tVKxnrJ9cf7IQrp/j33DaYbwiB1SK6nfickhnHwW2kBu/mko4RApx/IsRFzpZmdZyuULHcmQ+Yv0
EYlsjCFJ99acLwrLXFziYDBMgFWPNsKwmgyN4tlg5fDNlDRycQjSyUDUOi7Tu8WmCpJD9nlHVKds
ZuNYhpqtWVCqltBWixPtvKgjUNPoUwWaEC3oQnjWnCASgW6k7PHD/0l7icEAycklD4GOeuTau9B7
XxU4kzcU07ui5islhSxXk4B0TINGiN5gdJGk4S/WYnYolmPnncOwqva6T5VQ5IFMih9XNri3SnHo
1/Jd1jlV7u8ZbonE44A3494KZSEB+SaaQN5wOO6gOT5eizoQj6gBcIXJ2rxiZ7zak3JEQrePDRgy
zEo+3cJUFn/MU8HMjvOSMm95ePMeZJzBePVvZhlgTK2+0igTTt5neQXgdtxyGZhhu02vLafwvoaO
J4v7hY/usqNXYyOiT7nzVHj0vvcqxWWI3HO6AXk88/Hn7tB4bAN7PMn8XBzu9GSJdQR0DqKXEOQ8
goNjJXyqNIg8KbEsrDyM0P8I708ZfkqegKlA5p11CXqF1nr68N8QL8nLqRbeSwx7fWX/zeqz/xAk
sYetwyvnz5rQCcy0yn3lSQcS3VC8QEAt/hdXvJQh/gGMCOUZVMmF4nP38v9kRElysNqt5x1bufh8
h/kZtsfuJEYfUTFSCbStHveHivdraKZhYFkYLhCsDrTd/oZvGpzagW600zBPiA8GJ3thVS2R9gsP
GTyIKYHAsA9Cy00nqIoSji1WtH9fcl34tDjoj2ki95KyctNQ8vOFSLEAT6QtrXknbBKgykIMRV53
sS8QYUcFWIvqS/h10Kk8Z5k6DupV6Y7X1pqbBRVRboy4AyhqfSRZ5+xDQcs6RgWNGXvZIuaqg2XM
fiSBGQyXtFlHDwXW20VhHnC9HglrULzj3e9HPfrmGOha31hCdcx/HAW7QUCv+M+PYKZJDx9oECDz
dE/vrTAjIXN1Wa8a13NWax/1O6ozbhqyZ5zpMMdBZ21OHmzKDJ9O9hss/DVC+jW+Fwt0Y+aoul38
BKJ+wLNv/a03+fbA7ALSj/MEPsyK7nrztC2Hf8qe91ZpRXOEZaFsVH8WJhqGYoNNVuzEbtGRNbHI
9uWqZNB8UWYmhjPiPhwjawPgxFWTgkQNNh28zO/oop53VzlVWKlbHPaXtCdueBDkN4Ww9WPei8EW
3cov+4lJ3CRteh6NcYXk36nfE11dsihCVv0RddVt+upLuF9OU2P9ytx1UHBywyw0FSHkSKslb9CC
4djzxcOF+jbe1XTCGCv49dWEOcpos3GJ/vbLzOysnHoT6W5T+JUJZXTq4AMI9/hWaqEnCnNNWQha
ux2uhXW6msqi/9RUv76Lm/NgDfmBbx9Sst4+fsn6YGeooYDDRKulCOO4YpGzOMtslilhqnN8skoe
VuRdjeeXa53S6b6cd8bsv8sxtIS6ye9VRo09bkbl4ii3mfImOtVvHsPSp7EGbOq52S6A5pp2tjV9
e+K4kBZDdFCDx7XoIJK1Yd30nKguLxNIH/e054OlRWO+kovO/W3ULe5jpwB4HjSza9WoFcwg6Vfz
REY/ucd/kuzyQl57KJzf80UscUhhf+dMYkE6rKnOh2nPxs+5Fzk2iNGFSt/DchRQnYnCH3boBhBE
xSaq5OIeFGHG0i/hx/tZiYzM4umQc0BOTc5eCN4WymTLMLjd+7FNbEyF0288db5mqe9RcZy7YLwI
T7AqSrTSK3RbDFSoK5GY0OFA1DhA9TOgzm6O40+WiCRMmTmPsvri6vqmAsUENbBT+fjBoyeXRCTP
wcb2pVtmHWU9ZKJptNXsjzDo4PJnv/t2pzkq1GbArayRHd4ofPXjMrMWsDURg3enPza7+n/EkiFz
SrBEA2dFEZOeG2awXAuZGo+Koy+TeZwHFq03VemWmhLWPGxuBEMguHfqAsAlkGAdt947VUo6XIAl
xHev6ZVdfF3dBICP84K0YSb6eeZO3tIYXxsBZAJ220i7wB9EmRJ6vjixwVPvyltCTCVIRiWkZjVS
+iFjBdPXXGxpC3KNC3bcwasP/pxXTgt9ilz/kbeW5OhnH4zOTzJK4mf89eyl+crInUEq5QMySTBO
fzeCm4f9dX8aGWSN4RYXrptpOP6WM3whPPbuio3vLuY3jhUaBgimVW05lM/0k58IKIdJRZF24JoX
MmzDnC0Nq2+Mx6+xxrM11Sx+F58b85GicBc8fDHuIFKGkP7hJgB8W6kjBLAZupSHH4HZPBQKafX5
UubVceuJHwjAuEmD9YumsoXDMQLiJemSIVrYjy6ABo0pMJbH7I5tHo0F4I/UTjNpIABg4M4qrF2A
YEL6O3uvpGJzqQL990emG/19EGuK+c3QTKtXDtWch/QUbPF26MwYWT/m6Gfuu2Jq/uNnFCv3nBCS
JdeQhcSZuZTafUJQoS6SucKRFzMJGTNdBP8GvocQadQKslRN3nJr8cgD2Adcwzw0MlFXYilzM3Fh
LbV3Q2txiTxUavHg3Jp7HdMV9UMtWc9PEmuPz7R3Ke4F0BC7k+dhl4PvNw68zVDoAM/TBM3wde51
rV9XJ8jNodICRw5CFu+yR/H7STGO7SUpTWaiAW3PIAdneLILUJ3ZxMPCYNdFMSiKszy8tP9ad6PZ
5q7IKpnu2wJN667yX/j7BVuafU//10U+1K6FekuNCMddh90eJIv6sXvzDfHBYh/gZ3zG7vAwEnNW
09fvD8FLCFlea/vmeReWAH9dsER5XnbC5KeKsPcMBVkHEoT0SlO8UPI+43MexFg8Tqws4q3lQXXl
PrD4X40SyzIVLzrbnWOINmkhkF/hDXdKowLBHotyhwThJ5N+hdSJVRF3P33mK2rIO0nyZ4hFVzPS
HzllI25pi6/u9DlgJtepLYHJpzTPIJxUb2TDwatdM9aWKMZnwsMbvVLktG+nNykEZOXvl5ZNxC1o
6fXKaDl5GWbC/gODft/Yxp88+g0VAzK04+799e2ROICNwS66x88Dy7Cpc813XNOPQIkaMbMNTeIq
C5WltOIx3ZjrNF9xDBQeJB/Wihb5NnU4ElCuM5kZFuYwRg3He0ZZUo0Uj1/ahjS5KF4pg5/msSNS
5zipAhIRde910hhFCCTGsmoH9XQdl5yBaAKjcg0ESoeutDdRYLWUjfDxyBEzR08jDSv+5Hf24fbT
RTJC3xHOlsFw2h2PWRpfNLBE5HA1GbEN3Y+LeO4+on94vwbG0JKf6A/WkZ5y+EPibmWPD1Udsns1
2gLr4wegwPJqO0FkScPJXjC/tL7LRdmFd/P6qAAUO986HGWIuhu9HDFt3/QOn0Vy7/bH38TLci9u
Z2aiU7ZxMqexlI/nOjYgNd8cJV3s543+H/NEcccYfi1X9W7cpX1EK5s3BJOlGnybIdpxh8vNh94t
ONz2cc2OCa6dlcTlcRxkox5e/peqdoyfCyLUP8w38a+THrbnXD4I5dBxnUH9zz4NXSuEGsQIZbtt
nrnHYxzHR4tj2wyzgsI5TIlSIJqbmCYHTSgm1/oWdTbG5z1PYHRnZlsN+Nzl3VXK7YQKgPZ91teq
hkc56c8x4lzxSkm7X3knbh7UZkzjA4q5WANwW9obKlDbzmpP6eW2oGcwcc9s+SS7Eluf0cjPXrLD
+IMRzbqm1TYoqBeERDgd+J97VcM5tUD58VFnVEFrkCH6o0K8RxXbTHZTaQLOmZcA1k3TciwHCBYF
/Bkoh0seDKsEbBV4nZBTfsX47Lf0dCuUUwkzFJiG60Zz+F0u9LYR2HHB5BL+RLOSiiW/y/JCj8fb
3KEylEyn1B+8/4Lg4kCbcXh5l5X8daPE46ePuih/DZfbcJiAqZ6hRDNz7ZY3PpImHyCEWV2F2PRc
95OiJucY11UFj4VPAaV7ikObMlG0Bzmw73aaQAxnCSdvuLg5m0wBQv71RQeemasUX9qQ2Qzqv/hW
9/RWEMazwZ0jJOpAUv6RJhiEydzhCr2Yurlqc0yFygmS24vMSo16OVfQuWzr8jFCqMu+Hh88mwCy
4PDd8f/D2YBOhj4+VJ0HwV0Y6Q1sbueTXuVuRDD64IzxqRajSXIo90F5pU2wxXzdi8b7XzSrWcX0
wZw4GF2Dsyng+XWHZmlveQxpz+FSxXEcKf5UZ68s39SzxPWOFJwkntX5KsZKzXqJAIPvRGiwnCrJ
O0ifbfDpHxn5tNsALFdO1Oc2eYm2umuS4nXWHMtTsBNOrXbYIeLebaM1Nxtn3+Jy4IPSnXt5blaX
pp1e3+xa5JWX1a38IDrsvSHoaGNx6vvCPvXmSm3LYIHdUnD1sBRxW+4n+gEM68t0/gqwB9Enletm
KQHqHyn1oGmMjqgXvBJ+tC3jZ5laWmnnjajnwceTp9YLaGDP010vCagm3jPDbQRUKiQizxtXe2X8
84j42kt1pDhsJLTXwxEmM7+L9nV72w88+1rpOBUVQ/xwkmr0I+rfeilfUknZvYF2G1amgm0AhIG4
geHTr4MsOLKOFqiFyM5Nc0txTAF/k2R2Gy0cg6GJHQjlCtkHpHcSFmGjPAcOHsRQ6TVxfS4taGoy
TfP5xWhZM/Zht1odmXFiJZmTKCHRzis487bh7uOYp9LJCptQlq/8KZVxAzYy1FtKPylUXOLKi6d+
BHZ7w/OWD16eUa3+9QRDH7EDyNySDe4503VBbZuErulz6mI8NSk+fMoRNucnCyZY81Fb/ediZAUd
k4/VNPpBC/28eD/aZnvTZWqGq11qx2sDsZM2e0VD1lfgZGd+ihoioIN9n+ANd+Ifzw2b3YWvT+hV
GPbsOluFe0YzlROnKhsKMs56YKThRZwdduFXuyT7nwR4PUjkLSM+dtLeVa3477QRVX6MII2AKqkO
ljvgeV70fRFcb+IT0Y9sOYUQX4MhsgmYmr3av3QbZnPrj7VodJcWO0Ioaebza9nLqbZqATh5S+H8
Wx7014trIqpFz+NI4KYhmNRBjMUBYKbobif1c69ySWkiWKRDH3drSFGEr2Agz6A8I5ctDHsIby9K
v035wYeKlx2ZbpRm6GphEElQVPzGj4zkB0KhQp15p0L/CA6Q70G/iIIdnCNgrFTGnRjSjw4LoPuA
53E1A3gVVy7eb3QhzvkueElH1SM1q93PfCvXGih55Uo7rgtplP/X7ratkeHX0eazNir7OhP4xFNl
pBxP5vOqnGpF64DRmC1Zowbw+o1MpFRDSGxxZGl9A2jehUae8kdBvayriSNT/Q1AWT5UkcivEBBB
DPr3MixT87NNXpEjy5KBGj34F3bXEPDGySk+4NFy+f5/WyKbV3s/0biXmy01lGq8UJ0zKpDnTtDl
BPCaqmF/cOyUqVgxdb3w1baBfY7xCvBrd9rKDj6u2F4DEWJehNbHeWWBHifWGN520nHHjfG7QCaQ
F55vdZ8d1vyYd2z54YstvSm5nm/WT+Cl5tLhPtPNKYx3mUXCQsqkzTm8zTBFAOqASHvLvV0MfBzq
Q6C8gMLIdILv8lQSSZwQ1noM/uZMDd6OEHPWOJbXDwpqCVspLxx0s1/pcDyzgQ3IU3c0FEMgOU0N
yV83MXPw2yP5qlm+RvIxY/9A89ude0QxRXfR3lUeREXig2qhZ+ksiLz2dGsvy6HOy7hvplwNuZgj
15oUF0oji9m9yaAyHrw7Dc+B/RlWe2txEZCZnyoG6FnphbQj2c/XeLR9dq6aDhIQuW+KQQP6qnW0
N7VYiaKb1TDkDQ5MDSxW6KVawh2Ggp3ROi2e/UU6685BSUTlJoxk2sJWRkQqKys/+TCSyIlsvu6R
U5X3TmItdPWUM05FSn6cqf6eFbVcYMc9CAFwuajoziin3SUfhxFdNQrXzFQIECnSiEY5nDqg7BdN
JyRAD1f0xsjYSZ+KDhKmjjs5FF02ChiQoxfdFVPtmbYSiFjVlOyyptqT7giYMwHQdls1X24air7F
UzVq/VQz/NgO5iPjPVyTIU2amj31P56dQrmO71xQhRAzRnXTPvn9CSIkbPJ1SVYlv9cW9b5ePGbB
x3Y2NK78MX60DjrAsv2PcYAvPxyEQybAZpjPd72nct3HRBx0VfzTZIFLmL9RXFq6yR6t0pnByd9C
Txy3x0ZAn9y8FaTkoGmX+WUVWDkxLw6zTXT3FVdO8c+6OWFiIcNkgy1BucyenmnFAG0jIDbaNvdT
Dfwe1fZhwzYPFhhPK1ejYopJlrCVCjPqzOcY9KYPxxqw7NvcgSCpMhuq/Dd89MzGIMOwt6cMQhEv
bo38yY0y2SIkh+Wau2G3YjeiGeJ685Ty+M8CjKQJHz0UOL95GYPNCOMlDW+YypfXKUBztwLm8pKL
iGvCVNhJ4h0sL6D2pjd3wIqel0A5683oWrynkDgl30rGGq2LvrrbeYGtJFpaqStM5ooA/2SEZVZx
4o+z+F6kssCpE7XtsiHWNDI9ej0OHRTZhJ9/9l5rbqDvqjiM6airOBej4QqZmpOghO5fU3HFMvub
ISU2BBqxPcTVcTDpO91IXIKN4JaxgoX1GRjOmENPqzYtvQlwQGMRJX7a7uaxiPGHj7F5nEiRW25Y
L30G5aXoEMit6AT8/rT5sTAnQCuEaPosfhpyTtp+vObggRpxqAmJNeMJnXfiGi52vbrGZwe33jKz
+RcfAI4D8FKMVccm+psLwaBH08lQ5rliHBA5kCskd3BstQ+bSWo8EW/SFBb8izOoTZNyMMYYJTuU
C7QSH2MLd/Unr0Q6Z+Yxm8f2ThbvXcq7quy0d0ZOx6bKb1beCIla89An/6j8OZ0WndXqRaKHh4Cp
y3Z+KryZBSFBTdBgFAU/553im55eaOQE5yzzHwUqtvg0bsCSSqqH6fsjoN9tLvHm4o8a1WMjsWQN
liaeNM1KWHRxmd/HsbjFYbOA9wdhGQ9sr7mZyEZ71Bc8W35LuLLAyZDiUx3lIzmW1F1NaLXDwMAY
OigFXIyq0ce2WODNljWbAt/uoUMzRsM+WdrrNKE58V3bj4uDzpRR5PMWXmo1txrJaq6REvIaoqqR
iNusB0/r3kaJQ9HEtbQ31kD1b1vUrAJx+NL8zrJC+ASLsu6AYRpwAf9WR/4NLYbZ9/SH3DkM2uWQ
2jA+w96nPxJKexS+ZdmR7321FKY5tD5YDDn3GSFRoXA0qjDjGox/kg7E0JhPPLPPb8Gs9whychPu
/0IVTxcE2kDXCSzn0Ei3njAJ99yLGtO/ZW/CaNfdri2rKjeQzwf2F4o/VuQ8pjshBpSRsLrPuSb+
bIv4QLqTpsBC82JdW/Jz/aeko1+EVR6XBvxNJHJH9VrxMIZ/zZj6rytiXtEAUFxMsOK6xdkHX45l
XRTOHIQnqY8Vc+y+LMuo89g9zaMGXSAQyQBc7JN0cpzvymCHRhGi4HVf8+Yi3qd6ES/pFpEmTqef
EEYYgxaJT1ayuKp83/an26Un4qMfAfc+6AgOtzRFFTFxmekVanPo0zlv+FOuID+YIh4PXF4TfkG1
pKbvpD9u/IGCfdgsmHbLUTCEswDGY1mkhtAou3xoRhNErDjdyeyhkcs5wGYtsN2WpPjTcGCGc6i2
SFY1JDEmxx97Oe1dvjom6Xslqpf08mRlgbxL7zm3sI6DMvkEXPHXSiRzjaKmE3WGZms4LyefU1jX
X/HszRwpZQ43N3xIw+hvGgaqybuzug5uybL50qiPt+nNk38lUNyXLKkMYfwQW1b1/FgxFexDpxPB
MfRG/UqSRRBihdF2yj+O/Cw7G7jY20ME2yID70ceifksdj9XN40t6sEvFtuW7WqWf5ehzZNhFc3r
ghzUfu+EG7OxAXH+uLDg33aKVVCV5mviFGaDtFN7jMTEjBa3M2ukxTmvcez11vBrsT3shW8lHDNC
RPxvGx58C3Am2Ln86skaTRmfcQfuDcMmS3XgKxNzz7sAMoCk3Wa46d6NAle4o+L1B9mFXexa7Fqz
5YekRn4BPLm4KSyJUZEuaRE5r+6hdwK2SZ1vUz6dNFarKF4SpjckIxDPUpE7cDaGjG1FikXgfkre
JlHfBP0AUOS828+OZrzmiV43YTBYW9qlleX2bhxPHzRd60Y+3kL8DpzYmBp9ngG3djB7q1UCVt6Z
VJHQE3jcif1dVaL8KpQQPTxS8epVBx1G4sb96+/8g10zq3UqgnqNCFgde+i578tkovz3VbioZWj3
LtkufvZ3tHU/TbThhk2ofy6ce1Mg7Jt6NHA5FLE6PI7nfaoAV2/Mz+kmEUvZFm8NdAUt64eQNJ1b
wPyoBUi+vUbXm+SEfxN/ms6y8wgE5CjRxHOlvnFJYINelfqi6l+3G6tujpKGsBfewRZo+sp2a28K
V40LalPWqHNiF/cUesp2TAthUlWQvDjC6IvRcBeomnfOmjCRYseXXANb8Ld7bvhBOwMDglsQc2ya
5B+QJVV8wogduBmQDaYxaIFzXVEMc1fZdEBBpGjRE9TundEHfKW3BBL60D3+Py4KGxZw9jZNs8jG
qILObemhqmf2kg8zKvj9ikvjMcmjj7H+YkbrhYXmlPhh8VsKzX1ILfXHgOI1hNRbi/NRUffpKimW
LSPXPrwJ6bGPo5Al2xCRvPcXiCD9nlH4DkOVaF3g579R1bEb5Bji8ZKhd+8qugHdDyWlonaez9WA
0NJyrQQHBvj7/W9VNn4hID/2g9cLg49aJiettaqVJU7LHSmU6HtaH65Gy51Z6dfYfPa/qZYABEoW
mEhhVlPnlCmAghpF/T8O7R2gb7+R6pGvVVKKR6VVAtceOkh6Jl9UomY3LIerAcq7d2uzyyiiwQrD
/caKvdQhAPW6mtZd15dLl6BBmKUhavOO6nsOtHV+e90ZyspRvxQhhFVdQdjGQNlBg1gzizdUBylF
cIUeuQSx+sxelMamnC22esfnpspAHiM1cP0D0hejxc7R9Cni4ROHF+MsVb1buS/MxMZoQ4xxouuR
Qt4EHpxbp+bHnehC9NIeFcC0ksAQTvfxoahKWiJhwraKG/H0n+gTR784yqTS7hwjuQQbDysMpN1Q
SFoZvbsOlnYte87iIkWMV9pRasGEkNObgwNx4mxFv4CHi/RJyu7nXjmsL0jb6KObek4MBc6TwR3J
EgbnotNe2QbmZQotfEt7RANWY1kF246gSMQDjDw33hg0KvT+JEIK9R0O+WymCvD8FBLPoLOfy2bK
5JxBEYm5tPAFnEehqg+n3/2lsQFYth7iguJE1PeYspQ4RDhr17Tb1abs6dulCmXezt5oYbBZERvK
n1Pt1g7X9qJkVLg4I3ygMbg392ZICBe5R7AANUFnsYsjrdu6VRKczVt5KhmV9IM80z+HpEeFYE/R
M+gXrEJI6JSVcUvxSHRgzKMq5wcVkXL6PYP53n9tfYJu7pMf9vY1FSmgYoi8MYEmasMLcmTGQnl/
9EVk2noXUWFen/OxBzydGxle5y/6w9ZvFfCKTwpy8ZkuQj+5splzeCsfbix/TP6kYDGiuDX0sP2/
PnUEFC7I8jrlJ3dAAVuNFPm805ZJNjdAeEbBcmU92xqTy6wyRXM8UHKVM+Bol8z2MGBIpUfkPSR6
myNDsk6GbOPfmXAkFXTbqhzidxlVE/2QefUz2QudIVWVA4GgbkwtZ6wlU+6stNVwivfzg2ygJYHM
8MiBdKrfwm0GCa4UY69tnfMNt9gVFY+6lTkSFRN89MOj8DQpMUPFc09A5Xhy1+QpeWUH58zfblWQ
D9p/yRBwk6E/qoix2qkeP+Huv+PaQOu0KpJia7+PYA1BXUl/P8Ex4ABpIO/9itypY5HRu9jm//fP
oHJ753m/lW4u1fYJAVikVn8pJl153mGhARPtzGUBQY56UCIAbrrg/ZtXZQyTATR+yp+SwkaISA/n
5YEtmYu0rAqE3WqzcB9oTzT9ABde69wQCs3gI8ey/1ejjhNTbTFDZ6w3l2vbKuTy/LPhvMm1OmeX
VSwzV8KQGhL4KVVWJSmXWXIle0D/9WI7FfDFzlx18YETIWcYan1YIIK0JUTscq1mfnB4URMBXoxm
8clIwEewRAqWfX3a+Cv0+Sof04UkOJzahc/qr4d1w/LHiI98BY3p4CrKhnv3gBy4/6ee0t0ey17M
p3kYWXpEXzGVnoQAIvJy8qrcRuTajNnVl+/CJMOl7kwoUGDob+pAu1vC9aJJmHSGX1m181cCroAi
1CDJjITYa4NS5mOMkCVG0rm5cQcT1Dh0BQuw/ZvpEuxQMh6tAeDS5mv0rfvZ8BiHJOWkmt7sWFds
M7NahmciZxX7wtlj3bOpsHzwNFQ+KVhrgrVkfDTNSLOJHwkJIYYGGlVfJA9uA6W2q3l1WBiyXdKo
HXCYB2T6fpi0qaaTV5mgW8b4eJM94Tst6BfY/vwupYgfoQbmEHcKE2SZKK/6MzlDondunt9Tzzwx
qP7ZTdk3fd9ftJmydyfUCyFxgjTGWio9qqtyCwYyhKq3dgWh2KbkBgsbiL/tjwnphMi0F+X/PORr
OEAhsJkZHonRDa5Q3jyk+d2l5BMLmGHMkj7rGMgiusTeZpsA8FvCOr1q3cNhI8hBhpo4unnbRFij
3VbQFzjNG2p9l6XEQA1fvayq00zQMSMvgbwsAARzpkRGobvKd1fNmIli+96nXfKw3HhKg53mOpIR
Dr4ZaDTYwzchS9UCFOV2I5W05JgmlNikYJ2Wg8ONjSddRJR/5jTwjkmrJPt1UkgEJdCHFxebvnM4
r/lc6+Syvn44Fe5lM7bxfZmPzCtjfBUco/unYQtd3Ppf6f/z/nPrqnDzliuhS4ed0K4+1MN1WL3D
dDjXNGx1jzPzPLtRZCtvXaC1DeVNM9Nfum+aRUOjgaL6XXXlw5d1m3EphLV3aSlXAwS+wFMxI50c
JTpuf86iGYJScca7/XfdCFotvVCpV0CNvvLZA5e6RJ92F4JZynrdkuuQxfQqy6ErQ9/8CFXak84i
VRZy0apySbmt4xp89B/pE+Q08EcY9R6um1yiUZUNLloIdROSky2u50yjAHJfMOqXMQeF0LNG103Z
XfOPcM1WAOCFg5GMypqvIcZa11TP+Fnt1/iMJB6mPyF71sjrOIgVSAIE4S5xR2/iwvOMpK7r/VAA
tixiYuAJ6+fAoqIAAWS2PQBkgoEWUIyUqQOTHwiDGKWl/WTSrp+8IwYJ3jL4LPV0DEBVgm530Smd
URjMJQgDKuNc21PzZ66d1YwyngRqa6kw/9sJuT9RYogEw4HnO060EZ8p2itpvI4tNqobbNKc4Knt
JNioaBdNYdbgEXZwys7ClIlMbkENJNOt8ZUMFu0W1Pjbt2AN0MoM0q6uSwX77dOgo8n3bGr/ywYa
v56VawMPQzSChLPtCPriAvM7bfKYbxx3531F7K61WiU5u/buhxnh28l9pVrwz0BUExJZ04jgxfph
hDX7e1a0q+QkgjnSYAM+Bs/b0pxfr6wY53pEcI4qeNvcRssunyuDgHY5DtdDeyOzAAG/frqV5sAP
qao8OroY2A1nC7OgtOo8O924Go4nJ433qWti7mn+h/68H9ZxHInRiyD7kwzY8+Ac4/XL7+FyweQi
cITASr0H8DS8w34qHFL6yVB5WXGchdNGAfv/ISH5jNhA2AADvzOz7MK7FTWmjRjZRjf4yX55itxI
kMiiAMvjJ6uza6HaVetUUmkzW8Ns3wpKXCFJ18sOmjVfX/FMpTh8vDwq40eVWf5dLCuHHjMWae2p
u8xNYlUYn9cs7f7WLM22WTf9ViZXzD7Vu4TEsirN9aA+SddpDkPOCjXewcAG0yLzSkiuq6Y3DatB
lW/CMmtFGiH3qB59buFNqlfnI28Ea2aHcJGZXo5BZZSncNsHc73/7ij++CSL3EBzihklrPAKcFdz
jJESCCEK5ZwK4Nbm2fJlAaf09dbOFFJyvN2DV33qmnnabH213EqD5t1Mwrlbwvfcp3kTnwTD0Pkp
RHKrc3BLgIyL6M1GjiDZHNNpcXhnQJo17MXeMBTHobOcPd/a/wIekApo/PM5jQzdrK+xx8vPl5Z9
GMIvcTQJi0chZ/5LGAzxBC++Q0sJgc71Jvpen3+HvcrDCd0m8It/sNlGjRruwP2A0ZNZOrRgfRd1
KWWVhb8h8wr4JHzvvulRnb7WBxNYVKYNMoSp41IQ/dSCjHGgPVxBkDsX1TdbEuANOfB7/uoSNx5x
YbffTDCO+WP6gzrXWj3Pb2IKM+AKzcx1nNRHYIVJAllObnsz1cISD9C90R/BMsAfKvMjPw5RPEDK
h33zjd3tK5TnAVxMFjNDa8o9L+fl49hgwmoV6p5YKSefdBajHDlRpQrym+uUbZxRIpDFhsrXPXqN
jVeQdnNo07KjHCGhRz60lNOdQ8t2Sch0S3QEORFFrkyePi64PfqpA2X8G9Qk0rcZ829ypI14BQ0T
X2akgn3U8a8wotzvkCfrYJBLDvnPT2P0oRswJusigKJWmftZfUo0XjP59IPVp4+bizEXRddje/DZ
n6J2dn2jQHHnjTwn0A5lLPlTZvIDQd7VIwAu1iH2bHfTH/D3cjH0OUUOOhU3ztjtJzG6tAutLWCm
Zx0YoPpxIdHTUVayTkuQjQambaJ13Mvakw5n1vUauSeGM+gcac4hRSjbnyoDIith/90JR3ZXRNGz
NbSZRF9x3RMN6TdbfU+OjmKPBnRgE+keOTucyK37JFkdNGp6NbXSoyC8XCaOPZiUlQft5jSLlQZi
VAt5756WHn/iWTgqa/ktfw8F0R+IWB+HJPLoXXFIEatED26dX+Yo2e+o1TxB/bZ4SpO+62k+spP+
ZIYgtzCVH4sRrCHuVqTvJd2r1MMIfWLqsDJB7HeWwDcTXAxwckRil+YNeaxkory8X89IkPT/iBxr
odfokZMHshe9Mi+HTrwq6L1aTzmZZ7CWewKOvdji/YGwCqMnm5leEhltOhsKgwBQt6EPQbDvmBY/
oYOvsHa88Y7bg09LVLjTh8l/BI97IfQ2AuhKKMpMQF2F0fjMJB4JxGsb/d7rh32zlRRW78B3mpxj
BcUWi27rfT9z/mLOp3UFtHxKXCv896yn1In1ZoIWoFr2rKZ+0d4gWv8VBGhUa77vvFcWSVurq/EM
NvAJU/ZVNmkX16xDm/Glyr8GgF80mI5mJAK3XCtr8ljj9rAilC3GuSlSHraXS9GGhwxI1k/eet3G
4wj4TnNvviQ3Tpj15DrJnfmiJ4CSAvJIHPK6HJvvXOeTkqEzYtYa3xtkNxVOxRk+GU3PeYnN9KSg
EfmodcPCrFEkpD5VfsMmn9QwgmwN1rv+wT+aE0tRGLiyZY5TOZGj+uABPuFRukWXTYxY0fAScGQ4
FpxYzltEBLdA2KbTPhw4o3+6HafmmnZwWC+ZR3BvuCWKBoMjFPiRv02uXoJCKz1fP9bYo+Dk4s66
Wmi6GPRwYHy9KQXppx8UPnxkNOu94/dhWIjhnaYF5YXF0YA954hRHhboUnlXwRrrGzkeOFWwVYWQ
/9SSVa9WhfhEXCNd5c7bvDYpRhXvONZLSUjDuoWqteobl/yxawkh/6biQ6AznFXPyUr3ZmZRW3+X
9ldj5NoHWiOb0JIaRuV4EYmDmkD+Zp29dPxsVaWPX8N23qaUcpJ4hHYy/7ngTlzp5huy6tt+lAvt
9iqePeAQfNu9vUgEgJ2LoLYswbIkfBAALQqHttINPcTQ0RCTHfCW684ZnC8G7FK/bK8SbAScInqG
srDn9NtP7jCU2cXnLXEFp1a2LsqqIdgZh6QkrXKDmk3/xmb5G66TsX/Db42SGEJyC2FK3EMc4kvh
XUipPXIGzaLjaqulBPTHf//WGjWmEHpBhM+v1kOJ8WQL8VelgeVIqRnbyXS9I85kqjNl5R53V2Ql
UTABidW27O8Wc6G9xWhCSqqAk32kY8HJhkNgRflzrDwVi/cOAVCIAtNnVlFv9iqfxR1ekaMbMQqr
dyZL/OYoW3FGOspbf4agGQyWU29B0BzOjdV6heSb7EETkanZSjP7bsJoiQi5/JHpon731XfQivJU
vhbx+fhmpmZW8Jrh5RBq/bO1hI3BQm3b8YkaZVV7MQ3lGfKSE9P3Hh14tF++iCcwIHfY5bUEoe/6
GAHvZYqQiJOSUViEBfBKOIBscp8JHFNdw3ywTMzSILVrUcaRTAenwn5rgeLYzG7Tjr87qqT+ROOo
Y+cVZfOjb4Y2/Tc0xWw5qWpU9s2mS0TjBikb4pPply3AIBqctAS8q3+9muDze9l21JzXRsiXzZSy
UVuzsYRnL+vzxL0XfF4GDXMJiAfDyJM4m9frYbc0+VIT3eXLogz4Fjgr5VP3hpEHmkyWmnrBi+iF
em/ewNRp7j1E41CuZ6EDbViBm8v8epOCt/8iFvFZvOpfo5//npUQRsfV/OnKOTJKHSE3H9JGSQdb
djfClIC4pYp/Q01VLbC/l30kDKAy6KIpSOiSSOiZYgU44t0Qm5vjZzEQSIJ/2TjGp0C1634YFjlI
GdR8u2OXcWxgMV+hs1qYTdX0t1q5LoYFoOtYs0aj1lWdKxfG03b2GoUXXfQ8dRRldyyZiNIFI1jt
zjd5d/Cf9DVvIj2co4cIQj/7mKySx7IiI/w40Wg1/RCYrU81fzYq6eQS2EyHRO2zLDfbQGNiKg7V
EH9k2rJm15RZ/xeq/huKLwCOwFQE4G5YswEDgUbmzX76NLn/zEBw3XwTqB7IJnjgN7nVoS9ByeI3
+2dHi7Z32rI1KyxjbPbozGlrKg5zpCFS8OzZg+W8O+yDZGGCe/wqDC+uEtwRBj+Eyn3aV7Gm4w2p
Hb4UlaNAaF6a5nKk5YdcXrHQVPSpXWVamwHzOp1FsH8f0cLqq6Vzag2cza8rwsI4MPV6DChyhvEi
ywtp6ETwXpygPGYzc3ZKpOAg5PvbBg9A5nzuW6xXR3JOyCXsDki0d4m6e+4Uq4xQwvptID0yUw/l
nGeS6jjNModSNYbBJy8AUQYPzMvVfqrVxMvShx5E145g534JrhnoMm+X7BbkR2UWjja6ksCxbbhr
ZAvEgV1NvOnzMFid8o3PO2zQ2yqH/jdBRChr2NRWKE52C9KWpAKIZPZH9Wn7nq58Cv5uu+dNWazc
70MTuzJGaKIVcwUjcS6ZIYkU2w1CilSsqRdvp1oQQ6pBsUEnyB1lHUuulOgSyT7PodxGP9CPVvIL
v/zdpe6XGvJWekYmhNVnNWvP4iSYaR43bzGojUna+8M00WgvBvbmfVV28nkAQaHPhUyV9RrrDPuy
FkTutk4zkkvYlzrPguCm6tlohiO11kd3Tg+WWCQ9SiSjRPS77CcM+Db+d+LbKbwEaeWkGGgxo7zh
Lu91gD0io3in/Gn0pFYddffd/Kfg9bxn6uy95TF4V0t8YONqzFcJ+IoTkvhV4xadbgdxSPBdwymr
Qyw+X3Xqdg7Ouke9CKqVJ3XJlDojnphcgb9DQbfsgb/t+kvAtBLUwd8PkkbWTR2kopFLKMRoEvQO
02qYrk6fZA0zpZYzdh6PcreRUohF1yYI2QC2jISBdyJEtyHwZk1xgCyPiI7VcHFKO07r/8Olm5pt
PZjvdUp6g3VseKcdkJLPy30ZwQeOowjh4qLu+9i/zP78A/0sOw+mGJlF2YGvsY2t0ejfMjFkoGV3
ZiXTYn3FkME7unR4T5lC16a18zD5WO4JP869meUHO7ChIDsonH+fdAeqmXF5lQVEgZaIXK8vR31I
1mkgnBPyVnHPq+eQ3ScnaIupUpPdtgGl+HTE/6vHkVD96dAqm68s2iJI2XHwt2jPwOkWMbSrCLSA
GEAkjZbCz6JyNCqjeTnBKcUK88K4DJW+om0+vPbpS3MuwtB3/YwvYZCF8Dx2qIZBWrFr++3sNEbI
oSac+oDVrgb1FxRq8PvoHd4ncGa9Wp+xrtPk7BuRJqMmbghp96n61oln5tYnjG1Gnqj7dfPYElNu
bXTeUrz1AwfaTck+hpbH7GLhfXwxmhUmnvoo4tGul/asieDeQcsrhGhEBgi+yfnsCDToRvKWZt3f
xBxs7UiVD4cStqRrAw1LTclQUavQ9coKRiXM9MJhy6DSBM1L7D0CIboFFnovbQKT9JbQTGPPIz/U
yZW8ah9pVhwxveqMqal23zv2Bedf3manoXH0oMTRI8eJTEhCFuZbmwExhC76U3yzH9KzUwHjkKNn
3gkm1RBKZci3Xal0eqPrZLIl98fgaZmrP6ejcEe9ggF+Qc0IW5lHf78Zm1SibV7aE0cjU0i4aLkw
40WVsqQUH9LWc44sOVp5G7dvPdJdTYt57RboY2MSNLKh/sKmM4mRrdTbfxGqWtzQRvd3Y5btLbw9
r0UEPyXlUT/gyfa13nyFdURCXbG7bjoLYYdznwMDA1Y6WZbHBZn72Ls9nS9riI3lm++EQnnv+DYv
UCiw184IbZCmBfdwSf7FCRsquH/00qTuPKivhHb4Jz931WOgvLKEvI2LPpOyXgPxMOD2pA1FoqWC
R9rly9w9MkRrikexWizXCeGPXDSrb0ujPlvw/HWSXcFNFNs2ZGgQ4lR4ek168LOx38h/aHYkzS2o
unvikxDUhSDYMu47IFzNFEtkq8kiQj1jyXo9LVedBb3zU+uxicS1EioXLDd3fQd9lgtnwJFibZpk
hltXxsYX4k4xvjOOoFkM98mkxdSFw1gVKJ9a1zdstC+DB+2dotlT/K1Et0+T0Tc4YFBV6bmVi2Po
2U5WfWdBb9k4pLkAsL6gzK15MRouUtPLu58KPG0aBEsk5E+jZELU5R/bWsA8yE8zY+PWUyhO2Ze9
Jqh+Sw03yQJ/+zvzmKueXsa6Y+H7PfrOLT6l3nb/ngNSzHmQXFxFNNiGb2RdR3yg8l0JuknQUIGq
StcmuuaR0II3PxfyO43OhOQrhM8qNm9xjQ0BUtVLyjivxsVotuheM2Z+H1D4TCZm19CnvZUD1Nc5
hLAQ849v50nI56/kxmVv4/JR4eDgZRBLWyxW0SLx/HBN7Em7mfECPZSSm6Vbv0mjJ+MS8znejnCk
qeFujMnr0FnOS11zpHEJXn2fapaqfSBNVppdql2HYhKCKpLkMpFAYVrZeArIt8zzqyyWeAYAn3Re
I1IL/ZGLsA2pa7jb7WJ+fYeMLNys4wTp1NwknJxq3EtXwL/ReY6sQ1tjm2kaBJ6NXPyElVYVKUzA
bRWwtQr97FQDXIu7mSzHDS9CU7N25TG/7K3CDsP2UbDxHBDGlnxwQ4bdAu1PPd2mouSqTOfUCD1w
/wLzHdzc3R45TVELF2hDKgr+gHH13NQ4vp15HllGAhrCK/3WSkh4k4GgB/HwXigPrAwEkwo1CVU5
yQj1yNXw1r7N0f6V3zbfjYTySPOxlGQ5KdXbdje2wD3OrqBdXIqHJNQsfhMbpGAmfSpbV9bzr7Qc
EWtIUjjxNYhMBlx5lHMvzuW3DZbm+XvBS/4gqsA67PKEN20xi18xKh7aUBOSX4j5Sy8akpKb2ojN
0l6Oc/spS9rpY4XM4m5dX1HWzz+SOVjpR7ZbaNx5jIN5FJKhoHEFO+QLEmp7C8S0pp6ilpIFjktt
LhkURxxjV13es+uhDT/84N/yvLuz/MtLuFINWz57z6dsovGmgS4qTvJ58CL9ePYlvXY9GnA54BcG
1YOU1H06kKO6Z2Ix+Pl3EBVal0B8I6FFFL48DvmH1wpzzIs8VqhC65RLj1VkY5QZbFstVBgt2IZj
adcHA+NuVRxh+O+N86cSINtRy7snVLi2T+FQhc7yzj4qBg5Snxe9SylPIZu9EHDdiF8/jRKrYU6u
1Bnrg698T4RX80+SZWqHrwSyUCeQoUimeKHbVUDydr6EAaODl+egdFL2jITPGNf9fR9FhCN0zO/Q
uYJAkQOo6SpZVRaawKBvgCehP3YJYmt2Pev+c00EvWJY1Vm9dT6HMVl2Cj0gE0EKMKTDu0I6s+3w
yMNp9xX5Itj/IXKqzOYhPkOfusjwhPjLR92TJ39Id1O++ZzvrDgtqatXeZGgWeNlZ/EeeoYSwgUr
LijRylvAxJUPKPBKcra6qjgsWBYgKCj0uYqFHUOyYJ6PxJqRkwAEhPlLfthASyWO0RnpKjpxEbs7
8g22rJBLLKeqxmrGx3j/ucXeImLElWMFfjGdczGvtusL9w3iBz2RNrVzEHweIrFybz2tKbYTOm8Q
o2celNp+GM8CIoTwayZWh8PSTIrGZZ6fLtmm+sOkWVR0jwXiQZYjlAL0O/oXQ2mQAGOls8pxJmS+
QdlywXK7bMLMupm9gC5lSwiSA4coJy2D3qiiWHX84w//Xk1Ln8O2m++6mCqkmfwcPHdRMSzaTXqc
tlh5UAxyvsjaUBv3T8b5M6vC01O+bhXLepNZKNoXsI60iYeAI/hcnBmw7Xwv7jt+V2sryTrOlW5+
POR7rnhiDlZOU6+nEkaAOlERg+Sz7CjdFkgGU1eNpsrWMXIsPhiH3Jw4dUOV6vJh3e2lP00w8ib2
jVXDfmOEx+TE2cqUOvRfYmKb60UPM2wFWcOW3bALINMD3FGW21FVl0hmBdOej1M0FGzOmjShAyJa
LfFeb34fQXg63iHj1ACY/r/1QjT4CJDlzKCpv/ab3YzNZlj1oVLPJZNQBLqbFX9Lm2ZsSaB29oy2
kSk0N0gPfdZDTs1Wm+eLJoHPG8NbEZxphCCXL+p+cMb/vd3JceH3UrvCaZkdct76fWgr74voByzX
afMpYT4fK47r/Si6KM9uLdkTBc6pmeAhEcX1vCE/yXoJs4dIvndPSjMerolPdrYGlwoYusl7rAEi
9Q0EAm2DqYs1ccWQWAj9fB5bCRKZ5oSpnBruoPxVdyG5GRLWOqEL28bDkmGPIOCU4c5+QOxA1rgf
hWcsxYiGwp28n5KzkCgWte7dv+OmCpU1G0oqgFkYLAPiBlBoYoLXnE6ug9Wv5dHwTrOKqdeHmXUt
S0LR64ynLX6PFdJysjePU/++iAykMY435EQqTeSDXAgw3LZw9uITACn4j4Ni+G6LnXnH1GRyBeEh
7064yELvwpUlWl1xYbq81uc881QhoC3q7LrcJj+o911iv97bmoQmfy7RhMUC1z2dFm7YL3x+Wqr1
fOBNA37l2fIxMVxiJFo9ORZ9vMHWSpcgtC6ohBgMEmxyCU1/BPcfkLROutAgCbNh6JVkgy3YNAMU
zzMSsNtw+FN3FyxEv87x3KUwS0ItReCvKNtUc5ucj/TgO4uDHpOyY7lXBA3/pEoug9yEhKXvqs8T
6DLchqVngxi93QUeQA05umGYSWsTf68UCQgrQCl0Y9/zzvSvPJN8wFHBYRzf7Ia4ySUZ6rx6bk01
B/lheDuB7uv8yEKTUxBI2PZ/DogOqVoBNzZU5rVbi2oHpZPKjUOrbho8unUIPN3uvsv6g0GPDe1Y
oDxJOCW2Gq3mR1CZbTRXJRMoLe9IY2ZHe1xLgUDgeh1O8A08f/+qu30e3WKClp84SfQHmaNTKy9S
juQeVAtHMY+OggaGYNkXdBKT5tHN2cOtZQf82E+kPSCsYCndz09T6Oi4VPW3qRUvbDZOx3xMXeqN
wsDKsxUGmIfLd2JfwVm3WXUltGipOXmqNdDMQAXCmZafO/0lOPBOXBLeReThmA5yA9li6RSYE+vx
INbCRfGAPqbm0NDM3zgpPuSKYxERkFDM94kDDtvWitDtZB1eTt8jGDIQrrxll3imXwFhZe7iycjD
16D9gmI+V9pXUPI/MYdC6WpGckCCA+oem+ppFnDYJP/vwNujZ4mrKqM4FyJPjsxS3LttP+mak0eQ
NR8n+bY+NQhXuAYleJm6LHR14Rvz0j/gdqSsStak/FyW9JZ6URZzQA7gPILXn7YYY6mJ7t/xK8Fu
8ZwbeHTBATOqswXu9Ss2Z8jpPXvbYM1QhT/GX+uofTpkkPNC74HiEUCQ5Fg9ylIyFTiRWk1jtved
VVNvKvn7ZLF6GUHTHjNoQKF8j1y9d+5O2aW8ke0e/CXi1n/7ssuOvn5vSxxkWao0U/XFODYaYKD7
5l0AtLKw/js+hryuopFIfJf66rXC+ONOZX5SKQE/ea/lBF3Jt4UOywVv/gbSoU2Sfh+uKT9+lF1T
HcDBM1/kF/4FMA8sXEvzM7E1+IcRFQG1KlD+WAr6LWJja0K0fBB1ZMaFhl6oiIDLz35jCjUTnj/5
LPGxrKyeVL5NTVBzArnPyecw5Kub8oGdHF5oKXYVQaEpa8MB3KLArdO3NaFVmp2JwtyzLJnvMVdY
p4cHRSOf7JDhDMBtLYm8X8PIZgFEm5d2YgxhLhkFx7yQuSi7dPVsVNPQI2LMNOiSdKbNhsJr3rxX
2XT++YTVa0mzXbghSbFxx7XDVshiIzWhgZ3ISv7DlR/ymgS5igq4tdRL15AoVt/T0mIWnip4KCEY
nSoWnLNYtW59mwbmY+cLcjwAVqZpgTQ06F1Mg7sJCPYwlthMxoTLiPfn/dYfpF5m1OeUj1crywVJ
XAKW0RfhIhHuXMLePFhvcLOTBoyjX82/waH7AAMKm7AqabIUrWSC+Bpa3Em1QsvfOYh5R4LKdVDS
5m/IAUZbT1yG2BWnjn/YahInuSf1Bt2vQyDH+Go+H4n7MFuPmErBCXXVTew9etIYmdEpYtdp9WA8
hrnLbJ9+o0Xa758NU/8blm3zLuCE6WVPhNCfcVJamtNgvvJg6vZuvm43Up1qjHvyE1CFFHYG9NDF
LEY9n/EuAmpJYrtGyDS3CXKMY7rmgWKOvUBXykPzu9NH/OZBJyaPP10ubgQooBFmfaGy4kEPjuPM
FTNqw7ku7AdM+Dup8r7Mkt8W7n292dj6cOH9WIGQ18Bi1VPioVy+Qw7YyTG8cjKugCBX6kwJYvt8
OP1Fnj2m/vBQUKBi9Zr1Yi2pZztNQ2qVBzLoQdloCGqt1KzxgPp9/bmOtuF9xAmfDGlPYxkxtgLp
S0NSQtpMwpieIgwCizDz6/Pl3LZhBn5dMhK9zjfSDPla9akXtcH6Xgv2hApawvP6lOc1h8Z3NOY7
8kkuH3xwmGypRGJSZbwXl47B88/xVSdkqLCKKsmY7YqMEAyQWKHQ7nuJDuV9Xq37Jds1FsmgrYoI
VLItTo1f8ucgXXTJdk6B6UJ2AyCRjZpILrTTFv9pieyuY33VxUh+mO1sjwjYh8l/vqWPhY+Bep2K
jNi01iDwnEkZmL0yHTsjkn8qjOKAaqWhnddmFRUSh2/Fo5lliNd0RjbvpvcmBufZV9c81wdH0vIE
XGj/20uwsC2dgoG2ScLhUj4+JMtYmc1jizuk2rV2ZFfL0rv9J/uGpBoFPPPhuQhd+awMRceO4b4f
MI8khzsmxz+rRt1/2eAR4uzlIo39KdrjiRoR9ApRVy9oFdLwPs4JssGzvCCpnBZcRYl9nQeBEOft
CByxQnxddRfI12e25hQo8VQP5DHELLywouh3AevGAoCUqlyJmC/Oj4w6gaSU+MCqGlzdueiOSphq
lAqShhtkLS8rlryXrGKjJ7xv5HuTxtSAWxdVCL74Pm7/5PquwootOyyw2oWPq7ExaJvsssdXiOkZ
uA+qogsGYrbpa1IXhpVrk1m3aK8ipRf9iXlCwmMGRjjMhPFPWs5Z5uE7dkF8SJaqOsEblzknuy60
d4FQXJmhP3PKaAHnH7BrL+uzQ/Udg8tPv7hXOU3vcIJZrpfyAV1iJwNYOK0fZuPfeRZiQn33HgLw
a4MwZ+AqddK+B5CxqR30BxnrCRArgsQ0ls+wAbZ4d9E1YgVf2YHsCnHDxfw0BKcgKAWJRS70qzv1
8BOQ6HkIPQfx5wJ8fnIR26WUFeYYxfK9v5mnv3rIVz6kcQhzxDdGxUwFFH/qHhyQ5VLWxAcvEV14
lrZIuk2sH6oB4ALH5MjaeMXwzx3y3Jh2gW8CiyYgrwPur0I3fVpu9LAX71O30wMhGOOAj6F4yY3Z
yNl84TwfpPABrJSgbT1WM3xmDNUgfSj0brFzxQ0zSFFkb8cLc7+r7Gr1oCzHQUQrO54y525cGP5q
S0V67m0CA/8Wkvpvo6CF8ql9ur+5Tljha1v9LIlWDdTTCepvvodkp1cdws7Dv7dcfaU/T+BRlK8O
r4R1yHi9KXwcKfGs31zYdflKvpkONOgicDrlHEOEKxf1UE8iDAcVxgWEUqb079GURMnYbAYG4wQM
d+U6Inn5u9GIHURWZqtIFeMikXhiohKPNoroCih1JAQwSDIAmEyLd71c2FcDbxYEEHLRvdutxF2H
0RYPMaReB/TWOKEse43dMeOTRiRsyGMqMSY8H8a4BcW/nPSgdakPAKVmVAzcYcftmSNEOdEnyE/2
DRdWH/ll7ILx2oxY27O9310h6V043LiMZh+Uy08DHoWC6PcWtA5Lg7CzKCVm3cdPlSrvAzm7UVxq
Vt44PyLNXflXNja1Q4BKwihoIzBgho2V5FngghVt/QXqWjaH9yFqglk7lwdGhxCDq0NjrwCFRtCx
Z6Z3NG38xQveiDBQDaeZCz2cuuaQ095jhFXHYqtaZny+BQ4E/eK5+ppYkHFkwAdLxcwXIJ0Qec7U
wfAWfLwUDD3fT2d/xNDuO1henj2sFzQvIdsBkpY+xaEgxwuRKq77G9JSCMjlawYg6xjo35q7+R1z
pfa0DXBaISKpmyOcgEwlvXNK1BaZBZBSHsgy45oqiewUPhzBIaYdFh5J1g0MbYQdNibLY6K02gkQ
7SbSN1zSxwkfZ68FykhMaO6fWsYxjc15y0eWY38a72HSj/SFe19jfw7Sg0/v17tE0sAqT5uI+LfT
xxXq7KhioYn/I6lIalqGLSbxFTw/Ll94CNt0u4mzAW1x0eOT2sHwQvkc26z20jz49teKeu5WlpkE
eOuDm3cO826wvPSlvgc0SpOXU4uKg7IM21YvZVdZyXMKSD+EQmUDG2Or5dreQPTasUmJCdAULXxa
Pj2peKiXKLgHH6kyNS9+/sGy1hzvb0X9paJhAbo/+iaXbM6wqo8RikUItCv/GX0BtkAV/+JLZuBG
mzxuJJwPRFR3oEimqhMIygU/gNm+iQPPCoRFUAa2TUKXDQuh3XYtcbhtPy9SrWn8tJ4dqoa1RJNk
HDOVmiLOOxgLttdGdh9vH+Y4yH2+1JNd3eXzSesjIHbfoRhrIM83uW3ghwX6OZJ+G+O66hid5gB+
bGo1kDPH1v5YMlJ88pJiBc/cEFTycton98HQyS7cogETJ/as9nuU2jKJ4XTeNL7maM9I8LSuZHxL
YVwNnolZPV6PkILh+lCrnR4wYjJvkdPbVB8j8ppneLvLX8t1Z4C/wX/YkLXpSnslRvZ9nbhA9FOJ
/QNhC1bP7EIDYScPNnKf0mOH5R/zBEoKJr2oyQ39jrC6zqghffMndnhhKP2u1bXEc0mOIrpHMXts
iz/s5ZXTcueMfUx/9QX3+wQ+kDqRiZwp3PjdGLqEN+juPGrWLwZ55E5c99rXxjc0+lR6c/UCTFvM
PW4FZrgZ1OzIlqmStOatQECpJVk4Ax8ebxbVV7nqU2eLUuodQIXIaNYMDZEtG9F2MxZZIkv5BSct
R26+zkdHgNoClTHE07/DoNJ6+rIFxH9CMq5fm4sBTFsKUev4MlVVhR49vaal2EA/kWFYLyh2sqRU
oBEJm12563rt8hrmdoBXyl6ZxoBI8GsjpvOPjzDIQMWASt2Rm3k481qCw8iFuo/pBrJ8+QVZG6gV
f05huI3BbL8SUP3nP+uQybbwKeXRoieRazsfYVOMSXfbfEwIbA3biGpAJk7Oz+69NNgQW7XESSdl
mWn3igh+c3hltXH+BwOXWgQwXSM7VjUTdIerCBBh36tz55sRgGhgKSL506yr0+8HWdubC3vCwIgG
6ruALeoDNPEkbF2zO8DYTPkdznhLH0QKH1IK+MwICoeY9/vkreTvZ5qPLYfOaaGDOgDREK9K9jcv
Zi0W5o2MYpQTiqJ0BPnzCWtDxiIZisuulk6aABq4zmcm7fubbE/J6YcaPtDMyi0eotiYFYB9bOrC
tvtRe5iuNaK3FA6BahyVZ0MJvQeihGknlYI6Xj3J/FnkZ1gRfiTI6F81McdvzsYyLsg77H4B1ocu
R+U6T9UK5l4MN2QCdFjUdwTmQGKd4BbIIGWH0eaWv6ssCVKXuRy28fFT5iyHEXMhxXMq8cCFFVTy
iemfiwLJ0zYmPkxuaoDciyNc+4wYfhfFMKWsjLfMrZV7lwMcA+adva/hzuWEgPRW7IH27cUVe93a
u8GjkTaOQVAlC2ab6Rp8uVP4uzdX1lqCAcxkcjZY0wBjZqN9cV5FcegJ5aBPolWBTlsrxhd3QoCT
Vv7T7oSq2hF3P0d3Q9pIUXq623C+g1B/lII1xDcYrSqXCJf4iHpcfIAmF6OsxeuLUrJZX+usQjTD
x6U38l0GnOzT1SfpF6B6OJNOZMOx36fbVpw/ZTFTrrquLs7NaS4fGOXgkY5Qi2T2p4QD6PB+iPJV
SaFasGTk+U5t9NfAWeE8tPsQh9wAafrKYhEgYk2GLYwZj41NX0g0qNhC5ht7QMiFiZaVtHSw2n3k
Xad3VVzPMWznTfGifdiea6SzlJoY5d1KZIyTR8ZCUhXUbkQxaKTKm8rPuV7ZpwblmkZI7USJuqh6
lAyc1bm9CAeR+A44vwgWYmQVyXPPTn2VRu9uIhLqUtJ9Lh1Mcb3F0h6YXI22q+7SMxgYK3uY/4x+
BGPPSbRnKxlhtTke+Ptio6OFFHbeA5T3VyXUZmdmN9WBP2zDkgJHJKJUoETcorYcS14l2Ne1FDsn
f5GYnXKUE3znY5lMEXfPBke4R7AUK2Ff6oEA00lvn5e01ASI/GOqQuxjkVpYtdpJzfqJKyMmc3BO
TVJz0Mi56d7v4Q/E6vVhfHL7W+W9va49Ocp9i6CAq82nscB2qAqGULA2GmmKQmtK8DftwjZRrxoo
YbCHxBnunbCqHMElVUJqMg46Ltyn8lkDQ8YROZYSNmqR73sioXaBX4IOpH/QNOtR2/6IGVdvx6V1
4G2v2DNmg4W/mBlxwGuZpgCaw46HpsdenchDNYO7KGYPgKI1pYXE1ZWvrr4YU8hTVz79tnFxVR43
7/tD2ZT5rEDOJ4wOWTlFmcx6zJ0LCY1XtHxcKsXY4GbrSGYAWJ6f/PLFuNhqulNXMAyFqV0pGvXT
odw1YLOJicdSs8Gw2wS7l1PrYcxHFnCYWPBPLW6oQ3F5duXXqQ/8y1PSosgzOs8tmwDLt+aUrzHz
/vrNDufvYEPiZfvjHEkrCA/ZRHn0ge2dbhJ1JZ5Hmm1KJF7NicAxXA6D0sbozlNZy4AntFXC1frq
CzdXCoFoT27j7imqoCbyO22Wb0/B2TtNMSU2Jv6ghABx2e+Z2D5efEf8BvtyzkPK5ZFBGuukumoJ
yYKDdgvlxNq6leBGd2BLxuck/0HGy0rLs1Scymv7hmNiI2OMdthgkGL9Y5dII9MNubew7uhLmams
p5rfQmOG1B6Y/3A4eqL2UyxmrO7x8NGMCeRoW96obq0eagC+KcDupEVgEGCOfbt6KYOgJSH1FIrE
KWLxLN9l6S4WwBYfocoADrOJT8W8evYtkjYF4EkNdMof9+Y6wKRjSIYsW90G+yzikRMJuiusixLM
xH9GOF3yGKcZWiXTMES13cFldpJtde6Ube93tzviJ55Iiafp3NPpU71g8nlEkvYRsdXQvYwHecFV
S0V+eLHDr2TJMSjmMRtS0ZoitH0lGKrQnVpmyFrMKMuUT39JYIN8B9HYj5UOPjUY8wEJ7O7IS8SV
xaMgxzc8jhPhyjpicuIgiHSNg9oi/0fXuDfH37JiCuSPJggo6QteckSdLjA+bnnep983srLPcIeS
uZP2xUP2Xo8NzCttadWWfEDacXp45GqsD0Gj9zRPmFJB44KSlzyHyc/zba81z9I8c/CNQd9NEVZm
7EXzZTGbEMmY0r51kuexY7x5FOLBQvd347hhNUSG2i4RjXgSZfS9MDOMkb5cHVIwtjiJx9gfVRJ9
o5xZcw/SDc+uqJ66ikUWkBcil4axp5iEn5lSFMR9IXZ0e6qQGmts4xxII0wgD1LfO2VU+gJC/Re5
XJmMXQXe3++0Jv9YeJJGKI3/GhVIcSID1pyx+xU02ikIcA2q/eYJoe2ivA1o7T4oHNj14vczW6cp
LG2JuQnS+PkqAZKPVneQanWRbHIbS/LrOU91/IkrdSpWWHFKNh57BB3QL/kLd9PA6/Bi0NFuRchg
vARoiPkKlNeF4PXEtWtuWOZ5LZkn6QsaDHD+3cf5Wgp8xnFsbHJZwY/qca8ibzFZIL2v6AnjLBaZ
VoPa8fQ7eLJWDMmJ1wAj+WNA2KcU5ecUBH50PNZppg7qPhNYKfj3Qz9gqn79Rob3rzzQ6QyxvbcN
AZ3Ti9q+u9koHS5LDY1AAPhDUb67EGD6rqSaHn+N0yWisMgWtHChJT8wSuPyOLg9+r7mY6vZW46J
bLW3/hj+LkH2P6co2APGPqFywNS0vVselsLO1uRSmDz6uiL9Dp4Aq3cvu4Pd6ELSakxu5vXZ8WNK
XCNe6mhP4sDSBzlHRrM2QCfZkl7y+G0kwyzJ7gQwbVi6ix7dM9sDXzVkx5YOD+7YvH3zHlCSXCcb
vOD3/tEVyejXsrmF1AXTBubLtPKzpnVvBVMKpxNU5qJ7Ag+37NkBb/kv6S2/dA6kJXWED5ST0j2m
J0XuMhrqhkZWQN9kFm97x/JOOT9TQeEV2FMGecZeWJ6+GZL109fB+2HUGsCQyTuFZsngMZOZQCwB
xsDYkoQ/q+YRBGgFh6wzfEvNlTFjT4VX9ylMb/pKqeSftaQNTsJLOmQYYLU89OHXntz7FeZNwyBw
x2lEJ+xIv1qOIjn1r1BUsC72dxeb0Iy+4NJ/Mz4iJGZNAQ14F5O26SZ7ENaUtegbCOqXdrKK69D3
7qqrS0uglpTAIe0OZt7grXPn/L8XSN/B00Cz5coqJ+4JsTAFOqvWWHOiUwLS6IYbdKmCnV2gJnNN
6ACuNz4I2niuq6ZoEKVC2xsveGNNbGFt2ggOjCt65IgNbwg/efCf7ZYXNOZI47rOmAlt3NeXtj2e
eSkkDkK+N678r/Ryg6Mg/SheZVRfqwAWvMd45I75fxgrYTPzp6ml/VmpeXZCZQT17HHx67/weWfL
ZI+LwJjSmZUiKvT7Iz1eaVVkwrEjIH1aDIMW8lABIHDNEB5jh0YmlxDJtwcMC854Lzo2nDQ0NsV9
maALCQMZraKRJtIBOHOjnrZGzY2SZ8Qsy0DGvaOyAhghad69Ctf9gQMjaVeE/Wo78ZxC3Ul/crb2
/O0dBxbukxTIRZNpUF7qRV6rJLJd+R+af4gGnSBWz6nMvQRURO+OqMJcCcXRwIHNBNxoeNuH0qK5
m/ABzS6DgdWbfgbgCI1GI16NO6rai68OG2noQXhaZA2+uGKHBtBlFDS4qx+MWl5kKQ9Dq+kKN6gi
3fwxrDWZx4Jq3Rsbqq/xPe2/PRCamYpao0JyXTbaWD2lx1e3tS2KJJk7TFzS/fejMJN9w3e7hmD5
3DklREVC0t8Yv3GZHrulSpyKe3pCtW1msT0uFRIv1WRY+9MOIKn82SmJBMOG/z9Z1FTQvqYCuuWK
fWGfa1octvMXuxBSQ50RFh74GVLLDe4NefdWyvX6iOUxieKN400IoLLV1r+9VoksokZxNGBI8/6J
0jKN/nnANA5mW2jJj6YyrlyAwlthj3BhLhuKSXdc8CHDTMvMAmd+FFml/4HxZuF/D9vs4uScCrA5
yKSNxglQaIzA+nQ34dmTXeMUR7K2S0auEeg6hi69vCFj1X4alDiN5JqrrXpNNke8z8TlaGtICaWW
htSK8S73vxi2HXkGijr9WxhsIgIiVwT3pRnG9di8wCo+5k45GDGDQmAvaeARYz4H/oY7YKGLUJWR
W0+CpWViAzQN3W/aLAlDw2Jdwsktrn34ifeZRa2S9kWmYmbYWFDya+LpWMjy+n+PIE2tw14GsaWr
5iM/syFOa36KVzPBjAWE/e5Xn1GH+t0Q9I5Fb74vQ3vck5jljKYya9mAH27U+4GLZjkuTsCj3jUN
fhGVAbaF+yivmUgdiqDJiD07hR3Ofj1o2F5QhNgs5zjLiii1bEKiY9hALnVjuEl5aqKqv4Hsu9yl
FXxo8cpl1kwxr8HRlGWGaLPGdVTpkIpBBsW66eJSfpNElKAqnWnmBDZzTBHtXHjiB+Iqg/1BVr9e
hA8vt1NSgnoD6e7Fxe74yHm4E4DLQ8jtkfYTnwqGkvjgi4shYmUGm+DfgnrewPKvdykFWqLCC8Vc
3EfnJv4qcg/bA7bkCl/N/qpAUYA8s1sakFElFfHk0wOLSU92IqhzvR2wq++tWY+4YudLU/kw0N9v
dPEG3wRjZoN5Tgz8lMFZaKtLKXn1hGSXx7aGZ84M8J25ie3xJ4GdtkbbiegBr0khQt5vFfCwHInU
y5XXye+UOxlDlkX/UQ6+vd2luszA3uK53oQ4TWTlTCGYcKrhMsuU+27oF4dK9QoA7FxZBClT/46k
BJ0ghc8PDCuVxIJgW5ATv8Bc//xQBjPDUsz7EhRVgSQpsTNwnE1DqLFT49i+nFQMp5SpLfUDe7DG
Inn8u6m9xoBtw5le77HHUkDxBWbZgh4wwjQSq8bCatXOpSb6Qnx6YXZj0U1Aa0RUIrxItR00HXsc
L3dhrUPtFl9HHapnt5wP9gmcWdMdhWw1QRaG2/CcpW0xcJRU3G9Di/cpHx7fGCjNKcIqfbxI4Hr0
1Adv+ZZNZGcyXxSEPAXtf2Wg7g/95dH4+6KAM4A7ZijppEr8Dn++hayxETtaosYCZ5Yj/9AKRHtA
w7oTaOqDKdCa2dhzI5iz7mtPbvEgdCw7ogSdlr4IXUshB+8UpHFDCfx8aWeryb7t9DVLtwlqD79g
VOdJ43dFvpGATlsnjW7kMUsH+4ThzQcLFKR0qzQhYT+kaVkjJr8nzE+LvSJgK7RcpZk2M8vf34Lq
UoQdyGm8ZccCkk1WHiwO/Z6uKgSWKIp1qwySZ032Qc2Ktyw0dGe5Ukl6tThuV2s6nvSHwbTi+v2r
fBFiYvEYgQ8HbePAce5sL6TKLivlSL4dFAvmr1VN0dHbt0iXeP0wuS6YEYJYI7WQrNXMbx7w+2FL
8u71KQ6g3R9oObDuNp99tzxCt0TCcJT5JFx8WKRK59Yw8OdtLxZN9Y4D2NsbWQ+pdxEG+81osiQe
iFSrnFx1l/IqXs3Us2JL4i/pMJKhY85pnIjbFBi1a6O3gtY5+lfVszaxTQFGyh1mqXIQh5UO4maG
u8IHRMQKH7l57BhWy6lBW53rji17Uux2yGLTLOLAEx0Mz8c/S21rAXT+XRHh+4Om9sGm32wF5ThX
i9v+bNhuCOnlEEmYx998Zeo7OFmBCV53++aFrO4ciAsk8tiC9Wvn652vI+4KMxelubyU+b2A1hfU
5P5RPXA+hQJP6r3bxXdFBscJbEyL8u3Ow56MT4lwDt78NwiMgj4F6HJIwYZov9ErdlWMetxHMrMy
kt0WDsUh6yloto3jmxWpHbsG+OUlMjKsVex03c13M7r7KRCwoXVRbvwFGmHjGv6+82+JzkDDFejC
I7HYjNRv3WgwfeyDiqj1KGGp6+GydfR57dOhCHrGr2wsyUtktSM5UpF2m4DsVny3D26WXQRXjXFl
1+cwR81a/lci7y1feYgn6OjnrHJ5BZdpj1ELYqFw6isxWIif7a4djIS8BDMPWAO+tdioV3EsnaE8
6rrmfKT4U0pAYDBYAToYpSEDE7X2AAVjeV+ZNpobgeg+3/7R3ltGyfPA/W4cc7h6B5WRjZ1FcPIW
ND4FGbFt5KJsGzHZj823jLZV7z9zyu2ium3VcbxRKk+vM+i7Y6N2aR5tnCvNgz2FAf/KjvRGWvko
KV9Wkj5EJVf+cJeQzcjDsOgGLtNtORksuRp9Tewsnt0DFBZigWzaltpH6CXoxRz7V44acb2mTq2X
KbxE6GIrnjoSdgn6qhTNVisod2KMi6wLqQIZ50dI5O0+AJhhcAXDOHyzFmJPbBvn3uC87wDD0Ygn
KKSngi3XaZuIQFMZYGHjISDbkXEI6vbwLAPFrIdCe+coxrIy2RIfqy8G3QsjZ5QO7S6mj3WA5Zb+
xvPTOukmOnEY0ouMgtFrYpnMA33+U/RJmARKvBBDqOqk4O4l0nQ+tIaBJlmves11ITTNm8jgG436
6t2goqVUF3v/Lus00tcrVxNep6FCHjOeZKV9n8JUYMkZBT+4CNg47yA+uk10s9CAW+JJu1fMzd9h
+9gjbJYwtw3oQRPT5ExYANyIfOE22LHUPFfNH7XxiuA8F8UXNiaJJp+X7wAB4PPEGXDJNN+kWKV8
vKbTTcbqy305O/EQ2yKVx+KZrjhpA6ITP3h8YNcUDMslMk5WiT/05ZUwmFSzBu4aM2gBYVjvHKKo
Lc+grshWIwz1oN38+gyj146D6Y7/S4eUNatu8Evhmn+igBkDPp3a25vupenlrZVb3L6oudreiFq8
8s1qhX2bfENhXw3+pDyddzbDwxkYN1PLDW92mUMLKYHjqdGkgc/Ni63xn5LV8z2sz2Jp4dqptShw
Xz6DqK4mPjkhpxuR7RwImUd2Zy5lsg8DLhsrr+fThorwSGL+uS/dp8Sj7pmV5yFpJCMSbjCE7jCW
dFnY9coPkaH5k2wbXTRfJYiD3wlpgAAGuSdD6CtQ2n3Rr6E/TZlSdbqfti8sv3c9YYhykHyUAqcB
K74ELKRTPfufTeYrmQx+/rhznnH3hBZCqKVTJE49r+4T1l8TCSrIbINfEfG2qy9q3rftFqw6Rl/N
xoD8jDJQfABIVV+3d3vKREoPpSQjI0qUy4ZD5gQgvKL3zFsQmk/qNSE3ru28npT3wvznZRvRqdDk
NnAI/frYkN91y2yI2JjUQJdwFWFJ0DjViDtNHMLZHwmdeGT+apfwr3qI30hijOaw7JV3QhzaWRbw
Hg+Z8Hc3s8Dyhx/x/T94px7fXrW+OvJrzrAl7Wb5G2nygWslgZe4QmU+a7ZREA6ZfhnMfbtBk/Uh
m1BJCOL+4w+JyWA7D17mnFkWde9hCWiTb3HT3exMTA1GenS30wStxp36POeR7XiWbi21ajafYx88
/NkOCNW/7PaTqJDI2aMN9yq/MJbZINfrBk3AId3a5g3NeQDroGxVNuFx4F4q0lP+Erxrjl1pC2K9
FFsLj4neHJcMkj6R8tTW4qFYGfKnefeX15tnKFB3bBuN5XPtLvvk8MQGVeYicNlHlJDWU7NVTiIl
srqZVdBOOsGSnAET6FrMeBPTqefAWYXPPD/Iq8wDJpeA8zJ1x1ERFqUiE304mk+tvUvOSsbAOS7d
O6DxGjit4xqHnwethjmt3FPRKZ8gPbfPHEQeCW/JfUczRbRB3ZzOoeLT38QyBLSScb57myELAAz9
hgYMTQOATqCQwIlnXIlGF4n/U6yNbIp0yyqhGLYnTjRLV4n3nYS+lFIR+WLaHMCV3bxF2263YhpN
RPqrHxB0awfcm8qJgyvxVaYJxnjAjuMXlUM5+wLyw0AxYgKZL4JMkIq5L+Qq8EBIqzkWriSFW++G
aD/961jqUvesaNzYaIOZ5ZWsLr5aFH+f3EPGSmt1vPXpEa/7agzsJCVDcYp/b11SoqXYhr/SV3+6
QgVUj1BKzHlJdOCexxg26cSpqSwGI5rEuFmLxgOHFRRwPqu3Ig5h9OqIZZkGIwSvL/+GM+G8hdIv
09CEpp0DjZONm+MyvOtLxb5buqKkKnu114wKRhEdFQvmOjlRE0BqALw3l9aizXPhUrX4t2xyj/i4
orxASgRYmVFZL4njsELNO0nf1snddHCVf0rpt34RkRRJqKv76xTjtluMK4mn8uqRGXpCaJRVJ1gx
9mwlO6WQ5X0mUZO2YxGVUlaTm8wTu/hxUiitPuaOzbzSBkoJv9/P//lSJ7GjmZYhkdcLoJGR5d4f
XRVJQcdsaVtLlkOh+CkvUWJqy1hUlf3TcIdBmCPRTQhPtB1u3FXOOnNVogfidNHM01oVo1Sd1geK
5EdW8QyUueP9mnjaBZ7oZykisRh19yB2kcGraBeOkYdcAnrLcd1hRmXqdZ8GcQnPbjy4sHxK8QcC
cLi7VuNlK+Q1hGvNp57tLOrYQNJcbm8cfRcLLv4XLu6s6uYb0rS7m5K5uyb+0dkcUhAIY7q2gxZr
iPKBvcs9C8xHSO6FV+2SqXovAITeu/sBz4SLEb+B5fLYqeSoW+EI9APO34qSo3B+kZ+EMTnbKwQK
9CsNZLJ3y7BcL4rk/keNJELYXR2chgv/biPxaEHtX5EQsSzkid78oqUN/RlBdCRtgD0hazxEkgZw
uvO5jvmSTDjrWtIpLmpULSHN8n8ggQBhVG78o3nuRqlVjRNg9I2D0u/qJ6yk4zvD5SfPGrCyHUiR
cqfqReDRfuGeiXfaRXu22H1Ik+qU3YMgUXtY8IIDSZMcOd/2NLAX68Ryo3/auAKvZeJEb7s4YXgn
QFblnYyzGGqzSDWUdyD5AR68PnaSE7rr/b6eEuO5W0J2erygAqu24GM/DeUCF6kfCEoCp7GJ1Lii
gYou0CqhHMkVkTi7FcZisxcLN/4ROQ69iasH5Nnu6nYiUmks7mfiD8z7oweySbTHQKf9SVEwFlZD
fuOUrFO4RC0uw9yCe+NPqzPyRBSM2LQBfR5GTRqMB+4xXBVCkxbHSwMowD5YSl3q+ICwrmCFT7Z5
EViz3+j8sZXkeX9ssjOJSrdz2QkD4Eo1svIzf9J6R4z5Asu0XI6HzGpN+bfyviyvySzalOIzJ+ga
amyYGUbQtme/FjiaXFfcmEec9zTR1PGyRX4AuTMNAMy6livoQ9V8KN3cRHVg6DdKvZyQBV10qiSa
OzGT/zHxgpGucoGkVPVza++a5sf9mFpISRQ8cQgpfZhfUlyN/OzzAOA27j+FF8JPfEUQIryyQtWT
9EtbtfWph6tVHImgxpBK4lOfOIHV4jEu29LZN4tO+NisSQ0vq7fnbXIfNtKFaDqvBM96R7Nkl4F+
zF82QDmqeYGOv16vravMOi8S+X2BV2TBOYbcazaxDHq0I2YxqpSW1+M2ZfApi1UlIEFPx6ZMqh42
qFYbesARqzYSu/o07KxgaOlCqdrgcuW2w7QKPUk65Cv7f0I2SSBpOn3vwVmexVhYdRGNLHYZDccd
6CZcUzZquhgADtnPGND6QnF5BdYmLHr7TApv5t2McF2nyZcWkq5ZXW9N+qBPNshcW11syUM2lhmH
gR05QJjopFTYeCSzhoHkwBfxtX/oWbnP+8iDqjqkKt9HeWJpS74guoLOmIYcVSTxc1FXkkNMYeI1
06MiWJ92ib/yrB52rI0rLcB5xNuzqJw9R42SOpUCFY8QkIwd3pY7hLp1G64C6UiN4jdB9B+lcj55
VNcQ4W6ujxdIeBo5kpTGh7IxbWVl73GkhMI0lAs4HBQfNGx31UG5uYtSppPZN3LYfy7UvgRB2H5k
WKHrLF/ZCzKFrayUANLfMoteU+uyLpmbbzNrbYra9F16+ocTgfajem2X9tua20oeSnKGjdMCfFAI
fNKzBF3PfpOk9cMbcrc+Z9oaLWrQbmfq6aqyvXAqR65wDowrqq1S9nw7FDhU3Hw2fPTzmLq26HFi
aXtjV3m8esfpLPfz3ty7MY3KWB3OzzsHiSYKlE4yhf/NGTmnB9US4N/SNIWdes/8C4gAT8/lSQNG
ovhlvVKu5jQLm7QC3Y66NUwNrYzA//DKf9f5TQPr7Fe/IkR5Kmm/6AuKr4BsITEV8PUNGLb1pYtz
1GGJCSuVlcKntgrJvkhWLnqJYACLh9v5UP2PJk799dslZecQgjhQT+oW8TxKRApBdU957vBXMUkd
J9KFVh+QJGzbenQ/PO1wCTrrNp1oc401yEizbsYcXbupoiQuLtjmBYeuHjJ352r/qR80sJAE7V1U
gpnkJ4KoNqoUAHGdQN8acKt5Ed2tqgqWW04sprJIEvvctnXcGBIffpCSYaBcvj3yegwnaNGub+6n
s+RC28baE20muX2QiunN+pe5rCwx6sBXNnH+Tg3jR0SO1xxWbu4d3suroSw+OYyuYIjj/UV34rHs
9m/qdJ8R13c7ZDbcaXUJNl4/YNGcPvsOLzgOm3ke90oF6KcDeO6ppktpYwV+tZMSemYMr4LKiTMl
XSYGVX/Cb//Xbac/8rxgkIBtRzLr62Z3848kB3LGjCTM9AwlLb7JQhfdPy+N2O4HZhHbgE/RYZr9
MWdeCo/g+hL51lznrue26YHpFoaSMGcWP+EjM+ybUB7idwZpJk1OhHazO3BjwSGWuzor1k/USTHR
9v8/SuXCIxMDGDjsNqzwNGLSCI+NeNRWWRDtCj74vNL7FVSH1B/hlHGQn+f6Nod5W4yhHI7gb5Ya
gNY5DEGWOLk955nwdOwrVPacR21RZT+9ka2b1Yrxpb7BgIAcESYrpODOVErAKR0FL7vxg0IvaMTD
MnCynqqaVcBO2fMsYAQhFcsj0/ltxE3Gwp30iTcGyQ1tQgYZfRCy9RgpMzkJXUpX8A35ef7mt8QW
eyWhdUx6SsXvm/68jCMiO67o9BqrfWG2XwPV82sqlXwDFFzTHP/D5zN5tNLAlcBmoyBTdXTLs+ID
meE6XJiUmjSDZZ0PGbAWUNH8P+izNMv0wAM3Tf8MBt/+LEEvxkd7F9M2z3dIhe67Irim1ReW1GJT
Vey5BS2mEYt+fYyYLogAwDO5cHgU32Z5sClKPzRAPAFzkArjOwsJZ2w60a+3G7sQJshZB7Oks6H6
iLO6GwmTHN+bnKQ2XdpjZ4oTnU0puS+2lyJp9T51TWDcsJN4T0lDcEI2ZGNRfRnMRct7+WX1Sf/o
avio7BVeKAtO8dBk7mfY0Dj+UIDPk51REH65HDcI9SI2klDxR+Dcdt+6DW2Dv4NIoR8PlaYSIv1k
2ZKgrvVQagqHPB+v1VOPXUZLlP8TlG3hM9cB6dl6VzvzIJAHKOq96NCoyucO2G1XC9IjLTOxJvza
y7PaRyuxCEV8R5BsJvBniyQqnRT4uyRYizED/8CPItzcFIHfhyp2Hm/gUMzR66AVN78y17MMAI3d
pEkaekO9wZILXPpaT+R8ojVo7TypkcK5Yqtqx4wsNRninrgs4UelVvkRPaWO8oZyMBLWSguxtxxe
c6LI6pUGK8BsRv5UXdyEpuqitTb+ixpocJ4kUGytQDr3t7erf3457Xzy7JvhmokN/v6ReCisBax+
gRh/G3zi3K8VoJU2YxpLAGTaPkVdnYWp+Z73ody25OvhkvVSCeGZ6+eiqYIbFZbp7REk0tUBne/b
+OUhLq/vCIz6jzFJhrMiqGW0z06+vbTHjD3ohXeBxqLA8d/bLiOLa+RQwRP/cNRiBIj1aUdhjFIT
6aAgSRy1UMblRijYDnVNOzUhbMZjmZJHnQufosYXGAxoEfHgZE02JWb691Uf7vj/5swRfPsMr8a2
G0Wm1OTOOAlVb3IfAptgk15mn9FL7ImQVqPwQa1hfsHU19ISEyfIl2cD7eR8fheBGuMyqYogrTLk
jo34XQodMcI8X2nNXs+n8y6+NpOOIyZ/k5VPKbhRCLLxF42c+EC+v2tA2+ujM5ebGFEH1My6oHwM
uVQKiZ/fMvzACq28dHMLEVYMSLrKvZl0Wug3R36WRpZE8j5MTzg7pVQeoDV4CZzMbPcooky0oBPL
1+EoRT6jEr0/2L2/cLPMubn7uj91XM/78AxGIBYQZdmFIgg4CdejdFbRWQzCJYoXN5u3p2Gwc3H+
khYamxAXnnuggQ8KEMVnY+jx+Nkp70qSvyvN+tqARJWjHExfrFXGWep0O/lb2yVlLaw0cRpSUY2d
OjQkkIAodpSYlGO1kibasuhslQdeD+/Y/1R/w6Ylf43leh2/YkbD7hAZu4/tVA4BTKmDhGbDKbjI
KhKNXhLEcjRpgJ2axK15TyNBLCmqpOn8O6emJHFTeXYEm9Tb+27YjaCooVs/2HXP58OdyNLmSw6f
753mqfP9tZMYQ9uvHgwHxjEqMvWtryqNp3M5AAIFvNn9rMRt2+CCBAIOXNHa6pNuAq1bAV2ywuBI
fDkVOeS4Q5xQRCq4Ibn9OqNh/b7YnB112Foo79PDJIpjMaRM3zxxXa5aWPEedyY0DiK4Kg+XR4e8
SoIF6EgrYESr4dASkDzCXZQs2rlfkYsrH8KPvwIYiZqi44nPnWv1CUAgb8JX6aopHKCUXiP0o86z
2bCLlqR6FujOSsBh3zqikiomcpRKLtFbNW4vj8VOhMGCaYfcOLjFR9IuYwRB6eHeonNJk01g2yhl
q0tYDITQgMHZ0BxdrzvyWbGmmRyTrw3Qn+ZCLXWrtTrJYcW55kxUpZejG1heDjHF+y0lcy/uOeYT
4+XV/4/bsWtbsq0ZWkaSCRGLtgUWe5HvR3FkxVpOFj9chfQA2OiIbf5OQXWk35x5wMvnU0ncgheR
g/wM9A75Ju9K+VtmXQ/YaP2WmMc8drQbelKJEhqm5Cl/Np/VvICCjOcUg0zcpZ1vzOlFMuFNrmJz
6NX4annmPNxjQQjLf4wkNHlOSmDeJC+l/xcnUO/kN77akiM21bacCwAaRskTBEwl3qgM0wcgfSSl
BlAZzd5//4oeJO7TnH+WMa55+kpslNeBAIfoPvA17WWsHabiJqXszIfupk0Sc2Gak/gyqfuIUX3/
ZW3m/pTsV/v33mTFD9tAbMma9Q62SdWlqsAGsHaSIqWQ8qw/IWVf0XFp0AnDXGjJajTw7ISZvfay
BPSXi+Ob4AO5+kupIk7umCwCCKr42KF8RB+F7Z6Jl6d1O2YHK56Ckrwbi6BIPUz+a4Dax17GeGEA
NCZQCSeVwlg9h6LjmJkEWrdBkwrg775D6dGRcyuCHwcVW0Kg7PG81FS41l85cElR4WV5s6BnF5j/
Iah84o5mSLkTVSHOWfZLaCU0EijE5jPIauuf5QZckuIz75KllxxaVGWv3mC+7DYLziwq7aYnyia3
GYJ8tdPQ2wT6yTV01gqWanJrhqdQPhBGLHV1eMXuzizLkEuElc7lB1ahD2B9z0PJ8NPiMR9bQYJa
+xwjzHIc4B/IevOGzp0DbdUXkRhi/GqBwJSfIN756alAimtmFFso9nGxhVGFIt8e3luV7eLxJ/AO
bslt+5J9YtaR8L+438LuDW7zytJXb+Gv5+Jzga8v2YYY7K/1sda/N4+ikeLOBac9YUwkJO5LDVw8
EYK1Hm++XCcUmdeB51hV/E7AIwbbzShoRklgWQqEBg/iOeQFVV5XSaO659qhIXhmr8d+V55M4EwE
8/D9WPMdYGzGbrCpkItiPet4P0Baxa1ug3ucKQho1NFhvykRa7oZuB627i4QUAKFOsafYdJhCePm
mHc7xEctAPG8D5brea9DXrp7fosoDuQhqulXAqwV96g3iZzqxtKDiwMOzNhftfPdgGQnCsG5QOc4
1LF+Dsepxv8UOQIZVPpiVPvDNsYMQI5GPNsHcE1oMJnjd8GtwBrDNl16AOg5rs7xDljxtZBx9p0P
2DFdwi8BPCUa3AlCct7A92jt+8i8DG2gJLu9EpryhKX/FgyIDUi9k7lkXvKTavd6hacsiF9TOG7S
NgM3c8v8OTGVa1cTM4QI5+qdOY4qtq/dVlJkx3T5ZmvEwhH2bu9Zs/Yz9pA3w1rhGBwE1KARINm9
7j4g/fJh5q6vU4M3qhFcrPHhWnKm8TrxyHre6qXqcTqALTuQUAGFYoL9rNlb/tcHpeFkDGi3fecC
onUukxuOlsyPUDrYY1jrKOoerC2lfkqW64gmjkXYcJYjqkzL/OxFykm1Me7eDy64qcd7Xff5QtW/
3tE2efRXqDKcBTBp4UtINULW/YXPtVBGNQABtbFcJVXZZZF+Q/7JgXTcGa3cag+la62Wf0iso4rY
PICWxdRholWcqDFICayGRaE5jX+gV13Obe+CqnU+7W4f3jHkclWaLLn5QayPbgo1zSbtZyLdjOJp
uo51ZNRIMq+XH3HzCzVmOXomzsyX8RJIWagBd0DO25CPGPVSgJOF8wpcbLM09YBw5SxLZpEt8Q8Z
fcVY4SlLAkj3x0MackxJn4d4oRKeK2Sh3e/t3Z4wVn1UmeZlt2Hisdd4RjK+snL/Pl3JX3vXhijX
DINA6Ubl9s3kS5GzSy5+SWvzOggfGiwcgCuOK3HtrKikV9ITlOt4cxrnmvKt/podBLs+BZStfVfr
vvcbSqIO/ETHiPACva7oQlzE8xDz7uEp75+aUhPYJWdovjHoI3+r0EYv2sOqeox5CbHZvDlC5N/Q
gHnKnuYcGd2Tv2EFtCASeRS7xYKL7QsAFJ8fJLnc0dabsGlKNWWnmBhkuhiOVxFsGIa2cT3Ceq3o
0q2T10eJ5EyxdqeQxSlTPhjJDwZ9ANJ38B1Ie1+mJOSRm1tmw44sn4skog32tmSADQcen2TWOdoE
3eF0+RC2mOaNBXhd9d3I4QnUj8fclfxbExJu4Lbw7aCcucUILZA9gzfJmIFU3vI0OoyWbN0KXmhh
7EftdwbSTBLiMWBRtoTBdIraRIBaJyNmvxpd89JWcD/71T08pqqq1V+uVADcj9iSitbxM59/QPWq
dSbdTD5fQAa751kT+2c6Q7XNJUHXDDtA1pCPnUQCFarKCAbIjjMOePPbM5L43k8srVb9RK1kedXZ
rWY5NkiqjZlcFLmvVYJy5I/uA6A8wA19t/wO3fjv5naNaBMvaqakqCcfbQUHeV/f4xUjcLi6qcye
4ABuSREqY2yfhAUuCgt8LnoV7KXj4yy3J199+oGwqzJRslbYwxaznyiQvvZr+rS+n+CqKV1CkkeJ
xQ68t3haTj7rq6A9p9pR8wfZU+CLMVeAh1vpfQdlP7V5ML/rz4yJTh0yH+Aefo9NOhpQJVR5V+i1
ovLgkOPwUmlr3bb1jMhN8H4T/3h0h1xfgmLvPymyzpL7ToMRpxcrCt5KujnpAiNyKWLJB5z9G/oy
s2+B9AN+huZwbzA3Ifhux31z6RWVW7HkVCb6ArvykwS2OqFRyCNRnhRx8UQ6/fp/Lwhm6ShiGnOr
mGUU+0KXCoA7F7nfCkWeDEbaPZCg2P1TN6BE6t8i9D9HZhB1vH4uNryzbyqP7Nisyl3hMaUzWi0S
WXWiOOju+Qj6lhnLHXeyDy8ahkBSFbfKBQV9ZY4c4prLboWO91HEDtKhEppbwhem+MLldcLOtG3f
UUZX/0h1sDoOHW0Uo1tEreQPuPnbCvHg3l01JXmgfBqKo7nfT2mi5fOu8CLXuBDGR6K2S8a/88Ns
dmEhgOnIlh6OqGAMlbhrVdAvRjzPo1gR7JoPbMruu7z0jtLchwK76jqVl/JpvRiwnFhGmjjGuv4K
2eWypDOciSMfiyf7XKJVdmXaiH2u9DDli1gbmrKNDUAk4X9QkdKnDkvn07MdGDOronHHj7/oVKF8
9SgJXGCd/4byzdhHhJU9iTd+RJXVe0eRCXZsAMMbyew/DI8KmrNRKb7AEuaCLyVmdjaZ3y9ikvq6
a5INY4gBe+3K3myIsABenmG1wy0+QQRmAnx8gNf2ZghOpWYo2CpvSb4tbTnSsASMEelOEwUDxLvN
hftzVyWuw6cl56bXwf/+Iz9LksMB7YpfCFJd4uSWM/AMeZq3fDtZEqRtCPWUJaVp7gPnNOI8FQLO
Qss/RuIxTWKP4D3rl9aDIIpu/PtZn1sauqErHw7HvhPTs+ZLK1p8OMRyV01NPrqAs3G//hfCxFA4
t87K6Ht8j3XKBUzjTApoXPaKqvs2fJGP3Rp+QJ0lob5AzZ0ZJldbuNrUcn1fFflpRkrKFA9b1bfR
qo9+VN6OVlZA7Lec33D98h4DGAf2NLlUg7eQB/4lgSTAdJXtaUmJTj1+AekHWerafMqe9e9lTk7J
g8dS1yKP4vJGGRfI82sjKpW2Rki+lECjUmNuqar2tf673tGFyaFkMyO72co7aLrO9rh0vzJmhRsb
IvPkRmSoj19AiPWDqO/ZbFmJ5rAtpHJJ2OjCLIPMeeSwwR6Qumt8tzzJibxTwjfoS35ro3NOrr0k
ME4XxfGKvgLBAqfvRfteWibS7gySPQkQVIIHP3aqhg6Q7M+dwOqihSJ8qvMH0w3YQYk6OaOhjwPW
KDUzVClL5XPiK3OD21Sg7y86y3NLZxE2jPYHfGX7upXCRecSXcv/lNYz8jzKxljm6WW2ObdX6TmX
J2suMjqyIqxHkZRxvZdq23OsAthSpOtvS3JM9xHQOpQ3peh3jlKPw7BNF5tZlFFRMj4qlVlPupBr
aG1s89H9hF4gJ6OtZIeekbs+19TgvFNfi25off5J2BoQZqiNKPDhOYnAx8XTixHDSQwZJqOi0ZB3
g1sS2uqnGxgZ9unl6RAVQDHLKkuzSrG25yC+FjZMqyc1SbJX6P0oQnpEU9n6T80QZQQ1/jb//fo+
Sux3B1wQfb3NxHw7zfDOd2PizQjGvQS0iIUgN/EGhU0kuSX3nQIhiCF4+b0DefSfDFbg8fGpa7+Q
vRj/G5ncevFQ40ev1sijt7tiLcw7puMhI6nGzYleKNpJduqfA4lDRqbwcCte5u0u0kad+1HJgNIe
sFrE6XjD8N5E8VFDJPUEEU2HkGJVdlRAHI37Z6Am0SX8BpXdNaqyHdqolUKLWvxaeySjJK24V9Re
nSItMhdZwznSF95tR1ZHuxQbcQYxeMzXK95hNGjx+TybwjA44WJDK41hAJPqifvDjwU0908Yg+1j
HJZsaMOGCRm+JlT1s1E32CdnPFjvXB3HlsBPB4BB9qQyLWwhZv0MUOc37BN9SZaqOjpEapaGrxbt
kmg0Gi8nBwrXGv/ZO9/ienTCcFLFS+WcdjcZsAdrkeGf7x1BUWzveKngoc357kP6Zq7sVhbGKDTn
ySvlWbS9DSF8fMfk7lgJTAHpRW0VEEtTVloysLE3zTwPqhK1ik8w0U+Qoso1KWza4/RYpDQh6Rv4
bhKIfEtguYaFRf38oM5H7lgfs4AGyGLuImPNfRphs+xH+19TjpT2GKqShjNT1DhVINts0YRM8QPd
gc5U8QmR+3Qd542R+aVyVhIUP5xPCVeyPPrVfg7SFOJ0HnUc43Gq+Bx4Dwc6MRIlIZvmFq+hU/8/
FtyEU/eEH5Cgii5hD15cE+dIxwSt6yYMZxfLHKSOJmfsNjiie+rWRWzbd9mKIqLS4ngzSy+WCyPX
yCt9rdWbmxSCt4rcU3Nr/l0LlOd7WyyNDrr4mLxSXbUyax2YI4+IxDzcn10VuPxsk+kDxu5fJzgx
iH38hohuuEuaaDYHWi4EtmBmLCKIfEBDzv8n1C+k9qaA2YZnZvtovT/g7FbrF+UDGSO+WkF8j/FS
/QUtDJIAZecf83vtTKaxZsF56NG0ZsgiOkCgPGm6isOIqLsbQhITqu4XzEx7IXb7h4ruQ7BaTtUs
VUmvLj9LklSiQRU+ZYzNaf6h5XKHS6XdKkou8MbPfWlOaQbSm+0TnZL8Ab3LIQNeA17ycZgEqIGL
nBXUc5tCeq7ntaMzd53ZHEnUh8YksmPUV50jTckpf38ZoMKMjzouX2kBKz3NFwqHwgG1BDFoMjps
g+r4C0yEQRrcpCiyt4VtxrYBeN1EmV3CtpPU3eSMSP5Xq38DPcIG14frRbA7m8T1YsHg3Vywd4fS
M7f0XPmZS3MpqxTa9PvjnufF2nfKrNPi8kUb895GeluxSlbp+OckXmQZq9LELLEbaLVeM9cvVfWU
90A30aDFJnPr/uM3TDfDaGRNL22Z8dnKr+xvT1+WzfRbnVr3Hy2TEkKRXbSp2IJaDNvmHEYUdT9x
GiPSiKM97WABdjT/dzb0X+2ttJLxtzC5lujESl7YU9y+vTecijh/aVdG72phcIYkCPJZSwSI5c3F
tn5qqUYhyM51yqKxnYY1eESWI4ldqxZ4ndT2R4poPON7Dm4eogYfQBJ6wCim8dmTx71EGWqERclY
Kf2+Jfifs3islazMyyU5FdcWpG2mvQtU9ZnXTes3Bya+SkKtQCaqBNLbmLYkW1yLiYjcWyH5lShD
EpHNxP1ifrasTGhcnmWqGo2ykwZhfBzwSfMDu7oJB2txOOk7wMMoGwEfinAEv4ok2If1hsLbe+S3
eePK9ZXZIbRrGERB9xnDFfb0Y4jw1I5MkrlASIu4dtYeFR13nQkf9Fy3sM3hjv6YlayjZwx26+R+
GuCNj3cq5ABARk4AVsrTn/urdR6kDJCeIjUllrLMih+697BVM5VHoTraVFwffyOlR6g3wwzLySK4
0DDhN2Mri02M4Ne7iWc8vZwHoyqBHFtEggQCYcMY8HFuN527Y8dlL99xcM9Eh9S+BI/iDxOmrIUJ
VoROAKsT+VRoHYYnsyKc4AhzkUW7kDe+XMhNWo620WjZdhfpu1+lZBFMmnHEc1otYvGrY4fRMqSF
+sStBO6/7DpFR2Ps3TW14rnN6mgUBlgd3QQIERmC78lSpyvAP2Aylt88vTdSMktjgzkXd16BsWnB
nbMUYwsSsoV/u+5nDLrUpJc5H+kIsbGILdThtUGBi8rxr+NPIs5Cs3l9uJlLIdWLMx9ffDunaS+l
W9OFRbevnH32mV6nnKk4rLj17v0F7qNEGcyntuKvvgBe+ksz+FWP/Utfjizc0HdgnfmVck9BzT4a
SiLbjPo62CdDpHMVnKOjoNEyWAj7rTNiBw3inqbWnAq12P9FAR+tom30iCHn+7uPDdLhRCiMzz/g
2gx5Jd9MTYbAcOjkl4OGw/ZixKydxcfx0dcFU3MGvrVaZjAFf2KeB8Y3aQRPqOZS2Na4Pigbfrd3
o4pYoIaaTBGfKQ0V45YKCbeAuNWQ/iAfToa3ggJNYTrXkU1gT3F8roTVcJzGPgpE8limxm2123yy
oR85QcP8UrITowwziMWZogz06nJBd2JFfSI84v4PvjqJKkid+cTePVLlq3jFXWv6yFTPoOG3Isgh
K3iNpH/gQ56mn20p52aOn53aH1T6b0u3+N2rJwkYnUSysPnjr9zUt83y869mz4nN7qAmVthg/JsW
y0aTAi9lG+JHZHfZGjYBWMSmSWsHSHAp7FFJ9Bnb/Eg9+MBXPetr6DR5oJiqfnj3saU+H7a6EaZt
mSVTnxmXXfXtfo/y48Cp+3VAxZB8J96hk5qfxYr+iOAc3AvqpxKLWXwZfXGl1WDecIN/SNYOxvVM
bGMRvVm14IaJ7KHcEvXp4u2bZVyphA9W935RMPxvdjCrw90FbivlBaLZ8JFE0COyZkF6oZRMuuzk
KCYc9lQi0s2TcatEz3FPe77htCyKraF5lAOPsSvOA9m5dMeqwn7npwIU+Q3UqZoHGWmR7evTG2EG
j+3SitB+DY92tcpIcyCzspFATVh8jkcqqOz6W66w9XZW6Ezpu7/NSX25airwYjtqmiQPi9k7zm6k
Hpbd8hHfpF4QYzpmKfs50iXkd78aQtlzvf0vjxI6mqSXQ7Uteop8rP4zBOvY0LXwCWXKgC+W848V
9p/d3LdlWKxvHPn0PuvVuFIrKg8dw89y1Nh1wscZ05Gw3WYGVIynABdcju1llGhqaooW1rKvsNnb
ktvdf0gisvrkn2hdPu40J1jPwAIVCMU6XM63Xldh1XD9KzypWzjQ68bqDrfXdTmMehDd8GCr1qOV
osU9QJfOWsqKA8WOga9YoaKk1+j/sF3KYYcPbJhgThI/UPoykiYf/KyR3mRn15kLSvv9/+wah8s4
3MC5qGgrWHciWN0J5nG02zUMdgZWeTJ0CRzR7fEOzPxz9xR+U76SETSuJrX5/gXKfzpTTg99gIK2
jyL26HeiNcOq0sNeS+gbLLxk7CbmP9vw0GFQucTYXpol2llnp4zLA58bY4pIoywHF4r1xfNwJl6W
isw/DeN4EzllgepFPoLOb3+jbkKL5YWsb2KI06QxvK1DT0QhnnVXojPK7oPDvDcnpHkpqizjjqZZ
MfHWi5N7yURDv0XQHovIYcUiZVLLWkEiIZ0GQB70fkJzZfYA4O03RdJm0r9bX+NPwSAByuRLQtoT
CrbvhKAXsxWcN0HWQMGQFCKYUwzUDzsjdxXlVJeT64xoXr4BngUmd6crq79vidtjD2A9BMgtY51h
j4GE2bycFXc+OqzS+aqIAeI7jqsBgOqwKM415oHLegN6L4tOQgBSsaWx1cCQopNTzRByyfqXvEhu
JPvH+iuxs1v7/zZEPxGVC1SlwOpwiLB2Nz59WzP4fDlN37c27iR6aoRVSdHvTEQuvTO3kkk5LtL/
jhWEmFGH8zl/RuJ13tKvsZXwEQN9wrJduXJPx/uL2KB0aUZtTghz1C7YVYni19ejwfAbipwy6wb6
GiJiuhNz+cEgIgTUoxEHMkYmduJBCBRGhZq4OW8liiEdUTKlHGfvWtxPn3ejcn7nj758/S3xFtUJ
PhKA5xOJFBtJd0FOxDa3Vph0bSsIVBaC3vM6Y3bU5IFowxKWSicjKVxRZY+2n/v0hLWoGiEQylMn
qIn6Sq+8HFIB+OMP/e/hnKA1ccYgOSTbhLg72+ctm0QEbjCcVgJQuZVLgJ/PYqVzouSeFobjaPlG
ItXRdm0cMwlTinBkeBoZ06iyER5DwbRAXVpEyC5v4W+1c21otf0RA9X2qKx8M5hKDXlPeTCRxA75
a62bC06QZLR2DPRDeZ3rSsnDlckaeWgY6qTr6bGl9vPXJUQrMzUfG3EZ/c2iY2sSM61j6ioKqOcC
tqi6373VfrwkVY/lSShID9BddXrQwUKeinvJ/4XLmTjHDPM6pg4wSpJ+Rb1gGcnIiXUem01QdbcN
woE4reGXvtdUYfkJn737aoI1FICD8ihodLyrhoOxoexTY+GfFWgFWpeJgc5YTQ3+V/WI4YtlDDj/
DbQuxbMEhugj/eAa1HyqxlS8xAaDeJIJbbAkfl9zzL0XTZ2SCVcyeIwvFBKBPdb9MsoZL+4ZDiPE
qhi7CD36BC0nxkToXYUzg5IO3IGrJgUBwMOgkw8O/SLbkfGuRUHhe7jTrNQ6gRk1fNO8l12TWczI
xfVwbr2jknePTZMkfR3jhUyUq5qq16yHRUnMrBFDk5HJQUful6+oXWxPJPmwjnIc/h4lhkotOMoz
UKVNemgUyjzDgrsbOTcDhaf8BBLzLACnZk1uAJk0scRV9IzNMx7Ey9fN1iz1FMTghHZf3bj4PZ0Z
8wWivyxj60PBJn+m4IPOR8tdgBTR9zWW+Cz6K7aC83/PHuhfWgMw2wFKPVcdjxESobrS3j6eHUu2
akIwTEo/G/7h9QPA1X+9SkoZd2GvcuePw2JKi8vVldP2ztIbUgSZLTnf1LiqN1JGSb9CoKvSWa5m
KcY4Anv6jgy4izJQB/r3Ek5x+ZqmdSZicmYbDQGo8hWprZSPEO3FBWEFy0YSgXGvXWc/XN0csQNm
1CVlvj6pkdBLiNHEWwXj0QRKsvTom+bi50p0KykyOdEMs3QYU1PvdHFiXvdUmtcCWoc/m5DOMn7S
9AN0IGRgh+XORRih946kQWFctHxQ2KLKWcF32rrhbL2jX8C7Tzd9Cy/ZQIBWgh8ZZ90DMUWgMpUa
PomdoKdDzyIPb08Am9MpELKCXlIF5694aVJEFucKuxq7MHgKKGy6qHMMkY1OKQFAZAnOAGlawe6t
0I+jv6/p4+1b+VWWchebx+C4kqjfZxb5gGjQPwdEoEUhM0lZJ+A+kuYOiMLjwklNntN8wbYJky7M
4R22F0Ga6fnXIoV9OpXiAdDYq0+IyQ5QuceSPPYlxvQ0lhDPhMCEnoCTgi2tLGKb2CTxOOPtvfIn
aoLtYrwIgkc7ZqPqhn8y1v2e0MIUGyhbl04OeVWQNVEaBMuOfV5w1VbHA7Xxxah6imWRKWRI0m0U
tIK2IXudBpOSr3l98w8GK7G6cXRhqV/XpVzNoYPLSGvaRXglYXTI/8+hnzS7OeKFO99GOQBk4Nux
lL1uldR+G5Y/F+l+zvhdfMMk0LoVP0bZV+YaaHwqc4j/kR6PmicE56HFueXseoveEJ2ANQZVgbHY
SXpvx6Vlct7c+FiMPWluqNwvtmTvsGlS2w7ZuXVb1FkRimG8B9yJwrMepsta93fI8GUnMEFnVCT1
nXM9mt1CNMBioij/L68AXfFE2de4pmWMgKPIZRWTUF36deVkqB0+lId2Z6ITvf4h52iSvfZcwPV9
9UvLEL2bo7rfU9TIl3FaCSTZJ17WICUDqtzo1NTLzYG4vCU7bLSJd80QRFdCtUnxLSECFNpSddto
haWaKu6Gg1h5ZJTTClp4Ivwjn6wFVXslfk5XlnafMsZI6GJgzG+xXrHjjlN+f2BkhEGxT7bNaG7D
N2FvRwZ31hM1IWUzFCYY0Ijk9Gm3bSUOCb6gOQS7NuPTGN91LlODzoYN2aBUPcwypugk5uqWD9dS
P8D0f8gAyJESrDbbnBw/AA+680sP7qqf02BIMRmQ1+gjMu9STu8qb0nU5MVTegjr2wt2gDmsBJDf
MzJlraICkcyqnrGHv67batcDgzCPf8lr9QmrDaDRlLGNE3tS+5D1Nzy1vLmtLhTJ1kkbnhcFnP8Z
j19M1mpq7Xjs0f0SFVZ4RmNJgTS+GIbhsWwM8m5ciVp+SlmkntR1hP0gXSNdQbc5sjAe6BdS7NdY
t/dUK9+e60LsMLcTZBo+VuvdrGkHbv5rI12H7ky9Y+2hagR2z2Mi7oqysrnBP8/F+/lCwOD5yOpv
k+7xBEQP+2dysTV7XoNGhQxin9SAQCHNQdbTzVQbZtAZZWWvC55Nh186BUDriWJ2xEIDgLRuuhc+
bj0DSmYn94omR0zSYE8FLvxtMwrc3pINwi67CnTkxf2NKu5Z4gVWBJj8tqMoFf6DP9cvleVUwM0H
0zbSddfyVQk7zyNinvqgcP91WDCuGOnG+gI7eLu/uZfLDbhR6WxgZ7lV/Ek2j2nCabckYvTr8B5g
dZW4DJxSXCKvOQqHwgAbNoH9UrJCJsV0DiKQtyaubE0CYqjJ1L1J73O9Gua4lc1cQbcCGNiCWoMq
5+o7+/KQoG2VL5NdY5bNf97Onlq75js4+APioPgJAVa15bx8YMqFxdosW9UdRsrDPSlEcWqoKwVE
a1FDgkkoWadfyk/ux4HFvHxfnw5zjoWt3HiuIpTFjbOPDqo1MrB2cEXCqPGex9S/FoFVLph6im7o
mIzvySiNjTFUz2dM66TLWBfmlkxBUntlYhARmBhtJIwkWX9FCYgZUl7ceTl6c2a6PXEEjFD/uGOH
4jNlzCahK8EOX0KogRF8salQu/hqv6cDF1lJEbrbvKxribaGy7vkmVCpsQODBMGC5hIsGU6/F5HP
UQIS9XyexjZKrndevgCRZFTlMZPNevJThr7xd6/H10KKJFOzKUlzxr2RD0W0Kq8GwTuWQbtI4mFA
Q1f/CfLiZ1sJCzG8oNrz8c0+U22R1Ief6/4RXSVbuACJ2Q8LDUdKRQG6/7hcLWtyUUj1gDzMPHqG
UQeJ2qVeLVrCz994tMX8CB4F9L+VQP0C07iZM3g5QdYZyDKaTWWCRSbdWu8OXo7o8siB+hbKgkfw
RFJ0dcJdcEjksdus2IEvy4JIIrx74SVDiWgpdgs8QmMVQzHeLgEHeSHpHhIPH4sWa4B+ol8iXxmA
tw6d1oXP5wCbYpolFMiEEeN0oZ9NTo2TnYJjt0vel/62j0uRBtvCYE8WS1A5iNz9RPqmSMce/BoI
IBu9dbETdghiyRZsmGv/whiVExlbkFEwTGkamxaWJacCEldma+G4b/SGsmNMoz0Ksiyotn6DdLIh
N1PJxLwGxwhEgBP4auPJSyJkyOwrm1lWC5hw8DGcgfFuoTN+OC9Ac7zQ9+1eU5zgWSStUIOwmAK0
wcq2C/79QMavfAy6sles+CYXVowRaHldRkiiDG/oEmCRbv5E9uyc+vfAt5H7e1ME1eOx7LRiT5F3
nlQPpK2VbKUW0Vkj9X9elxtRjt9IXaX7Y/cZBF7/XyNlo3Pa5Cui3Bv8qNAA5oWFEyEE1Isx3zhy
sxlKYDeTQHXw4DBp+vL5C6VAelEZD95qF7aYSaWjzgYVNu19RIF8m5afMmOqXcD7gCaCktASK6wG
grooSbgu0fygy9O2IPdtRatMK8JewfvwETVsJYGqTlS+wvl8danbtYAEJc9TUo8rTJhDahPG4vCc
PzPbJ/qbwVHuwONZSbMQkL3yWOqLftqA1N8548g6phsqsd2YaRfSwASPUP4EVobH2qT6Q2QdBv6y
ZqajPQsYnEUbhaajJC1sVS5YM5R8xTX/ItGYpV82PF1K5TaaPBpyVS7TNS1lbY4NoHFCxOax/qDp
SyjiW2NpSLBPzONsn9e+nLA4zcwwvzm8Hs+zPxRU5tEfnbJ5sWrHYlj5SUW4hBIVIDL18lqeVbZN
Q0RYHLEHJGs/p6BKqVAo76AbkCkI8q/221jjrLzVdCFfMqxViy3CKbKhWrJz9171JqRbzyt/1Oj3
kXv8BjQ+qU1ABUvuN1/dGke2KmOo9lIrgcNbQKEZJPDbG5pS9PrLeZFj/hpg+Z7vpxH4t5LM5m7F
m73eKVZo5Baf7EsAVxhNOBzC+jfkHTvLaOBs2XOulV8j9lOTYGkzfYh02Twl1lVXWMHCEh5LKaBB
bSW6xdAvfH19e/xuwEdEJE+U9gjPTm3qyifJmPc7AyN6EDNmi4tvWSuCk0aOY2U8MY3KpkWG9+Wj
CjZ2Slq1fJS7AWiehFOLf+VpArn9OXWF1+6GGqGKTJfzlnvtpMjLq6hgLUsqZAFyVowFKcYiy0bC
li58ICCzSocVEXonGnVQ7QwhC0RooB07YSCNBOq3nE7BgjtO6GTze2sW7VbW41nRAf1obEjhyL9Q
MM2wuit0eTpqpmfBoq9bta5jdkhJntU6+1E1P8dPxKJyW7HTp5yQVtqL8gALl9RTe5v0krrs1d+V
tlq7LvTcr6a8nm8dDEL2BRXKBEHaD49QrIau2wmqToh27Tp9RG3kvjUCYIne7Ejh4Kn6h7xz5OO0
A6c9TU4yxjkZ0PHMHnH0IqPOSy/Bk/fN7OwLNGUwsdOJhXY2ckJVoXleHZ6gdSGqFQqSqQYBfu95
Bmo9x+UCUcqXE2fxphhFcHUvOdRYssmXf+zp3aC0cc1nR8EVqf8VtjWbr9Xy3FzWlq/QEu6xt1j1
3xKvNX0XkSm6as/udil6h8fTvNpWD9OWo1E7QO8Ji10Vo7n6umaPkzIMX+i5RHXg3rUEPJj3Sb8H
vGZINDAoXRJrsYfYpxiwPikFoa7urDj8FOIu0dWScK6FVtbRSbk9ciqnrxjNm8quwPZ0QzMM4IvG
gBoChuNTRtLjTConFnNIkdHt9Kn+Mi/NCwIsGpDiyCj1ufKe3JOhTSAUYQ2gs5NQ4kMx+X5QI24V
03QLniD4J1gSzMiH5Gppy3XPddqc6ox0dBHz3iBobCzYn5Kcj31x18tl/ncZfbbZjbOZAO1dmrLC
Hy8QdXK7TtS0P6dtNTqxVIyrsDMlEi0q2Z5IAoYhBQPTv/woRBWD8SuFaJzCrblRJs22RV+fPnf7
dD6hI/RV14EuLMd2zgUTCMONYNR/smhYIA/Rmjy/JW7WsaMP8dUQsIoyMV3DloahQUvIBubq3G8C
xmL4jFPRzu5aOCHCJ7idBe0D4M+AKW+3IXmvM2ecZdCV4Ltst8NVrmvd/9aPgGuCQ6o1PBl01JC5
cMeY6NM6pe2M+n7ITXKk0sLxow3fef58CQ7ap3dAyOtaKtBphNDNNceps+GwjXIsEM291Q32mJkG
aW8JQqeGGZkymMPiTKoCdjVtJl+iENDKCq8CmHuWUSfKFVB0y1uXWrmqDigRKt7r8nwIF6mTC4mj
sNNgYPbN0XFf0YU/hqEge+zAEGcwHNnSfPuJIdmPTqlZxIn7a6oWMnSi/RQIRc1LQDTXsNmntQtf
bwROPuBahfIceEASclJKuiYh6+8OA3apUI0cLotdhx1ZQUl6rlLApJo1cxWoedtukAHp2Uuhc/Si
ERBhc6W986Zq2AMiG+vyBdsKjPvdHLHNxUj5n+wejU+x1d8bEATDMpJrmopDnuokcYjL/HZiO0Jj
A4j7L5IjIP0BuVB5+s1HYWueo67NuyStBenogFNhsZoPLyhZfQ6MXT1jnw1dMRjWcDL6Sdjf1mGJ
JAv7wxYS5pnwDiwtdJ4WE0WD9QDjRqkcCdNAIDBbHOvS5sB3MRyJW0fwMlJK8E7POqk2GJUq81cO
W4K2HinpVVPttn/JUKZp44C3OanUCdRctT5WU5io+sfQOdj0zu9JaVWrHJQspv9hsay9ZrWeKiug
tEFpORIHvD/XJMHZn4u748YSjOBEoPDfJM7hyX7zDwN1SJP9SpEdjcY8tlfv6DYnXkKMZLS51iwz
zJBAlOAM51yexSzcrJEVSK3+PxiEnLny/jodJlnIEDOZyUz2CYRx7yMVi2z7J4mJx4QmJjwjYYQ4
keCmOJoFt/MqCixkhXnm7CQvTiEWiczd7mFuQ41bFk0hnNzOHN+U5VsCG4cbXlrq/Kh4UP5456F8
AXldqC2qv/NF4fDHLVMEGXt9YY4NxsBfhKeGdiZQ33qDfNr6ty3lGJlP0EzbQmqXC5VQHSU3ugCm
3RJqZeSIeGnkJjMnO0atIvEgtRsqEMAdx7/WMmO+QjzOfQZ4GwAiKpqYJaMigEzlmwJNxZsizKdv
UdRC/Xn0bcC01WXrl2fEqosDPKCI3dBst98f2SeEVztTPwIy2hiAjKXsi5ZBmeOJodtZC92T78Pa
LfvEkp5wT2kAa20N1u+CdxXlsr+P0LLq2lthTRAy3pddXwiiicuV3+xlwfWjS19brAn7Gn8bVROr
OR1TDam3LkcU3NSlcPy7GljhBcbGZlKIhmpviHHdmYqyBThixGij8J3huzLQ4WMmWI4VCuS8fZ2f
ZPbUy7Z/yXJyQtQRt6Vt5kwyfuZYUZtHMkFfL12cCJWxSlhhmXqaChJvGv06Tp7lpmgV7VFb6yj7
jgyHD91whk1bIrf+JxkR/AQ28zQ21i8x6GdIfIq0VL9muTA4h78gFmi6+bXPUIXa6YnlXWQg3u0D
L1NIEs/j431ViwTvuEoZ4nWHHpzV3Kib9qSXR899dPgdelMLk6MPf04AqHuD4YlXd+M12kO5MSE6
eJsV5m/cH24UL24+pXV2zHaTTX4RtW81NXuXDM/d0XrygfrImy7AjqltYR9TJKceCzSesE1hD5Os
PHuYyBeH/dkurDLd77yUN5/LjxyIuKt05pRADQXauLI3WIDFSeqWiVVwIyC7D5LeFfFt+gTLSTfY
Y4Nw2vfCEEQTapEZTc20piExl49DpkzfGl2eaHJNYKxkM9WjW6itxdaGf9KWNCEKXQKa728HsdB/
dnvPJgDbiBazfp8rUW8/UOrM6Ykq1Vv1gDPkd8EkyjvIXTI67fEaFbUkEea77mClRntoem/RPejP
tvyRYoNixOsC9zb2aWy9MUW6FWKHyA0QzHmjP8MHEn6JPE/3hmVDmj3v/S/vLTbSrVldFMxA167Z
+UmmQDfAWOm0mx/kj8aMhFyKcIbpb3yorXkbf+tkEja/TwXC4Q4bR0ZqzjH85jmiZizpV3Dm7qIY
7L1kLjMPb+lOrPZLGhK6vWeRHG83TWgOUQOYiTIOooRTZx+DvgD/tMk2hJYT2+0kFX0rxXltH5Hy
P/1/M/jmB56wty+3ZZIa6aEZ980fcQORpbk3SGUfeJIvQagArup0kTd2TIDvEvTpgDlejBoyxlqY
o3wfR5pP6AXlYXvjEEKI9elw051mx2YTKgWg3R6h2TzLMwe5FJAsnCkzwp5ok2mPEftaIAfxst0y
mn6e+U4bWV8lQxz10zsFpQEzUDAaAUjeklbsv+JS9B4VYQCuW3EUcpkJTq5IAVO3JranO7nsJIEm
Hytd9oGhot6cHDzRDboB7zm9B/DQxhEsNtajSmWPnIYll0QrAf3EATfkx0Pz0PNtT86tkA5SUb29
lFofQDiYelFguEDtJmcksq06+Kwj3LXprQ3JUXsbVdSWSVbzNLlGC7nEr5WG9NMM0+JB6XyaS9OK
VIFR0oq1Th27XAlly4FrYc3PuIXaOdWPnAZxXLn+AZ089y2krofAOTodFKeDoiF4ai2PzfIrrF6A
UGuM6sEIJVuKP1ls5sD15m5DuDLWfsO7sjfkB4qtjO3p4kJHUJ/Op15e1AAqKIKSSxraK4Swxka+
OZO0vVrxt02Io7E+9S4ZNXK2/6WM3Y9WWQdi34HYSpRRtK0cZvo5Tm4sWjRllPmXulHsd05hj/rB
ZIuJIQ69lOc/qd3cvgfAno55EosVen57SbHjrFP47xZLH+NUe1gjbKh0OHBZPRXelMR7nsimJ1Ne
l4GwRw9HKhQWAL91QI1LexE/z6FLnCdMjtx/10SpulZxi+l543hUgQv3+slIkkXNwS3etvYE0Mks
t53uKNC0CQgVRJh6mEBX8542mX2DF2gD4RuAk9UTFmg5mUT+zaKe/TY3UxmyxDwjlQPAPPi2iQwt
5Qvnx7DNL77FElT6gvjQHZ3cqI1w6bgrpI8jksqmw48yJEBTKwC3ldRhHbgXBAtAg0+5DN2KMZr9
ag9dp2OlMC9R1OA3qb4Z5z2NHsIbA1prXJKFnAhqs8810wJDrJFojtZYLQGe1p1PopVjFowG/sYi
z/NjDsFTwjc3AkzIl5FTH29UljRwMAlMvQyB8eaWGfRxCORD6lp2iYNxZiYjp6jLUKuzly4wYj5P
2lmzENsifVmA+OW62LZxQHKaR+Ppz6HPiuWcYGLCXgb/exIoUoj2SZaq6Ih2C4lDgkb9ScKGGTYG
Z2YHso1DQFxO1nDbuliNmz6hOjh0FQppMwUHHkTMayshkJH82rtosl/WXYwh49pllAUR7edXxXmW
YtrfPt47Yz7u7KwHPtKMGaZ4ZYAZJ5gpzyNJ789R+LO+y6mpa7M6+Q9Z9Xa3wqthRHGA56QPyj8l
LqsqrtGY2Zom72/KigiNN16v5olpwOapDRZd3DYBX806NZVga8uYZ7r1kctm+/tADNSyT8LHH0Xg
JZ9c5yu+0gtitLmMapHxDXeRZix7Qm6pgUsGW5W3+V3q2XjZG8z4HnOOQkFTOSQSJWvQChKi2jrK
PUZ8q11oIGstbfWUa38Gy60xXphqondRTmjBTmWKj94zjlYSDRpAh9MSHGhcOw1/h+AKYFAX1t4E
dGgtn7XQHUy5rbQzDIbVp2RWT5E/XX1gsMwiqZsEzJ8KfoYqpGbZ6Jnlqs5He1LmkcVluSC6heWH
d6WltcGvL8jhyZO6sIUcwai7g5tbZAaIFgNdEhe2d1n2RZncZurixYlV9+sqw5FR7sO+w88ZqB94
3qo4bghyXa4T7i+I2Oi+vcwpYiTR8Ji7HWHwrI1iM63WOlXfODKYGZSP07IP2EAUQ8ICpQGMbCeW
9EJqyx383Kt4UrWKz6QNEfutzuN+RCiOuwpRUmtowLeipM9Nzq78FO5u1t1i9KjZi12Hs5ksXGbu
QkRzE1qsqIIuYUty1MKnXrMfkwRNxxyKjv3qMnQ6bavKcSTxQKuO1Pb0oeIudMLz6I2HjOBtTsDf
9+0JwFedHVq3eIqsWAzpYT8+FZxBE5Iok0pzDxhwRLo1OorwdHPLjLWnANJneHG4AHlwbY9BqgR1
TYyN4vyYaXfikXq4K0TAgBG7kiL+Kx/6tO36xC5O1ujZgQ8Lya0orT4rUyFh5/6R7UNGa10wnMFm
oPfPSrQvASpc0AjUXSQNdDeWHrq7GrmRdqr8UIUq9xaPUcmlIjJfVI+ioY+fGKZljTVtSveFIEie
oTsH7EEhh8yXBc9DzQJyEatnl95FYYc/o/6GMPFV8Q+x1SkxJj9Spc2vX35xpZ3u8uLYYAUvcxe1
M7Vx5+E9SXHVP/1LMJSNebW9RPKzjATe5l+qzNAtOTToVr5hJe+BrakruhbbmSv0LnFPbKIEYzNT
sN+YiZprJ44lltfTV1fkN+Iir/fr9mXgYVoDR3V/kb7R861gXgVwm0Gwj8EASeVmmBsXaGawWGmv
h8WqpR2ixSZumBf1eS/w6K1HFmy6kcRT1BxZZ9cFFQ0yq4igj0Te1IYUb29oQUY08oSz4YHIucKn
ptUmi+SE8JoT37EJjgJXv4hU2knMduKSRmeJ+SZeqkJuXliYkA8ZFTYHEPxuPwj+fflWjy3Jb7j3
yKLtV0pqTeCWKPf9107k2fhZBuXXzQoAIuBDqKwjf8e9wuhcHfsNJ9Z/Im9jCRwL09iPJy0jGpFO
SouEluBvYnr/1ThtplCBsFwQC5NSvNUcUadZQFctmD8tD6lGBsIfQxWyX4o67GAZ0hdfnE6G4seH
aRlVwpF782DjhDt1pJBVrOaWpnvxAsRYazk9UAgmKSp1eHaqSYcO+rfxDnKmmAqHTRPSHgcTl7Sa
DyyK+yhl6ZJdTJtekLI9waQIw8IAwXPeWEVRZI3/srkMU3UN3/Ja48b6Al3ICLK2TB5kyZvKCUAO
cW/7D14wQr7XWxGu5gvsYMw01Y4XYI+rVYWRm7yH0/fFs0t9JW89Odr+yQ0hienkuxhancoF0XWp
tw+FWgpVLs1SerD35EYVZOPbAh49Q9Yb26M8u4FGaDZfYtJEzc69eOYTgGxJZBQf1mzMBo19VgIF
p4/fW5H5+fLll5YS8AiKW5YyWYtutb+Ql/cU30F3neAPjFzBzKP4JKTe0eBVXnqPFJHiYH6Jr7ze
mdTSCmXsibtyhc5FV0uP9ChTsWtJUKKaX9JGoeqvUakuRTUdFGJhiI8f/S6gqZ7Nhh12QimUCaRM
pwX04emiUXpxnM1c+JnBNEfNl39qY25h9iBP9cGBSSNulGsI9yu7Diz5VSjCpd/XcfyEfeE+QHjg
+Cqzi+NVcRbtOnEo6yhoTNTgiDZCLGWFzHPw75miIA9A6+xDEJCWMDgHBOloLec898wD8J552WxP
i4N47ClTaXSaueCd4kW2l2DwS2HvpSxPDA/p+tOf0NF9peLkXJsGRku4Yae+qcpkHfN+nM89pbWP
YsCQTBp/p8Z4NRZrMGu4SoYB9+9nsE6tdJ4gxedjg6d4rzbBJ0s4k6GIk65Wv/eyNJrSJyhGZhbw
lvVMvW3yKEaqff9svcpq9ZY+YGvLuw/tS42/pFt3sE3YMtpTmj98JwwNh4MGHo98XRzGFK7NusE7
EQAqGH7pSzZsyMP4NRs/YyfVAoFpAHYCaPfpnWBdgfUe8hDj71ZwvVQyINum7MGFXqSoBICp4Lu6
XKKTWDRgJaJ9ov+fKSK+551Y8SxPKIIB9BjKjoSk9uajQ5GvPUeGyU9mxXXp7AkRmy58qCFoREem
TDL2Hz3dtIS7WR+s5SXRuQUgU5mq00u5UfkDzk+U4k+ClVQ/ambDHFFaefcLcQmoY83T7NVPah9I
YyyPiGI5uO6DWKfvmWVHKNX/wcOgvCmmdLLvXie4TlLsDExI+fyWcNOssz+1+i89N1eLb3gbPDC4
6LRpdGB+dMxMnlC9qeYbikRqQZe0ONt5uNKaNcREWxBZ3RN9EP1/GwHhjXupGKAt6dI/vQPDnTQ9
W+ZerLlCO8Tt2HGLzD52Pb9kEKXj1Ek2jx68puOGKNfOaLw841f2/xnHxjVupifdsHu96vHArwm+
ryZ60zddcnk7NjHNGJ2wjMfoC5I4HRpUaVgiakKFD02JCXAYQLeu4YhkgfKk911iNy2FhWB/m27q
Pm2KuyZgvW8GIThJQPGYAPi10BiRO9VIkPgP2hPykEr77oFKOFyInsLsN0p64Khx2H0MlAfxE2fr
dGBHzt2T2mkjBx6oDO0C3BxEMEPU9enpcXluddyF5ITEOCUOYswhp6S24oZ9vRBwAsoQeGxiFF+N
drujuKxZlzzQDMdwcjT1FydGIOE7tWJMsaMk7KjnZPljmkfVJ/UHLfRGiYQDq6b4mm12W1tpfjlL
EFLi87GZGDG4y1ZE3lczuEJ0o35hoPeZw9sqKI0dBZRLi6Updxlo5B6A2UC3iqN6iX++D3Z96fdu
H4hHTMKscA3lT7UGeBSoM5lISgBs/5mKyCTBqRZgG5hpLglCH5Wo5SSYTlb9xWc9sZNsWQlah+Hj
5Tm8S3uik4yjwjo3ek/TkN6MDUOlDcVgPO++ZX42bTTCCcboKKLt1QImH5Zko/RrqUjrA6K+Yg+r
JxxmIMZELos/2wrDFL1GAlKZ0o6Bj1YrW8wbP3u+blwMMz++Tgiy0bmvJIwME64eFcXohP9OKmHD
7d9v5smnk9spsjx7OxkCrxsBwaRCRPWLZCngR7s/6ygRmvHprdW941ZZegsj/3qv3JOHwqS3ajCB
mmMi/PV7HR2WbiYVER9quBn7yisaT4GJFu24P1/jWf05YyoDZGx40Hj+H4as/L3hr15Gg0BjPDur
NtM6DiLeWtEbmeqGA19PqGMnOnobMzo22sITeKdsBl1SP+91SB/OhF8K6A7pvkEzB4eiQI5Wj7R/
97IazQDWumMTBRVIgJKFWmfBn22fDjHdest4G4O+vTu7QARZqY5OnMzyn0w+02MIol7Gz3O/FOxf
5nqQBEzzgnTDmrWIHL84y2YzlfcWiAmOVlgZIMi9ej4c9pn9qp+y2MrpfCoqY9RylcA7kZWohxOB
lz8IIU0Kn8bFrq9dP/B6m+Nqd+9tRL/yZ6mNWX/NWAYdao90n2LjomWcCmYVcXlDAL7GjhP89sVI
JRg5JR4Y65NjRrfolVCpbrqDJyUNU8eJIXHSZAmqPtxDKqXQ9/MrcgdXlzddNC395yW8yETi1p3v
mQ4SUop482HuqGRVkF/WcXLyxIPhIRaUTdIY4aTDlyOeKaVznwE6JbqAFUNDMvc2m04WLpMysn3X
cL+L8wZlQ/4nsNeLxv+bOzsCgeh08LyBIOa2DmrbbBm+iznxTmqGoYb/RKOc90b9X1EerFWo7fMo
QLPPUjGPVl0uZOXysEtZmRfjZFt0fj2vzvfAApGCsMmcOXy8zQOOX+0b/Eq1VJ3oXdNhdLgPdgEE
ZSxdSLHAodG3jGurwpCXiLe2O8/zKsJtLmErpYPleXYcxL+W27tYQ4M0sfAX1TMFQfCLpYacLAfD
SgZmRkNobLwkpMmJ8rp2H/1+q42p1MGeMcqt8q5c72tp+uNBVOK5e5kGfTDf9r5XyKlOWlMn/zXd
QhSuKDc8Pl1MSNVWmkUnCUaIC/ADGO0ggnG2WrX0l1WBtXemG4rbvEfF+utTxvCmZEg55XMJdVK+
1rpHNSm2yrYm3jkLDoysta+kiXq6r9GqnEGq82M5VtsgexEsqIdrLYLON4HTcl/nmfNleABYMjBo
U7e76o8UGnJxHqsPS7e37UZvkhcPLLFPqWWfdD6sFR/HSQz5g/Rp6PhHID1Sbd/9b9nSOCB2j4ef
/tlAJ7J0RX9B8Uve2Lkp5oo16u67/GUdcOUzir9vjvjYFRBFw5YcP5Us6CoDH8GPTThlWxMb+Sbl
v7OdxDPf4d7b8X8cKo0Hrw/fEE9P4nO6Rix5iXITaKvMurJz1T4VmFUJtVv2iirvl7SXCG/wM+wN
lpsWYdEIvtSfvRz+2V7tW4/LdLvrLJsLB4+orabpBUFdMUIdLFKpKd71SNvTY/dJ2+B+kjErED8E
vf8bE+NtQQYiL2aZ5Dwc1lP5nNylfTPgV3YKdAPv2ZZyZgpgO2hDdfDw9dO7XiirGzPw2LFAnGc1
KAGI0SvY+S2o1jElI8fTDyc26rad3R2zJ4XtP/cJHkWjHa5DETZdAOMMra+OtisTdZ4glpVHtGVU
j76xbkyCwisEwahAqOT1yKqtqxh7AuKhylOxRwMBOcBVDFExkL5xs2y6cGd20q5kIWJVMvLzcYoA
LUp3pVK7CErJ62vsdE0mmwEt271NeZ3cJd1RmxdQ/SuVsStH5uRAoHXATPLz8LcBiaWPTpukQakq
LA5pmGsn7Gw+qyC+dkutgnsn0VJOcO7IrdjK5QmtQ6BicQtqTNg5ew713PqopTNU9cqYC0k3NZCN
XPV5KPoZb9MdLDg8c272IW+zld5VKfB78z245Bz274zoUjm/MEgNAB8+3mZ0g3cMHzOe4oOwETct
xNzIiJvVVwzVUMcgUfnT72DnxcMcmtt/FGl2fM+r9+Gy7QQxoDc54x6SCGL4CEdHOS3J0zZqx8IM
baDrEgmQkj7NDsw9iGPZOb9aURrbfDaqSo7lhtVRWtqdRtgW4QFh0C4TBmkQOH4sajoEe1ge6dzp
bi9+/UEDwpTYO55cpsaYkhcVhFKmy1BiCQiAtnm1bs67JVWovOr9cMnGLi0AC9EnY2o+30VjLNzR
oSzwoISUlMXUhlMYwnLV41d/qX6dtxD7U5FSScbRwLUfePNGqjkhAuo70cWHUpGQHAJRmP9kdQsa
g/j7BSCB+Z2g/nFuFlRygBGYaRvZRu8jTcyd39g8+Us6D9mJQc7QNWCFHP/pxIP57utlhz9eZAoB
GM7ZWqdr1fgmimedHCK/N/c0lM2iTzKVBWRjQOaa/2Z9hv1RGthcGwmqgB3F1do64tzr26Ss7UXu
v5Hz6UwyefAIqXLtDP+PiOJNXvmPW/kZwwPg6dRRJyOEgVsQMWDri5daWsfiAMDHtXQQ84AA4DCs
pVjv+e7/VZ7ME5oEh+XTfO1AKvc1rcVmsKWbTNTZsqiNZuIuKatGWguZaOyCVvJs7xsqEYSyIVv8
jRssPG+lW6jTZHyYksfZeDn1elYcGF3KgK1qtFsgsEyTzeEm9SlOeL8zA8YWxSIFMcmOofVNZv4n
ghzcNdsNV0C0wFlUbZDU9iW/OZkjjgaxuHp8Y76++jgsHiG7zoBztWXvFa1RhcWOQ/8jcABdw+vM
vKdjUKJaZlpdBkgrOYG1lSSj3Ri/+UK4mz3Yp3fw2fJcmqU4ZCs5PwT610hBnNhEGW45839exb7n
0QQu3gymDAoZbVRkZBQzYRtOCoSMbZTKScOIx6YcV/b/EZOHWdFx2svTbVRGMRNO36WwRwRFUo1X
kVBMNX6c1BmXvKPZ/xzCVNLxVczZe43VCu0TpV4r+WrodWV07Rd8ujqGdMhZJpFaNyFzGaYpBu4h
qKiGKn5z2I4VeP1tIkmyiSZkV5mzP6QwCsWxvOSAaUYe70nqV+9MsXn+P+2EjJMawflUldR9Rlg2
v7YXnh9rtrDqwxb0aE38OUiF+zCCLco0FO6T9MTFVN5n4H1qV80WrGt4UC4vQ1Fj+AXc3cbf0KAh
ageZxVScaSK92YMaGNaQ579vGp2bGWglaJe9u0231ptxSSFBs7ox+VVvrHcYkPUPsHcRpya0ssj/
x9mWWA5rkgcw/IJQ4YdtnJ6sWKLILVDGcvEswCL6YPNm54CoEs/E9CN/HQl9+F/S1xZmrMza5aDW
FTdvnExUTr9Er1zgZSIsv8SnS8XCl+oOuDD4D8HKmsJYeied+cjt39nMLyzrDNuW7E4B1VEKmDp8
DfidKCPMKbTgrH3EelfZdyDSttZ3lTDULHBHXI3T44RrSggEFs/FvBH9JAc/+LfvDAWBY/mQiyT5
1Mt9uOcdx8tX0A4HQcmqPJPFiJ+j5698aM8xbpCZ8g8v+ZEE+AQlv5zjoKw1yjgqmxdZAqLyTPNU
jvfUkyw2AL5vnnom2SYsZK0dx651xKhs7voKbzwkpYNGmPYgo+OJiUlYWPVtrshJryeM/lMKMqFf
c1zo5LMGVnixq1E84Q7y1XrHsm/o3LbjKJPJ56E8rXL7eCz+HyYeafaGd1r6GDFGCYswKVdxMIja
Cff9zddsu6dOA70Soh4g/qOm1argQMuGNXpJO0gLvTbC3u+RMh2MBCQb6Go+J1jL4njO+VTGVxPo
rCGyhYKxcnF3KIZxqsZ7XqZzqtO6ciRWL0Y1kTmhPrk/LLXYFFNkI/zk2aD1wj6YjvhuJ9YR9sX7
f0Pyv/lkF8XAT2xZFKM3pUIK0w00buJkGdwo2NFqZNK72QW1Lh4mAX1s64qzSCkfJywO8jrzld8h
XxQ9s7maYszyCSDb4nOQVa++qc5wxggRsWfN6AsDNJD2xjV+TlJrgYrj4K6WyuUgV4bM5aCfPp27
3ZG4vb4/JRnJfQbFxk5DdUVXswMuEhXcZ+MpJOlMBC92hHDfwEM2YBpAB3juaFtw1wKmTNKSJUCJ
N9nNfl4cAAeSQ+aLxxRNuthYqeFx1zbpnP00gdLfHezqb8dHJ0MR7Bj4aGWFz+BnTv9fAgfdbXfB
efXb1m1sJpmrcsfrRoSSbyDhoR55tnqAHc+fV4g/YESIafCfjCwSsMRVa0ET95DCZ3onpJHoUBxO
YCFD4ofAB5RhGEs3071vYoENdr9OD9peWALukbiIpSvG/3Lp6e5eV+IlZQn4/9BVLKWMmQZFPzRG
0hPY5iJX46i/vplBf++812rGFVus7YAznTlhskFADUwfrzu5epq66Te+BX3zxxAFAaARDeeczwHd
JwNs8hjwS85CtiJyCCOIuT0U0ZL5IKl28uqP67obuWGJZ9eendgCQn77AaXfUZkEKHhcWtCgl1u/
1PYQ1xKlmLJT4u3k4WaeO7XjCFOvFKMphFrsPLYX94/f88KOtKeNmK9e1cs7mKe4CRpq2OoMMZS1
akTi/BOtKhztuEoMJxY4JvgbYJ9iKtovjsfIXnwK5ATkd1XUuOumQoiFPtap74qx6WP5fPqcy2c7
rSTxuyfAuIugMTKVvgoL3SiITHki+OvHGf9OxwWaL+PR6EnDCr9kIR3u6xi5dUJX0nDvlb9yOCOh
ZiFlPqSuWX3V4zWLg7pWo6s2GEEMTAN6ahkjNIH8VanGRKp7XsiT0HomxyU3qpJNRK8dHpa4gEGa
jt/hXwJmfbbT0jOf7tPc7FQGnF6es5yMbIlK7u+GEHT960zivMy3p0PqFkKateEs5xg3DJz71ZmI
VyzVtF0Re2DUI2MDExDavrhIwlAuBbLhzRLzUedFRM4RZgiGjhJhnmcMkYOsiOWmQMK17T7Fa4Wh
+UUKJ8WVIOopDd2oivcQXJbc0JdLNS4K6Dviip+vQdgXKSLbBkmR8n2ZpLLTGcar3Fg11J40yr9U
FjfW6MBqDJqhlWst5Pdunm5VEJkzl5inR5ZXN9gZDMpOhphzX4mqsTr4W8EWrkFweLNujmjJdBr6
nzt1hAo4TvcwKKsLO96z0zV8bNh5wpXDdjOUkkmZZIFNNweXNWQXbKZems2GdhkuEK8OXz7YaL9G
IeLZC2HqRaN0OqUuLffMBWKoT26tZAurtOccMqZyxdOjScZ5+SyaPKBrCDPFTQMN6iUeyj+XjrKB
+3v7rAmc0F7QKgqVgdN47dW7ULOfjKMHH/6ym1sz3f3zftvu++X0ASW8VKkHo8m/+o3YIGfRIDdW
QR8yUJzpVlmQGx/16i4bA4L8NoUyydtUX/7NygBfqLIR806McZHmSLL+WfpwcL+MQFTEp2kuVOQE
QS+ZbBLTrXDM+wMLWtptuRJkz40A+///5GSDTaAB8XA3hz9Ks8UJdmhsRMDVMW+I4gULUcKMteFn
KnctxzSBSCcXgAR3E4Xzl1/F7oa5c7kRk/S+y/hA5Wea6qCbfxqnbXdM0+ga1ak3O1kryaHSElbu
xHy/1iCTKzdSSrKfwI/lfBfVjlvvjAkvd07Scg1iTZp2VCYHgx2c+0Ye+jzgVx7TuWfCeXzhb5tr
ikUuhMAGQXmcFfr+Uazk8sQIBvZ6MWk2qksWRyxUg3WFg1pO15aSB7zRPlLyvcIsA9aOlG4DGvbk
ToBIGVJlgAjQMYhlXbYIQdjfKy50ftUSqGuf1joXpGKZCF86Jgx4fugqs3cdx2AV51cDkxOeNcUh
eyxr2VcxVjiPGCa2FRMB3vwbaxiCq6jzEuZn+ui4XdXfO5D3hyNWHs/7BUuCWj29J7SwsYqQrqsV
21TX/yMrbg6U93hbCpS5E4v78VDba1oKdbtgoFzyyEm2fe6RyzKOILDODbDFItHvda2/5K4EPx/z
H5eFu1v6MNjBX0SB/+KHRbCapRAmrI7VuIbN0XdT6wbVOjkRbqhjB3QfHcyYgcY1mqklhnGWrcKA
snBXvwnlyAfexfjYrm5Tp6l64JlCOl0/krYIEdqfk9UiDzjKUzNov88GTpCgSZqQtFXLepEpd+1W
JeGzoE4XdjtYz5+Vep+dLJa1pCHoGh0jPcEGRIXqRSBUBBgUGVyJlXfLRO9i31+LEdkh12p2ngo3
3P0ob1UjObcHDYSq7WAn1+W+/DXqDe5SJk4mV0biLBZdn/7bujp2kiC+CDPUJyHf1Vf1GwUy9T0a
yyoQKoYmT/0JkzWvLs6xR1sGUkEfR0GBGz8CfUhh5IuP6TnG/qk1O7p8Fr2OKsOoG8dO+3iaz2kk
bGipAxGKHp/X04HaAN9jUKp08mCOoTgakd6smw6FLqaKqV2j99BUP9hy6p5TMIo80K9oyBfz2jJi
zSghagajay9jBCmONyOuMmUBg7V41kunyKNrsgzqW1J6Jf3JIWpy7rmYd8NXQET8NP9Mk00dAxWF
y8djx0380Lhb2jrEAHUCX4tBnQ2ZHOL/RcVuCk7cDLr/S3+CHT5vNdcslCqzghSX/81P9WOJFyKz
wRWZdofiDgX1pj77+gjPfsCPD2x5vPtnFi0QhRIAzkYor7TeptYu/y/KrdKS3cFtxyZ3DPSgvw2D
xy71aLIUyiaC2fIq2/4YFyup4WzhhOy8XOh7FRjxCjcf7Xmlsxw/vUQ45nnF8/4Hhbdbe02rLVbt
cNDY+NNcAjHNXSNBDl0erNxIBD9OBE30aI3ud3Yh+S3slJAjAdd9jL2yx8SyGdwbZ5vd9N4zxaJI
aj+Aya0/AQGehOjllQG284K1Ub1E/38vj83utYPeMK8DQB9v2WyBRvI3gGqR/r1bhp85MeZGEJUN
afgcqlMGCzPEWUbb+lMBUU1RFiG4KR01i0pGam8j2Jr5vJWLnp5LTjhcLyGcQvNjrvnpJzVZbj9K
1T2c8pZA5l462arFMkjN5fLJCeQTHzQe+kSUD1XTJYBAsX+4ar3om1L/UCKq1cTK7JKCVIbJicVb
sbLe0O1OjviRRyPYGzC4cfVnagnw/Lxt1YccaX5hA6SksMjqRn8cnuGUkG+GC5E49tWbAK/76E3r
stDxb75tEyGH2m2OhA5adOFcsJMMWSbHWTryUyK1UCHmJOA1qeeSeYjrbRtWhTSSWw8vY653CXkB
Gs6SrPp6hgwF1y3+craZ8Bo6N/gJlHTTu9WzIx5viuRUY1bROqEEcrXrhlUcSO9YcUu9bc4XGJvw
30CaCfouMxCXMsLXRWX6KF8S42aIy/d3f4HBEfM/d1MKXctECE5rvNM/MHm7WWPnDoiqmiH8Qe3S
MtKh/wkDL749F2+MPuI1P2IeEBVrgS2sIYVDurhdakPSaD19k8+W0jbFPm+LpsrQgVXzmPbpKDdB
6ohjxLeoagEaBYza4uen5pV6LKlRvJIyKLZnkLh5P82PFdmdWQdjaZ/MV7vHUbvA4M+WTYPXNcrt
5ufn7QArNh3pvmVExlRiOZV1wSz6z0yHn18KT9mBFTiElroBql9hfQbZnVt4/W8LuRD4dhciqMyx
R7iqlTLuKASKC2x9ZgNPBPj5XE2aRua9VEashL308UyzT/Qq66pK2l1FGwyVRXaMllhPsHUMxNSf
Lsmild49ONrRzvQb3zoZboYSTbJDC2SVy/OqDxq1/8LzlZVoF8jd6qr2P8ieEnlimb/pP31vkTvC
GtMuPFUyRk9E+ux/IExBiEb4tfDQCSSEIYycjfZwmG2Oify7p2g/nUKjjeXm4l00y9g3jj73oRAC
wfnRr2V6ZKyKtmYCQIuTlRDV4m2MP+y8b86jvbOYwVeRGGapIlJLnTHQMGz3/h1zONRyIdBhx/t+
+cttdZYpgdOaWuuDvq0FvaiMoRyYU7nYRQ1QTCXibA3gxMNhxY9E6zH/d7Am/HrvbIfBwkCmU7f+
Vad4w9A48m1utMJPX8j12zS4+KctvwZwBFNcpx6ChGBWGSq0melfUHMHAFc5CoBkqM81JF/4nCWH
GKGxwVC2GWGG5JqSvQKnquKG7I/ZRN9yPl24NpRY93CKaX2Rdo5KYfJkxDoqp9qS+56HRHv0uUB+
53aQa0mXLlY56E14wNasW5tSESzASIlQn6k4DNQCABdn9jbkLIbr91jWjTydxJahJktev68UfkXj
FWqggHc8BQp4xOHF2LV4Qhkl7TrzTNMNkPc45fbpcBmcnhAbNLJAo6Qb8i/9c8jJrPfDIUjFpJfz
mLozKE5EUK53XzC48rYFRfLymKE4zld8srJTlA1QjNAT4bdxQxWc3+11MUQDvSla6Rip4qHl02Qi
Ow1/PBbk2OUE5YCC/ReksdLp0oNNrZfsFJPDmj5LVj9rWZBGWW81Gqjq/Rh+u9mvHxCg9K9zyw/Q
6dgYuRtrD0Q/TlgHsN9Y6qfxrUppNtqa/xshXw+at/IiaXxazzX/bQ3Is9SRoXo4SaH2JDEXVCTW
YhZGzaYMLkEfFKhw95MmMkIawOE2NH43Bh2xCVHknDr97gczYNeN0qONcdDraKf5jkcYrKSWCYfR
M20MeG9RLrGgbTbHa2dTQKjBVxK+8HHwiYT3yNYb9/l76TsNsngZKEcKApqGd9gRFjPefKWE8XuU
1lySaGeXe68B3QbYSTFNL2LuFhsQlCjfpMcZqdU+gKRqTKuRZ6HaZt/HTTaPekTMycaNuCD2xcww
WlUf5svfYP+owGt+uRTAxkbXdu2/cGhI5c4/EPeU6JqM/1Ksv43JhqhF62vdbRuYWgD5VUzd7Sja
9sKBMg2gl19UW/QGvyqmI1QJw1Dg3lWX+x0ylBbiZMvqS7Qlc+5DQ+DTCa0W4H7dBdr10ZcR4Wfo
ApSyOvMkwH+pYvgHJVPyxMt2/JOWQuw/UJ/VV0nx4QCZxed5I/Wn6Xd4IpXJLRvhNj/5eEMcJxIN
ygGKQdiWDxoG0E1xu8Nm1olcaxN8OdDIM98lS4U6l2ix/QRJlG/K8i8TP3MTNujY1n7xCePIxN/O
ugg8xnqiu0QijBTNwyeD3i0CL4iqidk08qlTsbOng9oJDrGJm8qPale0itDVf1bmTjIFZs/FCWfY
vCISaLcFoQtO/J/vTcHIRXm+KNa3EqFuuRtZ9JVoVtWYBKYMJdYHV1mezarGePa/Y62TpEz5OUBe
KHAJr8dqADo4FahZ3iTDdyG0+8oySezbYyUbiEElLwBeJb8LHdp5mcmaDO3DlH25fi9RxO7HDHrV
kJbd0NBu+y4tN/NIkpXWKuMLXGvG/ecCPCjJ649c0oFMms1KyKTWyd6oABu1bU4Uf05Q5ckwOeKj
wTLnYM0n6d+x5bNKHCQDd9sDKzmlsu+Rt1JbhUtuns0ov8mAr1hmX9FGzJSsucorsHfcYHwxJ4d2
nROX26FQmr1w0SkgUvptrByVdzwkhPnUz4y5i5kUN1Qv11lMiIznjwOh3XwpkXj8ge2LLvQqSMKn
Yn/Ix3bgvBuA7ATMgHkmimkhPRRwUxqIIgcg3km8iy/nzj3w2nx4WDrwDTUpzLd6Jk++y568SMkI
A1a324ADkvbyUBHSnrjjkJQC5sV6oaUfeM1DJKPUSJElxT0kcDuYfyN/NOdqRHwRbs7YfQ72LR2o
jM426TVrANMrOQ59ePvVKH5NpZJQ5FZFxS3FTfQLkyBg6PuXbNberP24cdZqm653AEPJFdmejuQ0
zwMn5U6LzW5tp4FJSKYcCQ1FoTtoLLRYdWnSBWcChzegeZo+0CZRSVZNUw35sa4kHENT/JMZ1aX7
m/72zaAAHY+8vnRImov5bQjXan1vjl2TrP8iHlKhqfNBj5qQ7iET85pS+K+0yCn0g9bwVTRVghHo
98pwMxQTBixmvfP2PMmX2LVk3NzICZkfGs2j6gjEnH/2bqUhGqD+2OldOaG4UbSzz3hyzWrSmUkr
qneYNOmxLN04hLKPy3Z44F+JhM2qCb/sd4rhVdj+Pg0QplLSLVhuxa7llucvjxMBCrN8T7qxYynv
uT2F/Df0AORNKnZtAqzfcv8Jy4RmO07uFvxuIxRrgUfv2MVavsPgMhafnTz6SYTne1aK2L7emzhw
CnXJ7ZahMrxo0tQCotNPVQ7IACOk8a+X330DjRYDxFeS9KisWKmF6qAIY2mA3bIiqBbDb7WJs+kD
WbniFmSE8KzPDlhkoYk2bukLT9E1LN7aRNqPCoqqcT4Tav73FaJMx7v1Gj3QqRLMUiNUY1F4u/o8
ODJ3KV+VQWyjzzqNU/RqfSy03qSjG8SwHSizRJ9sWn0i5Y3PZm6WWvi1twBeTHYAOWlgjDeOptP/
y7ZMXpLVWwORS/tFIDtLooHjcMvcMSRBUckJf8Q45EZhLUsIwPBmgQ77f9g/NDMY5NR3R+jSsBES
KrL/OEAHgZKPUHBohatq98m7g+3yZkebMXt4njMdSrep77kZnWKJsaCTDdcXgZ62W7k91A0iA2LX
yJERKVoGYWX6QxUUW3y7zSs9jpjv97F3x2w+bQGkyeS2N+0qoGjtV6tt5tUAGORe9D3TrCEx/n/F
JZ1XXKZpHj51X40KC7j2iz03QMJmw2yyOslZpdknj0pBradwZKEUdH01D1722QvH7rjAn+FQVk9J
5cDPq3p24BXZEJMkfv+GvHeRsAPpoYC9G5XnvxcjcHpsJM7cz7bxt7LfGOQldYiOe+Wa1ykboSQT
UVhHCia+O8JEY4aN04L5P9TsksUFB7uon5lZ7aURxwwDHhxqT2yyMLkFzPKNIAjN0MhE2DwOwzX4
JMOl5WcVZSvi/bsqk43+Haq9f2GjdunO5o1nl5xwWepn6lmTxaurX+fO8LpciafVzugvEzcTBGsk
ITonzd+91Mmb+7A62PqFBuod3aFdy0GE3Icc0L8InXpm9dekOwVsNrT6piulDptHpE53KEPfZfig
lQ2WUA2zChjYLFVkMx4sdjTvF7SAsWg8FrXPJgOMmYfc4N2O9+g5PONw+h3+SdS0sE/6s03bnZDJ
Pz6OAASWjHoD6KoGIn4aDQhmy9sbaeG9iC82B5Ju9CymVE8NZrAQZuRPSOuxNX+RrN9SquQzNGuV
77ZGZuhjjs7/zxxteAIZTqZUbry+nheG0ulpXQEeQSNHuvSQ50YU2BDC64+reLCnq/D33tY3xCUd
CNrI7zrErJN73bpLn4S/1dU4ZEQlq3NjlG/lEXXdS9NPP3tUGRJo3UCl8QJ6iVyCcPjF64eeeoSE
WcI611UCMMFBrtlFB0YKfUhRHJG84bWytRNNqDp21aLBfQskZB2C6zpobWz21ifq5FlXyyUgUZJp
eFs5kYF8J8rSss7Qw9QRccLML7lreKNYmLKkB4GW7YpWFUWnsVBN1sN4epyZgcjoSJhmRIS58RHd
7TZb45YD0CAe9EYcWt35YUGdnBHwC/a/p6tgwavGxTLesVI1f8Q9WR2zqoy1WkMBz+wcitzxY296
hNhTJWfigSDqnF5JoOHQmKWloNEH8Io9D7dy4jbp7Zpu6dm1TbQAUI0ns0nWprNe3PIlCYYNO+9l
N+2UQeGu2kaAqZMnElh9tEDwuBpg5C2aTujcqXfg20OpWdrsk6iQ1iPnz5/2eYrQDXRTsE+9FCbn
j1erIxX3JpWeNJ1vaARFzov3kJZ8Qkkol+gSGb/mSLznTWCitiNMMnogh0DqL+2pGiggo/Roasf6
TarlqR8WQtCjqGcF8odKlx/w29oEfEJsbwrNghTw6f/T+0J6OVCGGoxEZRSnxZtiVK1xs6xiIVK4
5/5sgKfn2Yj46tURxGlJVsZJUUL4HGZx5ifXZNqazTfR3BD9KnCjIy2LMgsnhRgUF1ZpN2fB4Z8N
DRt99M0+XXQN6F5SASb1ZB9me3MvKSwl/GN9Mf6KWVtHunMgtt+RRmfPJxL0nT8wnkm5+gT7RZ60
7AnLbpLK9RQfCb8lDi5/Q4LA5NRI3CxvXs3i8apGMnSc/2sft4YLkVPRaANdKbzyXqW0uPoWZF/y
0DpQmpiJRUkd+ZFUlACcJP7wBNYhT+PBetVBAE9APS9c6cAymXi4h1c9Cw1x1dceBTkoqGszPXup
0DpUEiNFe+xPuQ9K1pH7w7SwU+pScIfwvBDXl8vii9B5k+MTfxKt1e/wcpnrv6LA0GOTbwb9oUBt
tQWS/ocbMEiiOnr7XxpBYzfAsqjE1FZipdIJp4GiA0rps3N9TjGk7vTK8Vq2huGB5x44BNcXWTix
jidz2RIzBZoqrjC9FRvuCFgMBEgXTCS+Y5Tt7doq9WVGvQBwyjY3jirFgG+UWaNlvuOLTtCaYYUO
nzte0DHyInuQ4oWIFlpK2iBl7AY2FDKTshht8TyuAyzXU1bRi5jBJvbgf8zd/vQvM5CbBfljlxg9
Pav+94lbARrubGI4iJfVxSmXkr35fIJTF/AK9hM4VnKMRn4Qo36fpHjPeJD6axeQcJ9QKnQDqOTh
32t2wTPNlE1/q0cUO6NQnE3JUEBYe1Hd2NE9Mpmc+JM6MUlDLmdRCiH39a9871pJFoNthr16QLHJ
r2ahGNnrEx19Q2oG6yiWInwk6+0EHZQC84x65WkQtYYWHArbR/9vRnKJms6UkIhJoZDu0yskusqq
9BmqYmIJgJXC5mq+v4zaoZLiYlRHWEd09FR8iwS6YmV+kkFTawMy/lTI4dkyJZ7oWJNwE34lzny0
j5wfPImKMhM5dfHyskhFRlOcVGmNJKlNio2OQVmdgGt95AMc79Mpxxrwyg11fM49VlklhOSmcnVi
fYJJdrQxhO6Y259U0Qe8TKKxfFMG19bREjLw3CP93QTrXgjEyixqiKrCwc1wxi5aIPYW0+w1ZWey
z/ZqNGNb9Rwrr0CWcIx614RN/UW7RFUEj9MFWBpvpn63KDSEGnFOsQrP6YM28QG14iGuu/5NU5f2
DORJwZxJ4B06FPzExLh1IAjqJszT7ct+yoezUdB22BpkRcjhojEQVRgaKAJol8yDPPg5WXgB3GRa
tFpKkkNsiwo7ZG+B0HzLTH/5OUxkIRz134zJNL89wlwYHKu5JhfKyQc11DKXW1IhRQRdwtH4sB6J
w+m1Q5w9V3zXkPxPZniGxj5rchsqnvhU+8xqRalvFFbrAjspvo1IZbal2zW7ykA/xKrRaDrNIvMD
X8WzSmeTxwS31eR714phSx7kiqK/rL4F3zrCW3gHzrdhZIU298/rHJA+lmRWxbEo1/o3BispiGNV
BGxUV8zFG2miACkm24qesHac0kpXKlQjwr/d8VnLKrvk2IXsOl0wRk2k9Ef9yZ8wN4C7pLI+iS+e
A2yqs6BOjYR/BQYDgVfw+IIRHj8vc6tjwBy2pKLJBSbmwcwWuavkpBgDoygcPVH4Kn5Cso7B2PyK
j2c4EN6iL9etjagzn4XC4461pKhoUuF/UHtoOP7kK/G6V9l4fi8Cw1sgMjYId0iDDvR26tAjD64q
VwzwYB+cAnX1uOXqAwFLlflABzzxWvZFD0CyuO7ta9dXN5HBzDVbGDNEHhX6VfjwTBEZv+1Nvg/5
FZYq7z3OsYvwmU5RpO46a05YkyfXkl9w6unjm0RcFihV1p+q5VdMW0MlaT+heH9cCEwaKBz9Bn2b
fDTCTFhaklG27fVLldMMKv49jk+octdgxC7LoSNpIClS9MZfnrB5sCiYsfFi1l4yo1O6DjXJIJnh
EOWLnONX0YJ5mS1OQFWhEhI0f8U5z7twIJwNZt2wW/I3yAgB01UksNq1U0jmLG5W6Netc96e5ZJZ
b64/ZHcwAlx7IA+Aw0a1IhLU29h/xnXazI2KoA4XbwD/aWfm+HSmiMSrvWUHn9GN1JwMhpOwL7yz
FZJgOdwjrE+y8+GxwzRLB9HJTvc3HDiotpuG6XcILgnNBtbzULsPCc+f8ivY6JLiFe/CVfpb+gU5
2eT2rWyq3d8NZ1SBNc6Ya7iS0ls3ENQU5EDTEjHNe2r8cK4naFTcrkGF+hqhLvwIK3klydEpDpU+
ZLRuRLKze+k6FFvclYcR/WIpkbIr6Ut0tR0AMTqUvL0uWQy8H2G4FOdKW4ptZAwFfvKuII6qT224
sBznIim/kiL65x1KkYg+IZ9pY5cR8lFkeIwYkkxJyudPWJdGncUIai14AP+H8bq/e5X5iCZUQX75
CEjaslVaxWHzT+mlsvLXlB7JBelTnVINon2DedQ/9JkR8TC2RMwcQ503Eg9IteI8G32qj7NtwlL+
u6X7qC7H/rubhmaFbmf8ntV7ny/C2yhbq0X2+UCk2Gh1l0GFrOY90MRHK9EeHj2WtUl9jQZgpPBm
imG2r6aA47HcwGER2EA2QYQd52Ocx8S4PnJhiBjNk1Jli6CEy2CJTE8OouGPgzz+u8SPnsuAvH8J
uxXWPVWOunReklEGRiSyfZZbLwg26dv6NHfnGKd2Mv6m9Y06gCsFo1ALRK9iZrtJ9u1T10gJ3cej
NIG1nn9Bc0UAIXAYakzize5uA61wVfMWCANgaaDzAfWayQBB20K2W3uYZdMokgmR727ZTRGoNNTe
c4sGMeBDuBmGIcHF2gMKurSJK1HclJoslZQRzL/riT9NMtugmYo9dV2YIlPdGXAJJr9c9ibj9YPc
F7DuW2ykUgS5mBKSXt5Wv7zhqi/PhmLEoDdiZW8lRkvHMb4+yZq4yGtFvr3nnqGhbcGYPIIKP8aI
/Qy6J/jdnkmSfZJcTZjfZBUwjuiFKYYeRw5mCUkXBD/pWW5T7c+gleGhKl+rnDOAmGFVGAEdIpKp
Q9LB08QWehMIdaAPsa/OZmIPmq+8FCxIYFgbr5JPZRjg3M2k3ZgVT+UzRGWuqOAl1HDMKmrzZr8a
vD5ad4d/NDP1nUfYuIwSGt2s5goAcdnq69m880ZVuZLPOM+iNw9kMry1lnGMNNgLmiisPfhDfQFe
Bb8tnbM3nLjuvwE57Bo/bxmjy2BbkacPHM18s41ggw5/ebWqAiXWUK1JHz1HF4xmi/rtNeCeCRgl
GcteNQBmGPKnndpYX+HgfJLqmHwyjR2bB0L4sR2MPXjz231NmWu3HLdJqS7svhXs7Ygj/BDTdVsh
uuaxsTSrS0K/RwFUWuBpjkVIqSHwjvXORYeT6EU4aA4ojS6fxrsCVmyn94r8cg/D2LBPBxnFQW9Z
L8Hx2UDmAHJECBmXHT4QkixTHqi3tdY8Z3CGr8YS6+rleXIKwG4GMo9Ps+S+XxwnUP4McTcNTRUE
XLaPYggwDjEpiGyp+w54Nh+0RHQIm6ZuHwP7UfqhvF740h5CXFDazc7JvkpXa0CP9H/KY8oPNqHj
WKY/QwVGvKI1b6sRG2TSzYPiQQMNi14UGr+jsIsHJzMsBDgZP7BAdPCT/s6u47sbdD8tT/U9fPTq
vPgMQDyFVs5otolUTsXoyuFxStqHDA+bv9nrnHqckT1iQ5MJo4VFuVS/fh/2BRJ1El7oD9SAPYri
lR6qFVK4SBf5fWN7gun86IM5xrI3Exiy14PK5KJnm+8Q7gVqno1ZMcUPTCBgxQNCyMHqF7oNhPe/
49LmTWcXqnCDWcIjuqZIX0CPcGwz0c0S7f2ATQd+/By0mR1vjC6sh9scfzTwRhEPDxOo0ZDheEpr
BlPuZKnPngkCY0o+75HxVsUq24zWmoMd4D+YzzYPrlNxbMUxIvkVHZTh8lODPnk/gzX4/wD2Dgyq
tKo7TmgZxK0Cnt8Rfeafajc2EgoyJlj9MunQ3VQkI5JCQuZ7xWKz3dTY7gIWXvCUOQNMayZJJcZl
TR/YMYd7dEFo1pc/YOcUVKAC2sPhDFHHxzK3nwjCXK15FiY3XHbG+UoaCA9HKWetT84HW2BYFxux
zULpsYk952vrlrrWjo6TxWM2guZWJL1iB55dUgpjN09lFciwH3FZ79omXr51ABj1IQsgs3MCsyyM
mCuiuBMJURTWaPLGExXbirP5vvM3Ya2gukX2rGZVa93/Da/e6KjYsxOHZ2Adsr0jYLINMxEP1wTU
5QnZp+oZcxghYaWXPn9IFkwUQmoJST1RMvSaGzKsl+0ju//pxR5vUgu9wWDqaRYqWQC/OA4hqyvs
xX1T5fjWV7wWPstB90L31zBFGbI/tfkjkNQhGXFOv+4H25SJdLSy6+d26MjATt4pjlcYXZFca96X
XqTol/ZLedCtMQK4h5arnQXZjMYgXMXsV+XXhOFUMowT98LwKj1LXicBYyCzRb+Pn3E0hqG46hAu
cIEgTzjFGt4JpCymQnw31KxgAcNKjIpMQvQmwg4Hw05SprgyWia1KCR7+go47d2kc1oDHP+iqyF+
DzuGGlnULbG2jmuw2eQxCV29ZJDeFnplz7WumUswwAxMw+To60vJ5vW1d75Su5hFlgJB8haX95oF
744RfGfzkLV2SAFOR2h5e1wMpoW9E6JNhbjk0H8SLACda2auZrywNSB57bNK/WjTnvdMDVqtXLj+
6c6yqhyfDOnVZkqZdzMP0si4KW2tTGq+wuyBcG4imov00HDemLP5Xpyum7nC4gA71Pvz/Das8jS/
JPN3cZwwc9D1k/Y+3I4yMsODnIOFeiKanfmAGSByYFWS/dBHQpJO2xhTx3sj62+0PisOFjJXheKj
dXict6EebpdTGgkCyU9PMq/D7dj0N1ZcMGdYxgqF9BFX6r4Gnh1q3ogIyiVRWdvGzgfZmOWVtJ7d
lhNvZR+65RU4wVXFXWGKXZYxJ5NwRdqM40ONTyxDvESDIvT22KYT8iE9SErzBD00IrrpjsmaVNn3
MV5LuPFfDuGjfHbkkmnkHN5attYNqMk7gAH6DxHyY2NXzNhI4jAeI5v/v72IhlO16/dVY7QYRFQZ
izgZUdpznVEyyz/90FELOnbmDlAr24kkohUb7iCaBKGEkWnGUDZ0jqaazgYQEw4GFpHu9skfuhue
vLTl2zKgM4kTZeqHjbpavjA1oK4vbQ1CxhhlN1d4SBNUEhbKEGbY30IF0lx/+TuhuVsT8I4kOMDu
fRUZwl4LMC/14s4AGQkYxXViMcUAEbAnpb8tAN3vRHCY0dVaXKBjCcFJALLzd6ng6TyYyR1XQKTi
cOM6H4WZSNA5tysaw3IO+29y41AXevulYzNqXygkv3oCykd9KPXgjjssSCMptxux7uo5Hag3U9HN
383E3deh/9Eo1PBp/XlNMHpOsCT57qJfipVsYOojGSwJotTKxXBllPHDvjVLp+Wk2s+FaayWLrxi
lQ55e9xDiDdUPbkahGdG3lKEmXpBvCWl9jTsMXlEC6kFJjEVp58nzTBO/q4LjvYAPtVgQ0WH2UVM
o0OEiNAqWymlFRAkeIRcdPGjToRKolXVN5igiUzX9lG77Abj/H3/0YnwGdVr/fP1PjT2NfOKIjkc
lp0HXaGkGJyhOhXc8nmlq3ZzwthsfCahHE//t997jRPMB1NZ9C+3XiT5VtpFnOwBQZXnVtICwh3P
gCcYuC3P5ZNHXLkp36ctisYLTiOgBCRXcLyzdSbiVwyn8gN6C3CmVt28+dAM8U6QB+bBO3TkIlli
qZhx5RomtyLScMqPbWTpeppqC4EP06w/diLWoj0oeyUoZNb/iewhWvdIA5Z7Do/I2jzYooXKQw5a
ehW51YpPUvn0LJPs5lgp/rVKxF73MVg0bLrN12HhFxvVhR9xt5JE5OsYqP54UsHZLaqzorRCyoFd
VGXmDsrCoyHNRksICSrdmo0jv9eK2TopmSiSf7YyqHby8z+dTt4ztIEOdxWb2ghZXf9ImZWAIoZs
6BFURlPaI3N3XwQv+b5xNv2E4m9wVH0nGVSoVeLF2A2sn3CGvdaoRfcxXZ6DN8llmQhJ7k1aDigm
OfkNQRH2KWXVicPVPO3kAb7yeHop4KoShPh3AYxNH6OdA597o/6MsOtL1FZyO0VS0B2apAgf9a35
NUVMm3uSN7xw4XzZPIHkipQdmDClGxib9NwKLB2RtxTP6FuUrzulefcwUhcNrMimMjfUHx6ignrX
7IZqqx0Y9sgfMNkbY3iLIZxHhbwrwrPHgVf1Xpn4lUeFJckWC1qkBCnRocpw/jU3wWgDlPb1OVkd
PK6QooxIvgC0b6uyo3fdjBnr+KZh6497RN7lqgcTsL/1zYoPN5EzBYh5uNnh+sHgb109t0buPApf
q3AskOrq8kmZNA/LtAdD17s6bh2hM3IWnR/PCYs/tm8kPOvbMK3bOpOTTjO0dL5ZgZnV/lewJ7/p
ttwQzhTTeZeQjeP4151DkcXGFZKMzbMoT5NasycLpXhzzCsoF1darVrJs9nCaoOShTVndbjGWfyH
/2T5Hc31iwtbaXdftC1IFb8SeYlHhnGztC08eAL18ytTqeFg08EM9uHN/b9h3PJ3ZwhkGXFFfre4
BDiM1Mvd3tLrqNs7iXG4+F18eJTqmbNkMEjdfj7YZ+txud9dJGp7+T3S5HYkQ7gmyREb1pR0AEKM
e5AzGfGXbHmscOo2bsnoZRmJ7LlXmkQoAN3onU/kJVlzN19jrhpoLV3q1YukArP2leZHU0lefgxT
GY6IQJPQOrRUuBkZqDhG4eo6PDIdydu2GDjJ556PXos+XdY9rZq25q5GMc/SKBMVAj3apTvWfi28
7vz76vioPASsmiECUnO3RjSE2iFcjqNcbV0Vc/LgdPDT8o0cfq9pb/NgXw17utMYk0ZrpYmcwe7Y
rS4LJ3/AC+5EI7f141TMZlulrlqG6tzEGE/CifawxnJh3csh0PoZYKH5wEiQ3yC85xoLXCvevgAj
WkdJxoqGjXUkbFltLvBVPPBrOfTRPdNNmnT0j6X4jAf+Dl6r9b4LAlZRGDTuft/ntJhEjXo3Eoy1
qsNwFv7mNyqoSIrYb00yRhZAa7e8K89nsdPHqBdPJ2FwCdnlp+7iIg+cgD3bJ9mX6WLCbNFrjsiz
ouxrttuAcMGxAqSrr2QhNsPEa5lURvN1oEHIZDQYatU/aHuJYXbeqYwWwyTnV8DsE/t4+KvrBfTn
1HrwSma8V+0bT0l3o8ZzPOawxTT08SPfa3OH+RB1C0D2YAQNYiDY1jlxXcCHUftvaBsunVKoZfOh
4S92dugG/ChBznc1fUtKnt0Zkthh9TqGEn2SAjd4wVIg6MDv7DuulYhi0iVkLlMvAf+/Svf3XqAR
tKFykJXOUoPTjR0ayUI+8CJ3LGXWjQn59XKPO2A9rXAGcRjEJ41j2fYpEkbuDnNz4G4a7RRe6Mna
42Z8977p2JEGbMh5D3il4aQ7wPp959rqT/03TAxwEkLICSAGU7aFXfASoQ7lOKprm64p+qWrGpGs
i1D+RxNXgmryOIi4gGqysr2hQwm2JdSqpVGGBbMaRmvWVPExySk+ZCZcFOwnJ+sRVPO0Vx1EQ5TA
Kdkh9L7mkkMP0d//Tu1dVwhj9ZXT5+gdGeb8xe67w36zBJOI4b4RkgEO8osnIGKmN4P+1GfQgdA3
Br4lgaKh7fkV/Il+qxY5kKAwz4zo0OzaumjJOGBMthQWyhe0LzRsqVrkYsPD8kHINp0DCKgcy+9/
7apcnSH9KycqryxDNCulnF+mnsfY0M7k6ZJmyNSmntLbWWkLwxGpeZMHa5zm+1O68Pak5xaNvncO
EeuSHnCiLutxqgLSBDV/7BcJK9xgW0qb/GUsPembx1xPUBb8MHKRgVkxtAnlYuDdm+Fu2/PidDlT
ULU/YNbZTYvZ3tvpqcMUTOuXxi1MdIXGyJB/Tai+tKEiQWVdP5sLlX9uUNvrNjXI2yKn7+zeznkN
3zRbTo9vaOg/07ra137Mrd+3FIZ9qjDGJpRxnV+QyowrSLrrY/F64q9nKXzl6IanVUKV2iiT6TM+
avyucZ93RCx42SvnMWFy1ZC1Jqpd02GGe9UtPku/yKn1F2ceMP4lDfZ+IBzfopsrPGIweEAtjuoj
AiooPrplDpRsHYp1euV+XRNF7VBJ/reTtefzKykRO2O06S24beh93vyFtUPz6nbMWzp6MDeaPVnK
aB21TiOKDEmFvC3FGwY+mOSeN/wtT+cVFd8I0YF+Otg/oisvvBIs4jOBVwrZG7NKTE7aXLHbgKn0
2hDt40SoeArY8AymOWrBQ0QY+3znCyTONqtaE+C+2zU4EisuFkPkgqXi1b2Wu6dvo9XZS0sObpZp
TyaTf/im8H9zslgrAS5FFCJEvIjcjv1AWdKMhOX3OeCv0dgHrcf4NKmPDHE3Mew2LcQ9QlAKBC3E
FpPRbPaP29Lif+CtSe05JKuR5nVyzrqvngTBdzZb5D4u2uA25qjVIxofUA6yHyVajvimwVwlnvRI
jtyN6xFTc4le3UIoh9sjQEKWb8lnKmNz7U0MeIlKIppMQTGy5OJPiD2p3ssqgVOWe2GMEQ06ISiB
QhM6fi+2hM5BTo7B5bpWKE6+t5eaaYO8vGn8zDaFgy/2aR3Tber3JZTseyxdfVSLTZeP2zYFuvdC
A4PJogrtwuj8wzSnrs2pnYDT/xdhjL5/LKwLlEkr82N7w3y8hj9Q9kyN+a3pzuXQcPClGAmY8c/z
BEjUW8N8qyCP8qKFxIYC5yGyJdPSwuxtPU1+DUl2R9AL+uG9uVW9CJwKtUVba+QGriLEI2F8+rVC
SosboiK0XVvtRC+Hj1b6iPgULrAoS5mvQxsZlqbm08pNOAFQpgSlzFDqehsAbXc+DCvVB+CzNeP/
smh60Vv0SKwYroNSL9TPoxJhM51enb0mIFqCYEuidkqbKhjv8QWMz1iCpsjQzcZ3U9xrY+91UEVb
IZ8rBQN3Y0fgPNRdeg+E2gMDuOScdSL70NgT5+bDftOyvhtxLSeav3xcA5hekPqAHkmKoaz2q+G6
r928exOu1CZQzZA1GCYFe6F0it55JnpkzUwLhbXn2BZcej6yNm4mlvESlJE2/NN9sYp/oGJ46f67
f3nncnnLVY+KnscB98UISlnO67lXdqhLZpWUu2UNtHvG1Ih4MbLakhYwBWi78V0NzNyLq8FlmYTu
ejWtYycWHozTOXdtdRcXd9iD/Hj4SfZ+LCM2crXq7aaOT9b8RrbbRlJPkWHSfPhMXMiMH8Jm5hh1
cZbcdPJAw0/WlxEsMfKCPodIONTIthOLTAVBg/CcmKSEXud037trWoYusohY1Ru51jaeQhIMqLKo
5476LAA6922JB9dSxBuvKM5fc3cDQRoOdxnhxvIg3qj+4M3IjPmXV7mRVkO0SRw6T2zQFA00z5Uk
LUJj57u3yuzbcnwCih5aaPx3F+lYUtIaGhmgj3eI+geD3z+g1trQaIDNPvjHusUDXNVxzcfgtFbR
nZY5vRbWjIVpzynoAXYx6sIBVxP2u88SVPaWM4oyyJCY9gttnS8WvKEgGWfYvG6XZcXgGguYegTN
vQyCqsg4VSetjN6W4ZP6/qr2TDa8+f0sc53uWXKCn9WlEoRd0mSMaMps4wWkpjo0Fpd5AYPtA8ft
93Bq5RCG0nXzAoNzJ/SDRzg4wLIESh1TvxmEMwZ26QLzUm/OS9M7MzWw7j6xS/vqFiKBDUb1V/Wm
xtR7Ko52gRNJvvlZYZ6yj4Z1MtBFiiWCT8v3MHeQYRRudAtPgPWU/dEvqQwMlOTk+vjkoJDOn+F7
31iCIqxdSVCWjunINkiYIH56pvrr3T2CEU7SXmoIGqTRkI1wXBmIsDS+1MTp5H7Byxy4J6Yyhbh6
FdVCnJRAKAZtUNmKetFAOmxYKyEY80W55ovXb7xTx9L/N7zMn3P3XGrcM4Kmr7PY5v7W6gi56YME
3FrXu0flLPkltT2Vk1GClME+Qo6Pe/nD+IY+Jxu8ux/o7vG87sO26HUjOF+46S/U2kRyhEsoeaYN
98nqmi5t7hTNQS35C7liL74N9gfIBK3QxHhTMKfpvOZOfsT+bI7BGWYEpNLwhVoC8xEpstrLVrv9
yT0pvOcS+i1tGITSl2oPgcA+w2OFMFHf5+tMif6GqZFErO9XrrWRryUZAv1P9pHRW5zhyXj/1T7i
FR01+JENJkMqY/0R2zIGqciG9nITw3OfnIBGcdUgTFd5HTnvbCj8tRlwMEXSWDy4FssFjo7hc4o4
kjtPuaeeSx9DXDgSUQZCuBaQjM4j13wyslkOOvyYhUNE32CMH9vyGMq7KLD8R6ewxd4XeUibKSAH
XDtZI9WHpGw8ig+CqhY9JrGjFwX2MM+lZW8gNY1halzW3aFg8PjfUZyUvWz126LSaekBXf2HbJ32
cdyg6hNvJTxGKL+XLFOpZd1IfLsvdh3qmidniw5DUC0GT91+KKy6Cz9+GKskfbXQ9zEoikhCIQ5o
MDA5KASeo6nc5srhIuLRHKPgqeGlB8YvU4A4w/a5MCtwoLhYpjkndcNpMu211MnmJ9X4GSEbejZn
b2uBBnXgeio6v5PcZay99K0YbWdspSwdAIquPrqsm0CvMsavx1ChLRzvSV5CutxJLky5N2mdfGhK
TMwMKMcOkacu22F0yUW7q+eCyzOc3LwcD9sb3c7QjLYLqVC6/QdMcaS2gJrB7X5p0nQ2pTGjkRWf
huXCWwM/rXbEu0+QwRlQl1BHd9u7wm6EOBtUjK2tGPD2/2SbZBJeaLuTdY6S+mQY3EKIUUKpJ/YQ
xEsaV8vI23hTtWALHykxbue9ahA7egMLfaNuI3j3100aH5pspqSi+l5cEWI6QJRApmDMEjPjDvQj
vG3W3R17F/DJKMUrFPox8gYO11Da+uiG9YSCshQYZfUvGvW+MBal1GVsPNRkch3Yfjo2taymsDjz
WjPvOvNjiA5KhXKx/baVL4U2xFHaDzq9YtG7SK58axk8TZ95ze9kBLzfYXdnJqPW/d41KcVFpNNp
4O9wWv1OXqxJLxUKMQ/vivVzXObM36ka6tJBQfI8+f2PUtsx4LVnh8mPJVk3LYV7b8On+GzfShdl
0CYTIzy5Ps+OZiQMUI845wdJEu922GnAeMQaam3mpwyjFEwubJzKDp4ExirdY8rvKTc4+5TDiI0s
3S7AwBCKtgZj5vWj78qV34G8NdEOAu8/Qzrf+pn3d665PpTKu+GwudL8MueHCvcswrOgoInGiQKD
wvWv2KH9jqvLZP2wNZwePCwJkeyDBapG74H1VUsWRUejWNx3VkabcTdhu1YuphhwAtwGqIds6GA0
Ai2mdEbqxDVFQufUEXueYHP/JoUukJvJQS85Qyai/mhf4yRmVUFU9HpR9LX5l8p6DA4InTTwde6J
SuL7iCOVXE7sfdO1FNC2krh6uiLovfziJBzhdrCyvvvTKSBBUdquSCuvMljbHxDFOFp5GJ/MnYgb
h06ZxmtTnIhV6nEXdG2zrh2aCOmAzsP20b3iDgeU8ZxXj6yuR4hPOh+y1ZgBlFEP1wL/7b11DZ1K
SQwGYKLDwwvL07n+N3Ma/ySQVnfrZFwbPFJXJkHdqsDYaRpymzsZVMWp6EFUnJ7Cvprak8et4gM5
+GNi5UNSVrgJLWyILqiC7/27qa+5vQBHHv6G9pRcroxTv+PWSPyAw+y4pf/tjaH+SQJerFkdEM21
+Vue1t/iW6PrnjxQwotFxksNzM3rt+ZiXnw9wzoDAU3UP8rZpCenTNT4oEeSK9xN2aJQnq7CHco+
IYz38oY/l+2rlTeXMP8PfsrdEXPghsbYQsr6hR9rWduWxf5CAkH1nUM0lqwpUTJXNYI0OoZMlBc4
b855ZnDidENm+nEjbLtbqden2CCLkrk8FpA1l4Kz3S6qhMp4+wAGRH/G3wSj1fn+sHCJt+oZD7OG
mqa62jzsPrYGiVsopsUVvvFcOWd9VxnmJUabKui85ZQo07ekLYuaVYxJB60KvJVRUC3UJlORHpYQ
eho816GwZVs+Mox21ENXThNib7m5V4oP/+KZ5EFN9aTrHhVO7zVvlgB+rR6NcPY18I9DGV29WdF9
292HcoxxFphMUEOnX4buzvSxGru4/waQjeJ+XjBNXLl9IeEcbC9NrkHO0UIjV++gkMYHBewN7IRv
nc4OjpLQzlLijX6+27oHgWNS5uY/PIZt68oW9dcYoYmMCpoTMpcRs6d+iibTnjE861R2/t52Yov4
Rqwwv2PxknkHRuOnYSAf/AxTJT666FpDPdsEbSZLUPWoxnHH8UWXpT7vNJMSeueuDqW4Yz19cdh1
tOuE1OY0y3YuMYiqRpjN1mGDJhIHjSRc7qiK957RZZoa8ASizgdDal/BRkJmYQ9cZIM09GboMJgq
bUWk0W44R8zvOaff8R1tGiMG7b6mBkaps+VA3gjsNuO6mOSe+UzWIsI1/HpPDSYX/7eMR+/l66Xf
zUAKF9ocA3ETYwu951JLSK6UMAoLRav0Y32dq4aJ2hFIzDmQNycusYZPha4D2JMx0eFtPW8igWul
8GrdQS2igcgUTeDdj8Bd402I6yBI1YVZmYEWafYszB4E+LI7YsPOGYuFOc7DQHx/dXJg0DUzLp7c
27ay+ogiTjAsKhPDVzmX3uK22TjA6dFvXbMFC1t3woJbyCIsSRZpTMXEu1mpx8XfOuLEKHhek+CM
WmQO4CADQuxREy7pYJCTT6D7H2U3wqs9V4dU+IcOhQwu4GGYtTOCGDMuWdgiFNLFiRYD5PZTWedE
X5XvtilItmGAVDL8KuO1EXDkNYVCGqHewWN3s4KQLFh512XPCTO4PrmoN/IjC0ELq/jwpVU0/FIW
bi48lNGSztpQ24ipAEn/eWdeZ+zHVx55oQTiv4zG2BR8Qs1DQc1RA68HJ9pCK7s+8T0gkfVOQaAT
vSF1AUGIrZk+l/wMOYcqcm4QAlcCzS7QpaKB8ro/doP1dfco0L1D64oDUaARKkFwTdujoRMBSnH2
agk2pmmKBuZANIVgDEMlM+n8LNC1cC+SEVz3hRC1zHyHGGYXgpsGTX9fFzVRoNY5Xi3WbN1EkICt
R/bi++Sq2gJDJa1IQOwln/hlZgusqEjWjIieOnme2PPZoa5w1dVwTep6fsFty558t5gFE9shL2d7
M5Kqk3BWEKRX7w1bHUFwC2I8XpdZIMN7J4XU6ahIYRwMLL28MmEy07D9War8gkxwi1rWMjN05yBW
OgoXBtqVZ2TsZZ0KKeJm4zRaGdt7RnMkA37377WIGJquEOXyOfooJJti9jCajEB8SxpdrhPij7ze
JYJIZ+cBffgEJIZdJWE0kQBmH7U6sBOk6MR/oZr4SbDjm8POCQOLFlt/sKz6nATkShM/2kj9Hkxf
RDFk2qZaDOsUTLZg77ZWrvYV/29l1tqTd+WtcOUNujTYP7BGoxZp9XCiEsOna/JC3IxmExcDbXT3
OPag0IeAezPYdmC+mq2SyJTJZNGqGeaDUvluVj8LnJjyj5PJgwYrJT5V7kj3WHx6eCp2Dl+VzZmV
EemxMxE4GM+FpX9YgrXG+b+H4sJwespx4eHXBHsLAZG61GMOQaf5xdRL2H0/wzUKhRgcldBQ7+RZ
/hs8fS4Yza0vhuukLVYQwtZ2tUBDHsPP5bOGDfZujZl86J7YtOLJFFXw2/lc7p6gAK1ifGjpzl+v
xhx0dUuDqhkHzaJQYA7A2AKBkBs30/LUb3z8xXHoFS6PWY4a1LFDwAn+q/s7ZQ4zHAAxOKEn+bkO
g8nx5ACJEuqRWui3rFUp/OfxP3lg17svGbhlA7nt/PQl8ipOsPsX7j5Dz9MCoqJuV1voCF3aUyjo
fQKzjB1fJDpT8eCJyUFI7VQyjDSJ0aRNdKhZlzwIe85bT3c/AAgMt22qxykxHs6l4fRPtKvZgYnf
8nmgqL/X5uYwfNpPHZGFvy1G2txUjvJzeFZo2MnnK4WkeIRC5HjfLL7zoqvrcIq3gedgoivZMyr+
mxbKxPMm8M9rS8tzadgEv2JfbhfietgbFXgVurmoWmOtDcG5Oe3YuJNWx1WXuUQFmOBAU2Ses4Od
YLxp0pgsRv5q1qOXjLserG7q2PrI0dVouTVqqZ2zFgLe4eBX34W6txjqohF+3sNeOwM0EbXACJN2
zAJDsuplik4oO22u5U8GsN1UXG6W+cWxknmWf487+1NgzGalrxtXw7gKQe2HiNUsJLv7rwaqlMLK
mMTJkPaXDDszDt1gJfMGoNgnpDwrvsB3Y5+DvJ1zJm7vP6osoQLHLEuNmwTqqhxUkbFUmKgcmyMz
Otv19mUctuZE+djMmvQ0FiB5Q+H+9I0I0H8Cvh4i7DzapqT61i19kffvXUCl7Bq/KxN2VeqjTVS9
ODLjTKxCoVJqHRVpTEyX8NAtre3DhZtnq2glbSoHP6B2OIH0lGhjTUCx4rpORXMaIrRUl1jPKygF
DyjdPdk3vimCCCa8rPi5AG0WR/2HRhLUxEU1KBak2EbWBTMKzWbdGO5i8cghra55rOF+bL8LKbz0
q12mpZnoc30k0KBT/aHIuR/ilj+sKBZDoeq7huGMmtDOPpmsCsIbJKJj5IVoTSNxw6yOwFi502H1
MFJQiCFebkOp1FrQSD9Kf8XsMae2oB6E6ORvhF0HsI+RKiTc474J5PAH+lvexyH0CoeLGyv1I1oj
p+kPx6H56b15nMOkjMJpyGmOcJQ5K/fe8PSFx0XauQpVKrO4V7iCpar68m+l9Z54/2RzDpHJ8G3a
4KSesBq6JOx++6Cu1/mbOT8NIyshdUnkhp8QjWVlyni2ma8gegdznzbDK2W30frBG4kLVU335qH6
vYu9kVii/wZ86542qSSzfNbrSOMXtf6iy48+sGpe4ZFbgb/8P73IF3TBEHwJ/2V+sawpqsu6CReE
vcdkqe/nl9K34DsImHul1lUlqwueeCAJocS68qmqcYUdNzUn2kdpqTwe6mlr9YLEJ0nYIS9o1xWm
gDSSHlPVl9UgA/b1/MGFkqN/1lRD2LNeyfUAAMz/N1U1LA9Jghagh7ORTwQWs/XcvYDQ3uzUzbbz
TmoLZ0ujcj6/xWmcDhxxGlg5nCRXljlXL/tu61xbWtawCH0H/cVRTIdpGk+8dRlbk1ss8/KhlxVh
uQ6/CZGbpzNgFDGbJymgRvnsTi+ohH9LdV60lT28+3AA3aPLo5P/0rk0upjRLcPKbcu+CXVIeJoR
3b7fY9/FyUo7AlF3B/UHqwoT1UKW89no/REQ48fBWlzRXETmRUeSzCt8hRz90x2fS3VWanLsJiSc
Ar6nB2zVCb3RcY0IROfcUaE6iyio76umRz6K0Ybiaq57ZwFoi2J9p+Tx27sIOKKn7O487KvKMJ8r
H+1S3mglp6jJeX4YaxsuHp9GGv/GjMp0ubmmRM4uXzgtPoNyRjjd9l2XnAgTymp4l40MKQ/+zHGF
5ImTXmwD2+wR+uG8mJuyE66QNbnXp7GKr51o7307iySBBflcnQ6P+2Z34raVb9tKNs/0RcuAL10Q
Oq7iCBZgRsIS06NkPPChqbnd3y7Rp58V+rZJmO8lVaZuf29iWkzONvuYak/SSG0ojqUdQzLwsAZh
Pf+IHdmrnaVv81UYOxuAzkq/UXfw7f7bwGh00ICRGuMzvlDx5bxAYCoUHbsK1ynxrzcAaJYIYvBg
UIKn9Yxudp3rc57HHFj2dIG9CxfDWBVXTTGs2RqNnPLwn+0tp8A126lA5EmB0awHVn12d+MH4D7H
96E0mHWKVN1nSeo8q7v2ZPIhrPHqXN6NgGaLR8W4UKTpPCr4DLXJRLrTNYx2OXJBkky9rNPAMOv7
pzmF0RnkIxTSKaCUCOHqzqE6/zv2Fd1dIlzVz1S44iM1186PIsiwr4PDlIvKB/lYTr4EUa1AIOdh
RxXtP6fPuJ/n/roCAoFjFY6NRa0I0zn8L2TdwVv/eTJo2ExOdWWcJwKnFemzLW3EhjLO1arpCUJK
Z1ym8l5jSRCTdKVHKj+dByYCh8MUqFlCy6ofQK6K2ki8NiBm9vOvcondd38aN5hQxrkehRC9xWkU
BvYwqR7vh93kUy0k5Fhrnftt1UPYqQvEvvXpasbHGWrr6WEDSiIe22c8klinEmxZSRhKsQlGMVnS
lGL4oa/Pjy/6BYRajqQx7iJOnH3rVR0a/dRdPJG9G3bTzbxg4asAeS7TrMbi/LpmBvqK9Xqi4sk+
eoEsQoDmACwS7jryWSp48RW+zOqu2cMSozwRW4qSSxL/CUU9hOJ2aUK9gcV8XaNWwKdYyMo+kWP7
btquk3SgM87IEGBL+pkuEhUnA+NL5XtHjr9LgpDYKx2ovxV+XXuReNU3jG3TTsXjYMYTMYMmNwg+
5cJwfTcnJD9hXPnJPxW4GSlhVE1EcvbyIgaGTsAsk/5AAAGCC4Yi7Dx4QsfVnlPAcqoLK0QrMHQ4
1hZWinnktcPjch7m3HXwVFJQt3SQ9HU4ABtfj57z3ntpEfjbm+Ka8M2cZtwvDhD9MEUdq3O/MKZr
4M6zdx/IB9QQs4HO/oow45VprY22Pnk/OWTljA2knSWbs3dHL5auYiSHHfJm4P+W1mminDRyHT8Y
l+Z/SMIpCdindneN9j8Bxi9vDBzksEHR1NkbnUKCa8c/A5LaT0QGQGFx/eCx0EE1hNSxodyvZeOn
4+SomX9PnF4k++VIJ3H4OPGNDuICF52JQHmGJ8aEa08q0XNCw/BeL2y44D+aeZThrw4pE0dwKUWX
W2kxbk6XIDgEZxKeR0sXPuoDhPLFkbQk79nX4966vwH52XS0KvrqGu/YGs4OT0RhExoe4GICXFWl
djWGL+eSYHMP1xzSmaByiqTTfo6xPAzFlwYQktqapLlqzKWe7b6y5FRs3eQ5FYrKnk/Rr3m/Uybc
+snEkygZSIIqs0F+fNmwkg+BLpqqQYp3h3QM6nIRytBHqa/dDTPaJ99+J7hsO0/KFyAjJ8ixGU7H
o52ddS8yIMgm5VzAKNUTlmqRNdTrTgR6h6xFeVpDgFTd+tBg8Y0yFrb9QOmSmef4lBQ/Y39MUj2W
4QTCDPSdsGnRlxQ/M+cPmLcxffhQxlKv728NhRYmQSPIK6iHtK6gB02qjVuLZF0mZebheCV5EhNY
zs7ZMmHH2zY+XnEHM0skjBS1dm4vHJZEY52/K/mJDvoB77h2FSgjPfPL2fle5PO+5KPJRzh6zEyp
b4PpmHNGl3cn7dKrIUg1b8Du+LquwndUJiW1uj1YTwNQ8CFKKpX7MdqTtHUFIPC5COcIqxTanAco
87OAYR8l/SDI+AlHS43gzOJSI6m9NiVCIikDUsmD0YMfZTirhABVETflemQFR84iGGC1kwv7aFAR
8JAc6Euq7rPEPItruemGWlPOZ5RP2s1Qnu6rvf4bOZ1OCzsCjhsx3vmzBNP7dhUv+kP2AX3gDfEY
bMSZm5Z21Z4fd9k2hdwwqMKHy3dz4LrV1Yq/oqnhTQAGTOCJIKRdAogswYWOv/10Utu4ExCYCyqG
UMpsSgahT5tiLaj17xjt0ermejIOQQgdUYTcuNPm+kz0Vdgg5lV6khFUE/4MVLz8HAVJo7noCMeg
QHW8vKEr5y1h+bV9wdgEptQg+mpfGsBGglWrBC11TExxYeLAA9qEH6wFtg5I0BalNklE906t1X3Z
joKefb1PimTqwYDTzOxzuAjqJWtvVjZq7vaV75yXXbsUlLpU1Tw9dmJbB1T0OKlUgavPWE4INH2F
Iv45k7t5P9JGQm7g38q+w6RMH/Nx5zhPTtGHXCfOHyVt49ApTteqcbKt8kS4lk7/lndzub2SBl51
q9xD5gIDBqBP9T8IBVYGz/+Q0qUTHOVMOnxbSo9V3d1txbdlspQuSsrFP+aJ5TznT+m8NNSF3DLP
0p162pJeZ0UX87kECqbR14bO1faMeVA5wF6Mp16ZFxO4+SuavoxzMFo8atsO+F+C+rktA+9I/Obp
43T8sWHHUb3LJNu0AqfZdrcfFRSJNE/S9AjmpbhGVreEgXagVtqN7vSeVo+AfS/PP9ye8JY9cTN2
1cQRe2qZM4tWFZomu1gIJUD1Dptd1XyLi1sOBTAgKr6UF+2ICO10I4D74O7mo7newQKS+RIeHmiI
V+RL6pKQu+Gtgv7UHgdqSxvi6eJUsxXEQF7EYURQD/nC+xuh/e2HIZyM+Wgf1xNAGZwE2g6fQnos
YorLjFLQrib2niaW6tui/4JDbA0PO9iJpzXQtHvcxVwomtfle/kI1NtSgAoAOMs1TE9ybQcoK++R
TAAnKSocScQcAeXBxF5P25E/qicVfzgLz52MItzC6SzpVRJyZahXWBInx6NR7eDgo1aSPN6uRLYF
wADn5GhYePCsCqJtPEMN3SwJTA0zsHN7fmlIBbu+LV9RllGM6gyXBnWMgd8KohqRyE1+92I6ZEqQ
cceeriHZs4E3NIEJ+BPPyofjTIFLLVrvkoZhvTTUekEXhqFJ5UlJ70CosbZ6hb3LOJATpSLoi3Xa
o9uCquRgLEPdquZGnBu3Fdpw2amjYpi8kcznnnugQBEKPDS3UJEr5BUfOTVizBRJOIETXpPTx0Lx
3ko+heZu5EOFOhFi8SmcdCE/y/hK04KnV4Ai9lDVc1b05IWWpXROtnlM5I9MpdiLPp3Xo815vzU6
q61dNc0hoRM2abjPv0kSv52eMw/Itva++jK2Bf3NDflcxrj8M4o2w2yZd/BusPC3nkV0GobKFxeP
PeU6Wt3LJBSoaHjn8HLl1g1Y/SBpDt5voeHNHE/I8CmyZIMK7/kIRZ6EBXi66Kuw42aXUqtKzbmN
Xyhz89ucdwqN0YyiLsyRc5sdLNPcXh0U3Q8yGnPRUUOA4W5A83/uWBbsIgfbgxum6CB0XohGKNav
FVSco6OFrkLFwAnidqzISC5f1XTzqmbxbh81oy++1vtS08M3YRYu/zStNMWVjamcKG0zQDzYAsAO
0qv/8rB72E6i2ESXyHhYJTafqAZ6Fkaw/AibZxcLbVz/T5RN5xtO+4lEL90xWa+zAPLSjRlU1l/X
TzT5vXrKJg7axtrGMh1GcHdO0l2DXpvLUOdgnWB70qEsHPIMw+eeFlp8CEE6WnAXz3FgUVYNagI8
6UOekjgwZgQPNyY+6BiNZSUxL1PpdQYKQegS5xYoB80r2qMcevF0u8Ds0Yw13QPe/Er0reeNtJbm
oh2RIyPTclQdTcYBbBBa/8arqu3YsJgyKahxTaSEe3ZPMVyEzwN+CmqFz4pt9ymhVq9puRDcPwaP
/1vOFNlII3kh1ZZ+HcM+smYAty08Z8o25PNfYI1+7lbhJNyiLtbZtQwKcvC/Waoq0EpcIe2MPKSK
2+WG0LwJmCssfttX5CouqQ6G//TMv5CdJyLuWZuFsnIsCuVxf2rJYSruP+06jJ1ozBZL7CKn41gG
wBONtMVAI84gnr0bBQYRTZbVqtFvhS3SV9MXwLDKHJh7b/7oXv+XeF18Ji1twFYBYBsuXVr1N2Ch
XyXWtLyime0jSNE9MYrIct5bAx8YIuTObB4ij3D9JwCqcXh+YOc3BaRbR3qB1QYFsN+7flN38rgf
s7tLIBp8eU+mLXXvdRMJmOH4L0UgRG+xp/MZB2H90Pd4QWwmTFg5OwLaA7wyK0+8IgrAA/5elyNt
bPSlL/kmqadlqqnbgY/na2n7GmMoMoP+vy9IRglLFmIKI1CnBvSfBhEHkOFWj88L1yjtuNw0hVyS
hY/OrhCWNlix28MAIb1zmETHYp4hq2oST6LrM2JiF0CDSK6Czyu1TafHO4T3Kfz6kYxEciuBwX0/
vR3YLuT/UYYovY55NIibqb3TjWlAuGIkeqy2vqYf50cCBQEpgxh+0ds6jEUPw0ga2VbV+6gJLQZt
svlmlckRL0q1fbD68HEYniJcQl5mzTBnqfqLWGWCyWwFE/IUFUvdnxP70G8Gc7wb7bL+67zyna3f
wKmAk7fQUgLZIZ9Rgvj6VuQCYY6NVrXXHzyOwWwAYVQQYlwmnje9cn1A3oP7JhVv/tCzOo5aivm+
hKc5Qt/knVHAMTyw0BmoQJAUDAFWWUDac4DtN9GeQ5gRZIZJNjwL0NurLM9UMPLiBNJhbRHisjWb
igQfKPJQYNa7XbnfaGhG2k1FH5xn4wWgLC5852I+GTmXWc+bWArHE1K/dNxReXMEzgagG1sYcrYR
M/byrwW/n26c9T5s8Q0pxq6VF7oWt3zFtBCOwHXPwXqKp7Dd/BQtFgi/pgO0P6Fda70m0SW0mhuJ
SDG1QN1RDo/1f13R4TN5KpnHoD3BcfCoupAGDQ8Vz3YS2nwlqhTJ6etUYK8kj9orzAi4E1x7kRio
kAQ/+z3dM9M+A/DePO5WQMKDOYy30caDmziyGZX7ckd2LlYOsp+TLqD8MaVqd91h2OEZQMeb8i5C
0I3hZ+zuwIf9QiBrwWLBvcozigCnZvk7GMcU/mE/r0g6Ptsrd4EaiPpvHIoj5Llr8FYpv+EfFN+D
wVs4HiFThRMoiVgvsB+vSYHocaMt9MO3qBrIsqySwQHhdH04zkEDltYyjGXUeIjz7HWCI8M6TzRj
qLHeBc41eU5oZoAjDYhUk6dDLRVRK4Hzf+flK5rHSydi6fxT7wzsrhdT4bE/UdBBajGiKe7Ywnj3
6HdCPNYHSnhuo8UXr1+8iPuMPJuv9x8jiTgVSWacTph3H7uh0oIaMPDdq/vPt8ZVRHzwzmJSUtan
d3u92i+n/0niy0WzsJqjkTgGvJsm2Y//oMMMecuUAjrQblgEY9Zc9X/YEzzGJZgfykr6ZjyFq0fy
s6Lbt6fSphWMvIkOlAV5oO55iL6IkQmi8KzaC/3wNIjaE7O5cB/3z7wL+YsvLfwEAPCd/h6y4c31
Lp0eUqSGK9fFyQCOXuUPJh9HSNs0vuWSgrb5PSUt9UIAAxdzAtxxsVVkvz2EtlCdbx1HlMgDZRI8
tTmdhfTCzshZlx6jeA4Y3AWXnR/0ADP2BO1oEeaIIjUYWX52pBnVKN9fFDnQugymEjBHHBv0l1ta
1K9ZIBRTI2f0bvNyGPIoAK89orXaznYMIHJgdaSOAx1UDTZmUvELTTW1JgLpPZVO+mzxQFUcu+17
f9Bis5P0X5y7lrAM0xTDDKL1zX57bqahIdy5Dz8zjoZbDNF9AntQQZe6P4e/Mn7wWrcUeHSzwql6
lkvqm21MqUH9Sgk68IQn7RhHK4qUWu8nIDnJeQ7DqYo8YS68qhN6iep8lzUlbr4GULz7L72xef/m
1HtTgwr4+mP3+pFtR7iwKzWQobZ4LxAV8/hwKrgqDdovAt8rFXVzMV8olshyMgFO2+PfR/1k0P4f
IBn5/DkXKeRt/9XKt03UgP7I9yM6Th6vQQBKPnvHqmTHISuwcbS7NGoYnUEP/+Hr4RYaUUIoDW7C
8ZMaS5JSwuMxmSWGs+ohyhMbY+tDFO6bbEyKrly4wgrvo8wpHbOmmAHKuHo1yP7XiyiBmXKLX5CE
bXXE1LW5q7MN1LfFwzxH/JsvzMD8mKAyp3wkGVoePVxpaB7dFZM1egdVcnS731Ihkfka9MDqHqJ6
Kpp4eimNfb4j15LmhroqHFnXA/f1e2+/c+v9DNp4SDPsLQpRyON5+FKfvoQnvM//LEMmHa4P48qo
HaGvU4smcp6dwQKt5rpX31XnVQmqsy1BTEoAREtUZd5H8n6qHOHWgV0seMehwxRldxRK6tvbxbGD
c3nBdFeE+RZv6UO6a4kbY8EoK7Cc7ErmoDpwyXc1qaOnblmaH+tyVHaqPDtPdiYPrtopzq3Ln9MM
8KVfDSO0fZvjrJWN6XaNAH85zT0onQRXl26sRkDikBHOHuXOJ7VKU8/QhTPMiCSmZ/9pyBz7Chz0
TkBerlL39fZqf1AseVmxW1o0rCpLVMdoAnOUakcsLPs6O3qA0F0t/ZcUt1DxBL7RLu9cd/NPJw8D
EFBQ0weH0RlIP/Q8JM/7KGkXIiQ8Jqbo4T51dvaT+ImZXC/LEeH5rI6vpWSneVTxg/Ossfadd1SO
nS1G03VJk+XvVxcXYAx4vU2oDfch68FXHVEZmQJG/gyDBc74CXl9G1Gtc3W35cC/fwq5TiYesiY+
y5D3K0uz30Vbht3dGR6hqW23bV3mOyJhKuIhk0YMZwgs088DHI6ZktImEH70dqcbqt6gGRnH4b5O
g+jv7mZvnppIJP3gXXWAtLcQtdbT8KZYlO3X4J8S1mMcKAX6f/YYGDjaZ2kKgc4KajRI5OnTq3Qr
a262dwUhdemG3wzbR8CjBFMZW7VWck+79Q6B7m/I/NdHrtsIG3wAq42h41j7tKvTtVhAkqMqbPIi
BSWWsPymG1+PMTGtVU7iU/NaDy4VSGOrIUgs3BE/eVYx07AxNrwQjARrr2nN8Fx1fee2MiDOu/XI
kEHEvMB5Q/hCUqPVHP5jdfGHFxWssV215CvPlTpU3IQwTFUo2r8dBQviq6ooB7z1dUE+v5BuQ60X
q6n9oUr4YdGcn0ijq0X8vwwY6cCg3Hs7blxsPKV6BM9rE/G3H0nKZEtYvIFCTyNpvC8UqFvAYWJQ
A1vPQg9KCZNeBjhijqVfAj4udFqUJfeD9WYKfUHOxIK9IY4fFUHn/uylSS9EvJGo7g+d6b0awNrU
8HfIvdgGP/6oJCfD2TNcAz1+fsNajw/x7oWMG6W3uefHL2D1GabBeEpE8AH4qgLcxshlz1nd9g51
wCW36K6XMyO3CdGaGeYFZp+wQkDO+wobpla2LcszUxv/1/kNmsQ7eLRMaxX41yMjjxDgSOi9JIRW
VqNGdrwu3gfl2mVOadmWgXJk9hoRtWYj6fDee3VN5KmijlSAG+Ilh1aJHR768wontKpN73dTBtGF
9+mkmjOirPAfmzymGwBjLGKo9sH5WRiTen1REMePAycot8WnJtx4WR4zHHlLnzGVQSOlojN1rJl4
2u0aFeooHvVMEiAGdBiS6znm0OeDAZGBKRwnWZpN+z/9p4MJnBPTaaQfsyyOSzMrZ+nKr0w8ECgf
/yriJLc/3FrUchmjiKOtm7B/eoFeDy+TnrhHfBpeahkga/R+hPp0sPYkWqxzEMavdX4ZcuErDHEW
7X4yxqqTkfvUUUjHahgQjSmDd5gpzenBVwzIa6iYHFcVgEkeDGNxMnTxGX/CktXY0iRRO+AQOSBA
Ng2Sx6BzO4UgUjQ4AiBhccTTEK+jY9z8BCnmgj7J/1y+jjwyBqLKFqG8zgIX0EPQ9LZvf1dJoOj4
a6w7KMNVbB59dG4LNmBye/eMCaLxr7ikC+7g+AAanBk/JnCY3ZC5uGk+TjEATzkZQxEI7+Op46zX
R7djbAznyUBtW99IXuhIl8iUPQiiUSA0aYH5JOTaAkmm/M4tSRTkQcbYe0PO+12Gm9v3X9VZgDee
R2+8vFeUrGWr5+kz8bZeqJumN8oA6/zN6RlavMQGqOaXgN435gfiS+Wi125nFJFu3bez6YjuTATm
8xIMm03kaO6MkPYJRP4LvelG3Lx8uy+e2xzx4pwBCp7bTwQYGHRBcNCZeWAO/O3oRNq4QRVJmb+o
W4jJeY5q+JRiz2WWzTlid5y4WvuUGZDiZGDNC/2sUFIhO4dSOEUIG2YbvxYse8DABESA+ZwQ76TH
OHzggcB6zYNhHf0JFsEHTK10mWxgWI5ucoX2QYSprA7b/+883qBpXnwRTnz4HNPUjQ6Di/t2P1H1
c79Qysi3cTwVNMkUZJwWjzlH5fj2e4ZM08JX+4gLc0Skq4KZrrmsAGPnNTs+tk/pMxQcdXwBxpm+
2AAYQOa8ArTG9cQAY50qeTK6cPK5ti0NNJP7iczsPGMf6KK5psWLzcpMRxtMgaDR8/JGKOrQXb3F
rt9LSbVyE3nmIVVo+ciHaukiWsS+HeTcGLN0Tj0f/YbsUfNKbsA8ODdh4A3xZKEPr4vHnBIZLlOD
wbNtKg1gE8sG9PJ9dOXK25X/Ohj81ToROSwT7Hk3ZgiYvtL+UoZ1oIjMLRLM6VgsNn9txtHzufBy
5TyNlE+ISLbcFCXz9P2/QLQktPlVN+VS3uUrVbTRUawQAQv7w1a+0Z1zE5eIxvBxswvR1f2lH+uv
BjAwF7bWYizcXM2bSJh5seHXucB2JhZKre3ely/fyTw+VWKG2GO3EudQoCTr0usH5Pi0QuVGn0VF
lKm/HbMivc1+mcNpz6/ZXAOMK6fxtd7ATDAtGUQC6jBZz+UFo7hlV23qQA7QC5fEVPhwL17U6rWs
HK7/VL/LxHSlNzc5u6j9kHvgDvtEnQrGtxdVaICWIlaYDSefm6un+OvqjJxrZgaqPUmDH1ELKVSX
bHigdqcK7PKeSsPCU2HPFhllD5pvBJaaK6j/qIcEZ9tsBRo7qtJtSqcgMqx+I9BTu2wG5lQ/iSEH
JM3naLPJoVQIVpTGy0ekFrgnBzXL7f5ZXYvqSrqAVUadWolDDddLSYUjyyIEzU5sm/JdTBbdvp+I
DlwPgM6y0+EHFOaQ1M4LwecvQT8T4VFAUpoaV7jxVijvROwPLayxFqJYxVNfZIULR7ZvB0+slfSZ
ZN7Kwn7141kvC3c96uxyWcfqw+T3ZiIA38DVpNTB3RjZhIqZjS4AMMIOZJGh0gG4aOyRbv9JHGUJ
PXxHai8i4tWvnSm0cnQWoVGlyGAQYxto5T95DTB27ATgATLJ/Ff2Olm3tMmeU1tInCeYATnoH51L
S555rUBKd/yD3mX/XMp4N6J/GLbpARcSCQEOEl8q06cCZ3e1BM7lQWrKE0QfyB2cBjITE8oPut2P
IjIgIV5GcTypxwahAbezb8zyjufYuMCAWgZeWzYkZcuF9W+vVAVahIsH1hDGkzTyDKl9fUqdKexw
6q8uLVeHZcsF/43kX5OEgRS7B/o6JvN7wa9uD1ra0CTbcvcIoekMroijbTyAKsPsDp1ehlL8N6KU
eG00xmyQqs93JWBAIuZoAsUanKoVVwtJ2BGIFC5XCV7iVY6ONrLTMWL3XAxAPALw4Dyy121bDR7O
pQlBFEHaC92WZN6cbJM58UoWyn2SmnN1Ni79RsObk8tA9qXc08Veq4oy4/aFWx8Ru+t3fhrabEad
6aFLIjFfqLoDdVz5pFGNbUlwGx1qC2CBa1GZXAPDGx7LsMnjpANmed81//Z+H+h+zLsL4Ac8peRu
TxcxFBR+Txs9nz74vg7MexwwksiIO4uTe19434Z+XCbmDfmgSTQiqw3nRSagSDoNoEHDcOjjwStf
SsJF8Y/OTOR86B+DNtRcfsEaP0v6e+9Vr+9baRqNJySArzJ+592gRyGloxlDW0myiEfcUMoFn7i6
/LWlDZYfP1+ozkyetfl8zzDrpESp1P0RyNKMyX5I3bKJfvwUY0X6uhFn0Ps3xKDTVRnymkyYEAi8
VOGWI2d8dWSaPq+5dN/wKRDWbMu7gUXtvwMfI4ByN8vRjKTFFMK1HaZiuVBQcPkYq5gssaljPjgb
eFCwruX7HMWraEivBr47uYlAmsTho3vXgobwuk0DKoq8EvkOv8YzTmc6+8qwr7a90pxQ7lUaRPBV
Jn4BasjSxHpFCzk6KQHnNJrLkiIdUWnjCENEK/fZ3AgLYvX5Z4eCHAsbs9wHc6n4m2J/TLqkPImF
/6uApDiyhX5QfKhefUd2jSURxQn6SU5m9UVlA63q4/fc7EvFmv99rBKfG2Wp1TFNnlnvriK3SEpZ
PmMII3fvI4JcKLJoPzwyo8nTnUrf9CD9OPgtvyOLaFbW+436Gx2sdw2JTkqoi+nUsK4W5IFHqNw0
PJKwnfr0B2ZA0fk3rGxiWnICFXO7IC2oPZ/KvvaXxiXr2xvn7vAN1TpVd8waM7dTwTYu3NTgxF4i
Hx39gubHbpxz1nUygthQ0i2xTJ3cbh4ZPq8WBCsYe+ZY8hVeMhcNTYK4jFYDFYILl5ZKEupE9GfN
n+aUehMeYqAR/6fsopUDngbf045cUu1FSYe4C0PF3UUSG3F8M13jENfMcTI/dSvN3OdvXJRhnokn
GezffoAp8B+KCQZnxXndR+fxLIhMbHfPJ4cPJTYJ/TfGQjrUkhOq7noURE9uUFKp6v4Zfq96BXUO
EDRaL8AL++ceUABp3up07+gjyYmatuImYxiFhABBsFhEEmf38bd1O9dtTB/2oinOPLkFHQant8mW
C3/Fm46INoXxVs3H57vzC7op249mcY5FEMJDoMoAYBsPCpXZIp4JKG4VIdOHN6LB4C9niyIgBN9h
oy371tGXdR1YlwtTPGPgm1mTmSqLCtcXNW3XlQXVlyJmui879ILnLGK0RNh7ZmE3mVWRPkWtOLwc
1pxOBcbsJTWAGIJsOzqKU46xkOSnEmq8L9hrlBe3weywco4LX8TffGdIutjvoS1CdgDbdIq1NVAn
nZzQT+uQIUQdwtiFh8KB6vn2/s1zz1qnMl06XaM6IJjLoeIySc2eGii7UtcxbUtsD5U3/9cdLRaH
7VdRVuYt2mfNZFgPAgbsJnTVcK21LfgmQ3IRxMfMxHKBf0sKtUQVuYDEwP2Q2Y1ykx24Fj8CgK9N
jraK1JYHnwKHMfqdJ6rA7sJVAoBGMOAnQtgdrG5D+5f0Xok6t3gHBwsI1HtpaPpopUXQ7jfS4Xpj
oLmoLAc9fMwun5l1IkSJac+6Yx0hWxzn/dpU2x1dKZUcED9ZN3ht+JWjGCsx7XAv4M6AhrqAN7Rw
yu8BFEJbDKXl0NNsoXl2bp9oILufLIozdPlPqxyQWTsfEei6ExrI5F6Cp21eoIATG89KU0OQUfhm
TYze0lRaPqkGsceR43TsbGnYHDMCmPSvGzkoAA8ByhiiavtbBmjW5YeKN3JhZRLabqy1231SpYiu
EXF10GBmTIK1BNVVkY5RL9PudUCXSCzrRQIDhBeHd7zoHe7PdqYRJsCW/GCUW7fsLtifgCb1ueSP
YD9L5otjW2ADBdQshQgJ24sa3BmZdekp5xkTnq4zUju2DfdpuaRke4ejQnDgmx6b2E+MtNl3c8Zl
T/wLPVYruwegJu/f/9Y4wGAfIwPVkUuYI6C8asBcS+YLLdfsJyP/isUu0H4EGPVXA3cS1z93cmD/
KppbFjFXVxpXaDUGV2nFkgYHNpeQYhLq5ZounLcqWx+iL1v+9l9P4vJvTIpMBKfx0QRTZhDcXyqa
FlhiNmR4NXKOqek6NQOjFuoCMU4ceRmpvSZ887ARvQslFln/WpHGLASSDPOT3ZIFh+r9lMy3ksT0
addDMea+GTi6sweKHCe0wtN1z8hWJThCCQQGdD23AfVJdGVduUSVj4TEivcl8cVXFVt4A+LZRRW2
Jb56czM2F1OMfWkyjMS7e98+a2GdGZsjMbrCwwRoC5w9vkZHnm75gHZ1NdGCtWhCrVD97v3AXNiW
98F+Sbu3ajl6IL0H2Taar1mHnNyNsNZWjGUxaClq1KiAjaEXxQRxBqjLA9MukzVjKTfI4MB0/zqH
s+fOs9OMFNGsmvp6fq8dZZe8esU177cayVqQ7k+mLVjTZj9IwRWm6vYE45eM+KEwMiFpww6u7fEX
kmUOr1rS0zD9mEBLhnR491mtR2T5d62zyVKDpakinSfefVFawMuGpDu90Kv+wXjvOQyLuPnlY8Dr
ScRtkKT510Zs155KPL6IOhw8ocPD4+2eCzysbYgFsXenvwnGwRGPhQvymsLR1RqAbYxLeDRVR4Ot
TG58ESIzP8C9Vl8yGr/pCQfAClhuzUSz7B3hUcV0/7GAJYHY5B1An1gYkcbFXy79ZOcUavIMXc31
wc+cIRIiaiNkDL2O1XyQ5Lqiiowfe0HMg8/TX6qetFa70ACC+4+R5NVo15ySBjHGRTNihxvuZTKa
d8GJGFrtf7SvyDRx2GIOHKF46kuBQtaNQ+eMuq1JTZNhiW1Vc7r7jpxcG3SA8Sng7MaSAVUGC2pK
z6i2Q7/sxDq/Gy65qOp/aF5QtRtgxm4BJXRXWXc1Wly188BP+UJWwrWgFMOiYeVGX6uIPZY+Ei6J
egxfuIDvNhM0vOfl86bRM+3rVCOKG91k00yx5X3srYkzp0jOmlmdewGPC1keD8AJDN+HUgdfEnlz
+/oWIP0hEicjm000DF4GJh0mFG9NKmGuYR5JK7X5ewimLYVe9n1+onJ0k4IKHWjTjgc/BZIw9LBb
Pzz5ocPAy5HFB6RtYpoTLMkL8QT5IIu2hpHGbanhj57rbPGrXt5onKX7ItE6LUMj5rBA3BzQMXsc
nVnvO6DlJvl8p9HgqQg0p8uRNSErqQucBH2MVmnR1DhXCGfj/L9Jj1GSW+udlniP+q/RTOyQ+1ZB
usng3EWh0TLu+E4sePlKn2oW/Nhs3dK9wOs9bLzB6Fc+DtSIPukRFXskBoGzoqxPN8a3eoBW3up8
UOzZIUxfnGHM4nb4P3t0G+TR+eCOhn9UPZXtGW6Pxt/25R7xwQVX/W5n9LYMW/abxwhe+Dcl/wTw
Xfc2FiFuasI4Yf/KcCaVfHSYf/FY9Q6gTC7J/K/MEWNgU1uyz9AcNXczhGsKukyxPFGRiKxr8iYm
P9AI/LoRjn+EtMJ6+fFax3j5ZIE8X5zEWnjuZbXXjDAz6SKl5qBbpESxyPRQC1rjl0wcwcNYMtyW
bA/1pcQmJPS5iHQW+g2oZf0PKLfBSvVOAVvmxbgcW98cMl+aJKy/alUKzsxrCOyovkVo5wrs3mAl
uGXk8S5IgC3cWGyQQFl+viROQ2yrrZ297OeYLQH/mLestuajbBzRW8pHFyM3oJ2Oirx/0+bUxsMi
uSYFTgIAb9M6KLvmIXF479vH3ntuFSgpp1nidwxCNrovEuXTtszm2X2Liq/42Hf20L0B81Xp3GA3
xby/wGeW3zzLqthli+eWBsTb0gmNu6AULXNwm4Qw84lOsu+OjDzALM7BVlgvBU5y4l3G6QWp/zpj
lPdfjx0AdHSOem0+H1mxaV3BF9b4q1MdrjSeffc7362oEXW48OHxJTrEs3s4A6XYzPLPupgK46mK
rvxAroqTagaunWmpgSIziXnF8gIJ6j12apaIyOCzj9M730ZJquMO0fCR/+LafmIKhm9m2kkPqxRa
WsrVNUe+kijxp9/cgZaE0juLHwiubfjxKeSTcCFMGOcqY8Ilj3u0zz2cxB//dzOlRXpTho8cIrkb
P5xikm0DmrLFWE6w9OQL1I4sGrcbAURbO6/b608GV2UIXth2zi7X9ISr+p9HqrH16yI6ja6KAeve
Cyh7wih1+bTrmWaUXsj0Sbl7Ycx1k5U2mB5XlCLn8PiclLkoDQbNxUDFNqdE7CXG0roObLrjYlKH
28ml/rnZXXzEOCbQcEzHyvz6eMPrOe0N2iBcvDBRmmEzSHtcVoAbzGtB3XA6JJSg5Sexw8KrbuE6
xzKxMb0Q0lygczeI5cnaFdcECW4m8a1GXyP0YCZ4ciGy1ezsvPe0P8rjVuBfQsH0Ssj2aQ8q5h27
e5Q8Ttxd9dznX5c6sJkTRAyLCeinaIRP3L3oCUX6TAqtHbdY4ArOkV3sH4KWWZleSeJtmh/bTqWp
VfiMCUPdHug0HB8DBW6xe7Za3ddlqBmHYboeqI6Ky5LZ8ypT4AGaNDgGFvEFjjnohyieA9eoEboi
6vLsHEOPp5rzAgPobxMKCc9bILDybpt9Z6Sc01ibx4qtyFAJzApyxZBFKcHoHSBHiv7TUaCA6GDV
8qhH26xGbB4WOnNlzvvylev5BI0LUG2xnAwDgoavQVQlm7AgWfK0Fgu71Lmi5/2vo+PTclex+Pp5
TRS0cLeZnw3mb4FO+l/N+VXgCHTjWwwMkYC++rPSuPsiAia9PubRqQ7/T/IqMso52a7kDvULyWpR
4WLzivxdMYZCEdLP614OxeMoXP3XJupvDoS0bDzdpg90rW69s1lrzrfaqs+C5bydc8CWeq2sankA
ePj6mw2sZRQTp0Yz1noWb19Ec8u5AT1kXEamETz/K+Q6oHosAr8dmxE4opp7V/bSLQbRAfk+Mg9l
NNFzu7fgQHSHxi1Zq7EpBK9/elLDjLgPNJ4lxC6joiworLwdxIBwJFAKRFUQaJONdtzPQTZHAUIS
8+joty25dpUDXgAqsStFVt6WKVU+eJiqCXR9c+sj39YbUe/jLBG4wUrVeifcvj3getxyaotj73Ck
SXGsWuAy6Up3lo/jYfNoaRy8k2OUap564At9RE6TVDYetKOMUDLyWxqyeLoV0oNpagl7ns7+Aow1
bmcDBdRkUV/nZCSgdkwYudddc4nQMKX0mjJeErC2/+9PYD50/I+83X/XcIcFJoC8tF8ulSZXcpKv
p8SLvsRQ8KBxnJRVPIvQHD0M+mJlLjfGxSPb4P9fNZBegZXyGuHqT60Voq5ac4NS8cW/5QQQyrUS
EqgxzWJacG/njQwU6FCOAlpzAaD72baj+YAChKcnhdNAjm1j4QdPKAbkrrclamVeYQZ9ZgFl6Qs+
61pAtELMAuGx+lVZ9iLFkJd86u6P6Mt6g5q40nLYnS+joRXzLA17I5rdmkazNyVukFrS0NoY/fR4
Kq6mRpg4fLezevsu/lCrHAyz/Bv0ukqcTapCC+FivILDUMLokedDnn7hmWDHceIHpy+l6wuZAhkM
VCIqxsjqKOPxTiWofPLj9qE7lbB6ZwAOPgblGwDFDA2ZihWwjyzMdG4ll1FIdPuMzC1xFxLGtmWS
iszkiQkYibPnbVrC1z8nBg67V3lfjVEyItraUjYw+cY1OCuMdM6WFZEXxHKHFLalMXUKXbwfdrmB
q/N0DlEX+zw2YfBmbo5WjnVRsO1RgTrMY1J1H1kyBg8w9RuGcFgirb3O1D4pqlkRdLTGVuMNuQ+i
e9nAcofRIlDctU5XygKtmf/Irfjtk5ANG8PxhJY2dBPifAH2nus10bTQH/4Cw8KoEg0qFotMdwc+
odeoTLm3lPKobPCO33TBqZ07oiqWbto+wGg++qzOG6TAS9uzQASdZbCHEMIY4AirqcO9Vyu15L0A
HaCq8du/aHAFfGeHpnumT7loazQ61jXnCZEjnz9lOT94tWK/JIy/q4IFzpYpJ7+8uxIZNJTkSrdj
EfVADd74ZGGsXWP0ExaUJlGiT2+5F7tfJdMVrlg9kg3raz3lqcQzS3Hzph31HWPgb2wDog1Fi9Pp
0lDkErPj6zi68ne8J/yOxNGbnpo0UeA7NmlXc4AJuEN8hpJEj94YXmX/XtPohQP+DCAOnZH5cbaU
qxY4rwtGenOw/pUdASHjy8fWPWvMuIBWTgq68HeFI6Ikk/HoON8J2yXOH+UuiIlelqvfPPzLc0+p
wEeySD9TMrgAWikicwTHIz1fQKraRq4gYKIed3EtvrV4N2sIx+DT45L/PA7CxK5rK0/eInHIqNF9
mKmeMLMHqaRzLsRwSvo0hTH70dRqIoji49hIGcLizfAVKoxyf9t6HSgz6rix/RI4Dygx/ls8VgH+
SW2l8/AYmx1yvQG2kEwYQRmwvMwysk1eg8fh+KNryKj3RyYe259+UgV1qGbFHcWLjZVGUpjOnmSW
M8MkZIF7GKvw/BbwpXw7DUtcy78tJbffVDv72AaSzvxHOVOx/whtdPU3NWkAbfGMq2CN0HDz2WdV
Ax/Y9pOAw3pcYhwDjhaZoxXc0ylpdOjX8CckXwjQEdiLUNnveMeN1DNfFetOSal0op3BGMZwGV6k
fsDA+F6BxHTb9HUYx3ti4otpx1dNntYonZQurwjdDkmQY7nupA6uGmlp2a+arJipG7IoEK5cHC6Z
choos5fdSWGwC204WQwYqonoxuZlW0VF7V1fF82hLNo8JcK7XbSrXPIjfw9xz9qh/wjzpG0GntDV
VPqeskjKFVCZZJxkEW2mXyY73Ht5Vq8Cw4ge7z6vtRQvRcxExMYrxKtB0V3YnYj4hh8Jf8HOPTxt
NExRynPMAagQNx0kFJY/KeMrLl4FlS02zWktNtXaUgkjrYUp64q/o56XMjFqjTE+38EXmNU0fN33
lSfBDuaxYviy9NZ6N2Z8mfOzicRfUNXquzZrX4Vf/hhCoRz+q8PjueJ6nttuJynR0n4IXhf/DZp9
s+TDYJNN5JmMoP/OIAlXw/gBPIm3hBKSGGDhOq9dhaTylBdEGXWczsQmIw5WsK8ahApwOIWkL27g
IcWQ+PsFJrtZkj8zL7s+4gscnjM4Xkw3zq+sy8X0BvaqvDdIDf9s+ZgS/f4mBmdSIOvoVHxjZ7SU
IMGr8xFt13DpfRsCkfGC+L8BltVMBg0LRBz/VLEI2Qq3SNQMgJTiFVCgxbj2ChVqU+xj8FaOykXF
mJnHtW2SmxWPI/GXG9EMEXqoJbxAH4A3IsCtEUYmAhVmdnvn7QuQrE/qGeT8bTuQPmb1isxNW3P7
7KrR045uOKzaQRSQXEefR5tGzwr7mDGzM6q/whqKNbum+2KdZzwv4NPcAS3ip/iJuhJsrIzP1atX
61kVBG0JPfmHpzA0Z1Wyu0IqpRbLnTOYOSwumQMM924WDaJttFCfyCFANKHQFCXgNYNvNIrQevtg
DyIRbFo2y3dfmPHRDfkUBSDT1eCssUC7RnXort65dd4gxYSG7fUNmrEX4cXUT5eSPsDZ6Qt6qEYH
bmiKdgQzLWrk1Be+yAAba10v4w+pSBtk5/Vfdx5YkFAW2ez6FDDuGBPfkMAoXNebOmQQ3ML9sSAs
d7AAwxtI8TiBUXhevdSQX2b31YfEfMcqinHnSy/sK3hNnFXfXP4nhwaQkXrNOzGgmsLpQYLmqhJp
k6V8QZ4WOeZg4Haby0J8ac9Dra6CIscwmYFjcoc40NIyO3/1xg/Rwl2oGsEwnRkKSCu3w2HktrFC
6MbNQXwPZnrEGpXkT5YCSEgqHy0tcXLTohjshw4S694qFGo2ydKMukE8yrWEzZ/iRP4H+2HISzqv
IDb5bwEKxNu2TTUENPBd1b/B3d3WRQu6Aaip52XhThT4NmBsrYbT1DP0ZXi2yf2Y0NsL47jm8mT4
La7uPB6gqkCyK4rikaC83/yu76PYgH8h67ROPTqHJGXpCdudW86kR360beESFC78ANYIwoLmGfXd
I3gYE4xY79IswBSzaCAbDkhU8+rXjwP7EF2YNiUvSYXxnSF9gG+dd2Bzjwx2gJs10UTh2i0whsdL
E/eG3VQfR3Za6hP6ESRO9N97/a397DUK4QE4h3bRC+iLixbdGMg/j3tM/rRQL4BRNeBWVyn9UCSg
aQ7Z1RIqXnhhsXZ9vYidoW5DMf/zcfBneJSf3cgn+JqtiJS/NBtwSVi1hb5U31LPemrdEwYO04MM
TxrSxkdeh+GVkWpyq/1IE2LqeloE6Ct9apmmdp5jfZMeG9TckSKoAg+m2DJFpT1HWvP2wbfkj9AN
/HNzOtKxB6x1FmCjyjSaKhhvrppUcPDsH1yxWW9ikJHpEnY3kF3PgBQB+owOYwF9KcBoBZk/Z/90
LmOjsByQh2JGsEUVM9mvdXH4ANBVYxLSSZC5niCazKHgcWZvWEJ0yTWrb8/+/cmDRc/s2h01A3On
P97BNUfXorSassW682OtaOB9I8P+eIdE039sMaPkZCjouQKJMCV2IW7FdOq5engJBcm4QILhpEiU
azmiQV7YvteT36HY/mrWLJrjHM6xzb2KkaBSSHiV9EJJ6klrqGFldGNwbjMXgQWon2AU7JyV1Erq
fddy4sXO/+ifg8n685hlSwIKRrYg0GhDSuodNA5jYTARiUjO39amGd2DIFwy0k9Ejd4rStq7KOqZ
6lpI0UX0vo3p26aLr9PkWat4DN516v9/WxBCe7r06oIkryyO+YQ0QoZb5tubulScuWBV5rBg6fQ+
L+v84ggMixmJYD5iWswFJtHCAh9z/o//w2mAVlL0Ym/tMKa3aKnUkCvD8LoBZe4lWGmOzQO6Sri8
UbwuFFuIQq56/6dqDA4xCZ9wgR+TTuY3zDlfto1Z37ntH4yR52dTv9QYo1wgcJyc198gp0ivcV1L
9aaAf5dOS2DJScG9u4z83vv2K94mFGCCZfLKW51n2STjJkYCDj30oeRS23b4briLRJD/C+2Ye31L
5m66SkoK8lSOjfp9swaXiQPums21Ao96YcaYE1J1XVKFlfOHF4uMjjcR3eGVK+/DJphPLO/1gqa7
hh64NzO3sfJhw/8nQLDfNPI7iwnawgWcMNh7Iu+BPBuP5f+Iw4IhBaW8ZRrycCoGERiaIn3xWfPl
jWYo//3Cl5abj/+J1qzZKNwJHlRknmGCcMmg8QEk6R5qan0ET+bHGYIkQ3JUHJ/29naBaNKTY6XV
cpnwb5o+L0g68B0LwW6aGS7aNjm32O6+uthU6CPSTolf0Y/cMmG8IVprZIngyqTgUT+eueL2nzCk
mOXFehc2FiB9eUQ6HRYKt03CJf5ve4PsKMZkrY5/eXvNZBtJMrh+RFrPhSNrCTW8GWLSjP6MhPPC
b9Q7SVtRY8WdAtcbN5bM9tIDpvitEbX3g/HRhiPGD39/G6QoVPS9tQf9fXMZDLp1/aJmX0omMFJz
gCbN95qiMw8ksrYPE+2XoMymb2bqU8ikFiKS/D0DBpIvDfH3gh3Tb/dh8V2qb6G2X742x8UjglWc
W7zAQsuBz7w6iVvAHYXYd53uLQgtoYeIffsLVMFvbf6yfBTsB5B3o+Flyfn39kbHXZQdzsyfZSEU
Pfr6yACzI6qrjFh0v6vlYDdaI6V5rznidymtZp8fnCdyxf0AoXKXSOhLXjMsKrAYWOsFpE/Mpu8r
+GP/GknDGD4bqRt0gIf9kLDgm5+whNPUXG4NldKYcIYEjfU9k5y1ttDMFbwZ3saW7rnHy6iurq5x
/YKpoLbVMnlUPV925W3BWCYR+aK8ScX76RePsngemdo+HwP3G3VJKPvAGhpQTZLgiYczCjIZTynK
/Hdw3/hGbj+x24Jm0/XHFhLlBHlnLCFfYjuWU67iwimKpctcfg8TLFEROmQzyJiSat6XQ8fG6+aA
Pk8oHyHYzM05dzoXRsLNHd+lDHVqOdN9Na74ns7Slj+CESGNp42u0Z7a5rs/eIZV+aJiyo9IjJpx
zI99H0AM3ErZ792soAzioOdiQ/xMicUjonEeTfQx910/9lR/nLcBU7A4DqNrf7gOXp8OGDH0LjiH
XVS4RbUTabRrLG6dwugoqlUl/TGJrVtDjVObkLfI4Fvhkw5zmNij84akw42h96SQU58jkkF0dFuv
ha+WQitEfjKhU10vHWD8Hgef81jVt//8TL4nF1W1u7WbGCuyOW6P2QXdlM6Mnj/JMYk01hiIVCU3
9rytJkPSHnFFC1cripx2dJHKJGt7nBzAQfv5M/Bo45leaT3T6ChXfyBDY00bd6i0u66+YfjO7lYm
cnI3wBCHiCFhkMUv2U0zW+LPUt+LO5ATQqdYQlFw9D/D8uwng4u7khrDBAQI9vU/K5syaVj8Tpre
4dDIAN+T/Wkmr+72uHqCjubcyHQyLcOpVFnZ8LonFLAJcie85yorTok5mBieNiDoacyOPsqGn6Vl
SyvqtN7jEv1RboZl4i77Iy4mix3hXH8KIQXbOiUFr13baUxlbjYTzleHkJeHdTdDcJGj3sQS3BWQ
rCCU61qwXBSwbwW9dYcbVbazROro1u/OewJgAeBI5OMrv6fzbquV1ZjqbofzKZ9YXDno0cZzSL5v
RnwvnXVss1MBOo95jK61vrXnM/LzRQBapTj6FCJ+T/JMOMc135pZuQMkGrUegMwQgBXWAUQzx/LA
459a6HzlwIWYKiUdUL5+D9hiX4k8jggpQhEl8E/MOZuP4wCfkJYvk/ve6MDsA5vmxK933OAj2R05
CWGVnz374f58ON0ewyaierzVTar0NZx2Q4T3aBConWrVWUu9rwTsre+uGhyaqml8H26OxuWlXxru
HEBE1fUHZ7RuwjOq2Qv2ZYk8VcfiIwUqyfoaHoAcMR0JEvlg8BMuLyjSYDQXZSka6bXse7rKngPj
xb6MC7LNc2ECte5YHny6tRRQF8PIwclDEdTs/bBhNGCNlBleZuOvBtupGfuqTlfFvf1oZOcWesPn
7QgW4Mdtxj7oqklFJeA1cgh9ruv1oU29Ve1E7JLTVnDkNjRHRgbVQ5T5r2EqD7fb2Vy5UaUHxxDQ
i+9UEK9RY+2nfQSN0sNMbA8sRIV11sWnJgP8lPiD+g5WW3fWMUnKVteOG1moSqtFYYWE4FvwG4St
qIjqPcUpg+UPIKRudcLD3yBjxpiIZIpc9GTwKGk0jJDCiEp3XQUg0ro8eVKDqEAwvEk+KSuQbUM7
eIXbiPgq3Gv4LNmNWh22Pm50SyPAR1Jvn3aHKOTmaI4ppU6gGcWjIfyK5eb6CU9vye2XA4PIrOUf
tizB+ZQbehqrExEP2+GFfs2Q3osBL/tl1vHPXZNXmqBDX/ndB/6luGaKSxHEx/ubDfk/3gFtlxUr
Gbl5QvoWUWDg5lXYZSveMSxtHrIMX6OiFvjfDD+mzf080qzLtgQCxPWBuWUBhOwXz9FtOiVnAUvl
d6ybj8D0X2t++j5Ilr47+60ohKNG60sWAG1dL+zeIOx0d2dzPEYcXHOCUIWWpG7jbf3ZvjpChykU
2OTPWcYh9Anxw552ILTFrQpEf0NVOe2TJgHqT32eFrQTTNME5aN6UdXP5cNk2S9ZaZul2s9Pc+F/
+VZyIPQktCmUaZNCiFSLVp0UNUnHOG4yUdAYXgtfo9bIWWvXW5zb+x/KRhFmLaHxGVDCxJxffh8y
zkhrCprCCmK8Lxcw98i04uZXCmdjrSSMkCS+SNVdc1TAhOZisV6vCnlj8DqFORtjo8e6MJGDzNBR
aRlT1qihA1VLYvl8B9nbnqMc+suuxX3xwcURoDm63U9j6wONrSc0j5Ra78lQJoICE3VpdK/ahH1F
YwTlRFJ8/Ejw+/MvLvWpTbC4wQ1VY5Jggj/s0xGOp+DXlJuSCs57vyFsAQ/Wchxhruet7sSEA9R9
5HqRDQVoO9zoUNLhqim/Zs6Wn1ZGoF5E4+2GwyEJu8nSONmZa+mL9dN6bvkR8Gsb1id9ntGEJX8k
9lDsDPeJ0MlVA4yU4ZRXi5cDNAB4Kx6UOZH3a2EDd6vcyPhRv/6wkA/WQdEbiB+Cf8O7KO4pkW1t
P3fnKFP6wsOl1zGe7GWxxIZSgY4xBIk6D4jqYcXb6KuJsgX3C/a57bzj0/2LNKd1oP44JklrPefs
oT6QcZNe20jH0Xji4bkzBW1dQ4fSBYRmS0c0m6ppdBXkqoMfd5Pe1eKM/k4UFdu6sMmKjrQK0Pvt
nQJv4fdSfGFTFJtABWWFpzkaZXOzMIS4WipXmbIw7/Oxi5HqCsNfqitc4e8q/lCggomV4rXVMjk7
5HrLxyBEvcjThy8hjiWuVwE1dsJlJay7bgfG72mZhtdWdIXCDjID5aEpvGiGDOAEHffFOWhBS1o8
ZmQrRxOm9fiPva+VO5HbfWW5yCofUhb9FgRb90YypxuXFAfwC4NQ32ph9p+243JLW+45F3Vu8x7c
d1FKgSDykYXkApq/dJPFGX3lpDL6/VE3scjKCEtogcOFKSkSVJG322B+ljQEaYNiFy6cleTn2GUn
DlNi5ZPkg/ELvxrhn11/OZFB8TBrYRo8fbqDGviK9/uVsoikN9NDkCFJi6Vmdtv05toHiSVyH2av
v2guffD0kTD5h1RgT93i0zVgRJZzd2KdB59ZtWmWaYtDFNH688jKs/JwCINiQMF9ivb70AIEJKH5
wdQiEVAm/iK/TmMy4YhaBxMJN7Uy2X7Iet+NcFPGhuqOaOn/jV20eO1/D1V5Ucl/mAho/+FuWxvB
VUX7Cdakes6ufgHrpSWst/tXsT7XtjeUDti/o4gMI3+7XlyMBM5NNw8bL/3oJXlkvYo+2k94PBTf
5x8tySmN+xMULevfemJKGNdetErnota796iHv1P0GaDfDJSzP9n50x5pQDWMAynMl+bQ1DNGgW0Z
fACki9yEWhsTC5omioy+UwqUrXsKANaKJD2TB9keelsozrutToIe3uhx/KMPu19LBPs5wAOSHiMe
8ZtoM55Df9GRsSGfLC65Fk+JUzF71WoB69l9UWW3/hFRFlqqOmzPriFd29gQDlYWoNfd2i4P7ff1
v7qqTXRx8uCoLDInY+hznIn3DjVZ5sq7nCvtxVd3B2m/hhERJwUFSeizn9Z8e+Nu8My8wM3bfce8
e96TAZ+6KVvFTnequlJYQGMFGZd9Aj3KodmhiGlpt9qbXPJ4yvP9QLDhGTeIYdm/CtGPTR/cB9YH
Ju3bvrWrk9vIxb9qM8Fn4RHJlAh3VoPUrcP0jUNn61oiPTCKq8f5/HkjlqfKxps4AileTvgxjQgS
NK/KEEsGEDssoK3tEgX3jDeor21RMv7f2KHIDLTSf7epu080cbq1hX9q6qNzrdcuGYYOHMS9jq0A
e6TaJ3uwkriwKxOYOLwiXzFjMBXDfodgGz82munKScBZYFC/o+5kI7AjKuGwROAQixWS3t4u3nVN
6BFwyEM8uzMqqUknB5FCWWN6kjxvekVD/Emq+m9Idr5NqdAIsIZeEG2E26NWzH9FlTByuS4nDOGS
Cb5ebJhogh2+4wAi14I/9tl8+BnRdw3xZ7kh8VosHtsoHspSsOOp9fY1Huv2Wcrw7mCUylgVDwC9
QZMIeb/8F2bq6W/IsP1IGipCOFeqTVt0G+TVjuuyQllzfkb8dIsSEXxLDmFv1bg1UK34FT2SDmGC
2sW3aUbpZhlVUfa316uk+HgM6mvreja7fwbjEnsmfq7qPh7Zvswb0oN5Bvos4n+stJe73ukXgBCT
J26fnpzVYRU6XGgWmQZ7uhhlnDDomgpvWI1oPq9XTcLjKQFHIFdFdi8iy2o0qoem8W7XRsknrmB6
si1I6N/WSTXKOSg0SW9kwLpOBEM9QJDfiKoI7d5CFsicchfMCeHN+z+nV5rQtSXeLvwzttEdIha8
pkybr0Lp2ZU7mq/DqUYMR40RGCjjqJnDda0SrHeqpFarQ5MdifmrKV7en85sdC1fB/rXT7UYV1oF
S/S1y27etbI782DnCDKkqHiOLAPH9cT0OlDrNJgQSGIdXD8/YyLAgCyxh7RvCWdZouzQNDTdGK0f
S5EdqCDY9gk/LsJMeQ8v7zfsV8lAusmw5LaOlh9MHWbqSyDRlv0RGfGwmci6ZJc+gFrMroBHDlUk
6s0fEDX8QhNj9cTLAWnPbGinaCAwtUBH6dC51ZvVhZghxoe5BNzQqYDaPdxsaX7EsX3Bv8RVXSbm
4rEXUndxeFMVQlV3+gMVjJuOHbO3550G4LJ6V8VmY2KhTrwtFH1RDJE9FtRplrq60afIvB39KLFp
IlkornDfow0U91A2gLPMe90dooTsik+z3r5DA6MAOR/kyCtEUMqnTiI7R4qtb+fmKskcpWrdqKRZ
FrpIaL40KcLxFEvlraMesVZu7anIZV9ctMF8xV0RzbfLaRNrTO6svpDTZ1+ZlMcHfk7ScBLsdgNQ
RV5Z5oiaITxMRJPKohOgneoSU2g5ajijqln3DRuisSrjoJMuSSWTIGvbkVG4yWdPgo/EMl1DCUGK
6SdnYeI+zF+/kfVPnzBEtMVQo4Ol9sukj7XslFzQ2ZwFjRe6cHZ1ZY/zGZioqY+rc2P+zxbjIVH/
ngS7h3gqBRMs78qCa4cFmJj/L3mAP/Xwiky2vBKrTbNql4xU2OoyIVphGOWONnzp3Jo0mCaWT8ez
TW/nqrcsym4qtfi2qxzKmkKeTT46pNFbS9DybnG0k+xqqSaYlELO/WgDGlq8ZaWwxB6s1GHT1Ho8
Vh+sIvWwQLQJtSPxIZ5FKrj5B/M0BDB0NvLGMQuFgXmY+Ol8bG6mQ6dja39RpqNCjm5WXWaNejdx
LV9s41FOazLCNPr4BHc716NkpgT4BFvMqsN2+QeB9X7Y2aklWEwbfrO11EA2CYKgJVEKDLf1TxkD
gUyMHUP4vuuWE+XcPfL8ZechDZtVzFrxy98z8VbpEUj1cz+YP/8jfEboLH4iiSAGjS7ClKT1h93S
H9iYeTcUYs6t5heodPywPb6VK5GbrtNoc/vfzJSiab8C5F2soa5OMwJUUDAQSNiM5V6obIsMj8cu
r9xZ91SIKoBDBEIi+SGIoDXhc+DyboSM7bOuleC0AThZ4ffXmwwzlCm9B1ymuay8LeCi3ZJPHXJX
pQ6UYJoozz1WH0nsu6sCW5b60C2SjURfvxr1Wdm5PI9TfSQqBI99mrF22CPdwFoJZPTMQ+vvoOSB
oiIoeTNfUfOncIjeHehlXh2T0IWDmGOXky504PKvbICY1/YQGnItQQGtMPDExiRLZVlF5SATrLFE
Q1PbD8Nu2losCbfQwo7jK3SywFTDHwS/OMJDcqsaE4SbhNmr8zf5kqhkNtYGD0hH/rCzDSCmYF/e
KiHrUf8WWM+ExEi3hrU5zZn14yDTAlciwktW8+lpNYnPzl4M8plrf5P0mWSF6VCp7jQNqqhCzDM+
OXU+YpQjaCuRDeF50plAiIP6QXDzwI9K80n0NVaf2rkbrvNyV5ECy0+NxwULkcxdSbxjg5trbZi8
bsjNsFeuhumG6v4sHuiQyU0irqtsw6v7U83OCrfberjLWfo/cXRz3LlkIEqmGMmf/POmBcorWfRO
viqJi/j9wZLr3cki7dfKrhE2gAKDFg+2lt+ZUG8qPGuTdxmRDRaTzx6Ps/iNI6uRQYNziOCX8URl
wVNPIx8FpUh/U25VS5BSBdVmlr+nKCMNKTZO2rmLiklc4pIm0az2RUPsJyeqAYFVUwHkXr3Hcu+w
nATDU6ezYD+/bhuXsrsUYJHKzihRnlYwid0JyG+KCY7sMPpXz4P4Lj+5pFxs84y8iNmF2o+ur4Ag
D85EzoIXMpKKwAs+Mh2eE5GzlA+fV0uLoOdNBVlbyVQ3VEBPnG6EdkP9p7Xy62uBDeSV1BUDbBh6
j62lQJhO9tOQhpNTPFC5Lrggtnba+Cdqv509gnz3bPfoHZ5ag7KDV1+4EidnbIeZR1gQUjU4FYij
KQeb2CYMODWH0bbv5Uj+PhDk1SVoTrY5XcmsOWyiwnN2kGrD4jUXrTQgNhigRi+hLq3EqqPG79kX
tY7DSwvWlaFQsOw4Rr+jdMI/+3xwdxZObtfDm0H9z4oLJN0COtQQK5nCcevE29qdTHKA+HA590QG
wKEo8jn2rcmjDQ85peYbcAxQ1nWkhPQMrhXSxCVmf0mvRIdKNe9b7eQ/g6fLYqv/VMQRwpUyqznS
dH0l9+ged2P7wPx0SBcZeqwmK53auRvNLhf6ivzD5Lt/wTlHzvP8O0HqrRBJ5M6WyEFRw4Sd6KfX
O6gRNcXDB0B7XhYA6tbxa18m7qVSciOVfPYQ/gOFGSFDU9N71HeRWvygH+kBTIHe4lxGy4NbVF5K
oAMn/PYS8B3j7tvTy1bphnyJoI2xsJotIOgCVjml6Vyvk3CDW5+w4JTl8YqWrBSpADQjSmdX/KHb
+O1QKBIBLxBWJjd9LD7B5zqk8YKOsP2t0clvnpq5hs0+2Rdk/JkZyc4vNkU+zaQkA7m6akoY06zO
m37MVz0iO3bECahkBAJt5gexza6i+jWwupoHiaxUxc7Y0+7P6Blqx/dNmInsVX/tB58vRmW0LLMV
nqWnQLFBjmbRYQBgDZ65S1fxnQvFdfd/pndqrLcOXv4nH03Nc5bGUgI1/ngfEN1F3Lll6MR9uhcZ
zlCx+hGm17iHb1cqri72OfZjqzcdfhDkyDZ2MDNpFVdDH027+t8ax7BaypNBJoq4K0ov9INCyxpZ
1IT4B4ztUX5BpUkmY9/MreUBtbh8qleGgOFeJzBmoiB1VMJmIW2thuf0ZNs0A/Ie1OI56WHXsCmQ
2YX7plTYMxqi9ckKcoM1AvycQxTQTGo3ZARYAUMSjGyuN37+fmlyfjfdnWEdBHsA9vod5Y6dbiXl
uROVQn42eA+qYKaU17CYHxixazsV5FSNlm3h4ZHqSq5ugaPJt0ATDNiPwoBfPbnk1sQHjmaog7hp
5WDpSZKm4Ae1wL7Z/7VgC2OA5wHxcxK+sS11XD76WRmm5m+/mHOZHNO3Tkc1xt2E+v42jr/B2r9z
p1OQ8IbKWPqfZvvfKgP0u2LaIvUMBPPyAUBw9kqmw1coVXuFnmXaK8nwVZS69CBidQfsnZCJvXYL
05pCSys9VpWC5xjH2+3oLHyjwH8gjcHHlCjqFOhxD734EoPtjBG64AVQhcHhaw2RqkJv4TnJ3HiO
VHLoiqULAvfIM1VQ3Zy8bmd6ZYNJbdtKVAB33ARMkNAZkQxtfSRVPiiuXKxbInAnhRXd82unPj2N
E+Xav0oGlmNtK83AD8cdiZYuUcJUv2t6bfiQ/Gm6WsWPKU6Jybv1cvTlpJRYZcE1xn4H/sQOZ453
rUDNk25Z4wJFs8KU+gstKZuuVrwy0vYJ7xTc/myQ7YyQGgjuAFTIQpEwPvsC/b7tQlrh253phmPs
/wTBD+hw2KFkb6U2hPrIGG6mAEjyfK5BYkEKvsUTwF+pIJDroh4+/aEQWv217T3tjvu+6XlIoqi7
7TeXp6XFslt+hpvGm+jr1qLDOV9wjxaETZL2AtB7z/SSlgJLz10OlOf/I+l0BKqUmlrw8ACFEQ5I
ypswpgImSbby5mqjIp1lQyc5/8A7XXsrmejQOk3x5d3Ug51BIBWSiCr0jf0BYTwvoLTykbzNky+x
Lvqj7EJZ+nLi1HYJ0pf9vOst2YMWpBDMKkdnoh6R8q5JF6Q3jcg4Lmb4CSf0/HgKEWws2h9ijfA8
G9pQzEZ/8Wk4P4ke7QtofUFMJFkii9/aXmgRjIPzkPKnD+Taw+/+ei8CGjJH5iLkKbume/Lblik3
lcEDZ96CoFJlpS61/FJU+knXXqIEiheoAs5BgPeHiZN484lj23sp6SJCevhVS7U6hJ6vDprrzddg
zk+EPswUxo5yettWbw4bYyEzqOIBm34NRbhs2F1dYJamooaHiPvg3QFV1dMMxdQL6Q2Utv5KqNSm
stLbfvEFp+ocVczcnLbcSXtdWt+iBac0YQsg9kzwmWoNobR/PstpoIb6uv0o8ccULZk+lJ6RjWER
5Dp/w6M4a6LBreu2ksmCXpoI57NXHcAFhK9Z2ihLwVSW2/ujcdX8mlbfPmfKqljwcsSxEOrnnrvT
OD3HBgY8jxmhKW0Jz01Gf7mtdvrONUxflJhMu1XJhisrylVOLNy248tuuJ80XsF1SXqhtL2vyamh
wnaLYRZp95JB7fhNKW/9S89rddeG/yfmo7NUQaioEF1U6D12Jsl/LrVxsNMGRi4zUtr6hah8Q/Fd
Ap6QG76hAhf92XMf66t3P/TxOXEjLMSOBnuYHF2NRgDSKMAEkErCLKahBK/NCArfb+W/XzeKu0T9
fsES2H4m4JiugQnh4LzHign2Wcn/hG3xUCWvSzVJ2SI5wSNfDSqiI7hJKjQ+yt2YvKXZQlaDRotc
JhPmOuM+AlZBNfHKbqOzE2w8+j1ZGv1cw1wbmtisBC0dmy5J+M23Co1tx69cHLgrC5EQvcDY3p37
5vps90j6C/DK4ZK0DUxHF76TF2TRcE6N/jsky2yxMqomdADrsbEA0EbYtvVLWXbcqxo3WYdDgXZE
BmYw0ghgpE9SOsgrQk8bskeJwC5lnH8J2huSZwLxw975drvvAv/bZVt7sRvQNhPedGFkaEKLe9eE
H483Tm29avB9IxYR4Vucg3qqzEzKd4lASphoRRDdiCz7yssE9KeOlTQVVRWeR3rW2ktxEPY6Eft6
x084w41qOo15eya92n88Kx5635TCYA4l597bOn+2nQ5Ot8rmXrfFacKri0LHKbaJ41MqB4e+Znz7
WA88nHXiylJWMlaqj003wUWVtzvEcI75ZEIBuZpJz9alEOILdbROW3QF5lBYizU8QH4cPh0g20i6
dEroIw+omDXpfiV1USYiIqZg4D2HGMDyspMVZvgRBm6Wq47Js+OXK4Lm9bIm/mK7aBaGWwFFWgf6
Me+wmnzNeXQwAdQ9Usk1KQDh3aZY6WH+EkFQiyNfrZVcHuifUcpzXUL6w6qK8mvDSynW54SW38XO
DcTwOS/qa0d7otTrPyuwKxagsXiG7Kdf0jk+zBHKo6bt+69UM8Gzr/6SLs1+iyd1o5zaiNzuUiQk
wk8bQsWi0Jkb7SYqQ9FBID78aCY/bCndfQaTk9A1GrhLW4S9/3ome7Pk3+hf4kdt+dXPaUqUlXSQ
lHjOs+9z8q2A9VVPIfQvQlQxYPllwR+jh+aOtCBfQAMlnq1zIJZEbHgKEdZIBd6np6BDK7HJUF7U
A5X4ml1yRT87zxhDp05bSqLrXUmkG+C2UVqaxNAIKT8w0qa5yRvQd0k79yHUdoHy5maASLlNvOSD
zLupMAeGNXUjlVktxhtMDVoGP71W7vhrbJVuV9XT5UtXeqz7sRtcXE604XOIi24ulB1CP7fPzmyE
/cmMJjXE2GqS8rbMJ6enMKnDvm3JrV89waUfoP64dNhPP7jm9h1PDOWf4/JUs53PHw/NdxGknHmL
hFkTXvWAfKccCoMVul4BembcppXzHsCrvxHhtXoxT4ABSW0HrG1n4Lbw2cG7kFgRvlasUIzpQg8p
T3H4OKgq+2XUGfBleDLoxhKo9JNsQFXPiSiHYeNnRjlcrGSkYT61/bNUgcZetecDmF+zGFU/mnHL
uDoU88N9BatLIOp9e3jAGN2CZha2pmzsjo9oNBvePCjf5q2T+PMn5HA/sUAIqE/ZkjnKKNovH/iS
dlNW3LlIKtehJqLtGYrt1FIfC101CCI2gGuh5V7zGydGwMt7UoO8CGVDNT0kNJd8rjTZN+YkJAir
D1yLqa8TkajkBDsg3UlYaE1VBjv5EkkAQsezkM0h/z2L795OyATgTLhFt/R6Jo2zr60HmaJnGR8l
OYOM33eM00I9xtvPy0w2RYwoTxvpqTEe1Cm5HPsKiGvlGCK53pi3TFNSfKF3ICg2LNF16ej0CKy0
5uMele5BfF9J0LaUR4HCzbY5B117Il2MpfgMfQuNfkAdL7+W0xbhMR486FXh/cC/xEdp7ej9Jsfd
UbfrOZ2/OOC5LXYi0oXkzOh7Bv5KOQyGakVntKmRFO1z7Vc25g9jBrYMtVBoh0mQZQO2vXC5J4b8
lLSBMe83QzW4u3L7Z44QiA9il3p71IITgn03n6ftDaTUL+jCg0vAMuwxf3XL1ocs2vWLBMt8OKsl
B/Fp2FeaZWzNMe1Z6b16GcApxey3cL4Fx/KKUcGRTJ60yKc1YEXS37wwxawQvXytY10SK8FfuzRv
lBxLmmd/TCvpKF8zRSvGGocsWEe+d/MYXwo3Db3gUakf+pUELRYKqzpo8HTE35GpO9QU1byKrzg5
HNQuGk8Joe0vx6Vh4s9c0IXwrU2qKbnNtufFQTJYwBGziUvy+paeMzkfLbYqeZ/4qdJhZywFGalZ
tz0lzN0bqeDaGvJ8Og0m1iZ2iKuaIbGMMIsjAs8LRH4BOVWRtVNL5RZhTTFrFfbNIy4TV1gPfOsb
ln0gAUgqi9nqdPiEsawTW8JXNrVXcPPX8dqKyNTf0AGfAUfUQbwQSgPjg67OF5TeSv0Q1Au9yYNj
l8/CIjt01tQ9FSFt931x+FotKFakVwi1yaDbs67zdqF5NQmaR9OdwJ96dnCLdF5kfVv43Oa3VWv+
ZmxWIlMHrSw2QLoCSkkBGuPEhwROO/obw8F5SVs99yo1YHUa/0zKWMjbBE2E/tr4r7f5DEaA+aye
PZsToVNqHseK8xw33r5uDdb5cSOv0IBdjtvvAo5rbelQWLRzL0RZup8ssBKXV1A03ZZb4MueyxMN
GdK8Ixj+d+HUgbDrn00Zbd3ulKk9H4AbuIEZ65F4/6A1IVkZWb2wXAcfL3z4O4d/WGcwfln19UWz
UNHrDJHI1uoQ8u4/AaIUJObmhJB8kvnHOIu2rio1y3gQhz8/FqyRZYV82WPGpOmVjFIlTlhjHQKW
exnFtVBXYtgPTnV1gp18vleADjEEaBn0hDEOg/ZZzo4uiJszTRqJVq2D+jotaSeIONJzN4i/AJcU
eoiWp3C5Brx2hKdKiyypJi6dzeYNLYlBvHEs1Ul8q+/pwbkXQQsfFG/StOeNEcMWefXGLWusrmhc
1AbKpWGi42WC/Wiz4ZH4NxeCTynUrCVGpZkyqgPGDsrtd8zgsJ4lg2sluh3N0gpD5HbcpaZLfcna
T4dyoUJkAEkv9txPQHdileTCUtaRhXQP5rVOeHhdQBSgVrgCkrSTLRih5Sxv4BLIWTL1pGK1pSGm
iNf+cu4HSktt1gKru01LiC7RdH0SKSxFC9+gouAm/N0rLyyKQpIonDNcwB3aeiB4bmk/uqPElGb/
ZMPMtKDR3eozcAr64avZ1SRWIETNYhj3arPUO1Ys6GSWzqRF/OFRYxmVTEcPrfwHPdVFV5f83axK
F9LsvosDhx3vnrjegVZsyn5I0XktLUcbBWYjbfozdgelnUYXrTH4zJX13bd1jygLXqINsCA/TeUp
NMyMSKDVbJ5aVb5h9NjIrqOKymugAlxR4nei2t40iUVxPwOCvXnOPKA8HFgcpOyHiLvrDNNAtmJ+
iZqMUjQwaBTgT/7gE2Os8AMiscxGxrCRryYSf7PfpDVdQXDTUN4Tug31J0f2aS7mdsb8F0pMh6Cn
JYTPrH5WbnarH82GlpbYFzuciinvl0T4nL/+iQUERKF1NdOjFJqpEeSK+cUcdcQlyE5NKG0lBQKi
uGHln9zYYzEzLXKSOShXeOjJGiJioQ8kac1KIP7B2ONMkxF0B6f/4K2cHZZDV/nCDZoI5NL8sJxI
XvugoEfNINKpvGBG6kLawRGKdKW4HnxVSMzFF1C7w8eJA5e8/6nUlACtyZu6EVR63s41sbVsTi7X
L8vP197xUVqlEqOrRH9vsXTzAnV0OqZJD/eNqN4V+qXfqUYPcFl9UjfQMwYE/ucH0mCQ2T72lgbl
BubGdLGvV7NbhXQq+7kLtYUSEfprl2lpRb2YM/6rvTWO821xVzCmCbMX3WRwB7HT/dpbLXzYwsES
ACEpT2QxDfW+ncC+jV2cOq6/iq87fd6iS8EyT/h9I/b/bRGW9wsuRnrg5zWxOHVoYWeYuuib1myJ
s0Wp3g7zD1Onp0dT0s9Cg6FcdEO/NRxw1ZAOQ5xzjap+wEdlYwkfvdsnnFmFYKPvNmlbJecZ3qaF
RmTa+srnC1Y+mWyLlUGpOmqTmrQXkgTeUicmv+oDEq0zoj70TjubCE536MguovcISyPCAyAtx/ZI
Ttr4iI2vR+X7tramXO54qOYyanLVkKs7hCG/zSFNLf/pV+FvIFD11KuX2gYO75CR8fFwsv1sJK8v
xiz92wrPsi6CF2e/5HmPXUH9+WaX0tZKAeYbCO++3uIpRn9H5vLp2WNtPxFUOUevEwLZkG8ITIQe
e37zKQmNR0/YqvVugFwOtyS7/MRVMcDTGk8xpJeNJmH1jDuxOZkqq1SeDUiBDGB9ZgRRMxzIRs2l
ioPNxCRbdqN+hP0+LtGsuPn2EUbnDJtP5MCzDL/qHPnMrnjTbzDoThMdc1SJ7bmuN0966yUk1KUR
wezEVDxLQFgkqskYjwgvqwcwQWthM03x4KAoIbcCKqz3lyMermdmjTn2jogvrgN1rt+fvwBkLOOl
lXib2c2N69CwZ4SOCgQVebrX25q6+aHWfcv6YxIc7nP5l9zpiPuo8Mtc3DE2r1ps8fc13WB2mZaW
k5kTev+GsUicniVGiWvyPyNKUc37QiUkFJmhmrV4YJKdaniL9yerf3SpL6oCDEhcOnGjLH9V1Gq4
A5/MhLQktNnDOM+SohbSFf7C1taftQmucWxA9pODaiz3StWV4OMcfwE7ADCHvH81ZnPmamxW3l3x
1Q1LOv1ue7NHkHMf7laJJipXvz5iwbju3pTrE3z2fsuSDusdPwIilFZTvV7SWMlj2Nd5gWY+/7p6
2L0k5VpR5gg1yC9y43Qe5mDDyaDNj5lV4J4A+yarD3+q/G9MaBcH8u009gcMjHgOSHa+lrBf8tqA
C0pdLU/rVSMyyD6cuaQ8ZY6QZlCVMgqmcWwACoipz8TJy4Zqy2YiFA0HUu19W6UNj9vGAoGgR1Q0
RUcCa8/l4T29xW4zY8iD4w+eJBNMgATbqjR+ZMxf6YcuEIT4DjWtEZQHVCb1DlyJzz+Pd3SvA9n3
qEuIn6/dG7nXys6TfaThV7fAbgDGKdgt0P/Of0s7fizJ7N7o9BbVf8WxJEIO8f3PDWvmbzl1OAJh
wmIVXDdS8Pj3T+8EUt7rmQPr6ajqh5VBrcaZIGoYohYu55jtTgFHqYyM9907KzFMfu/qAQbXyt3A
LPwgpBjkwLcgeb8m6yCx9joPG6v6oxH8MRblXZCl+6oRxI8xjTcL5Pf6ADy3zq+3Z7VorEtvp7aY
0rHkKtzDQ+QFMUl7Yxun0Fs8m19QPqElGIB8oQDm8/JYjEumDyLeUzqLDdtmu/5ir8zMOiTOfQOn
o17eVH5v2W2I/9WBP8yEpRT02AYdlFyoPFYIqhBQr4N6PlS0p8sejrPSWVNwLI2QiwFJZsBzBrn/
XV/N5fbWuUlYy4G49sDbCiqgVNHbdAa/eLinYrgu0g/hVlHHSOxWOlJAJC1+8vS/iMpecB3L5b8X
ojFXiWkZO1oJGb6/p5LHr01rLIusqzN/eqS6BgL0FOrDtn2E1mUegsWYaxPK858WrUyQkwAQdYkN
thlLwOcZhhlwcdrIc98qiEbggBnzkJVkkKl57BFMCGGq38lfWLXF30GyNfPwo7iHCLDlUGjaFCKO
ZNyyzSHro36lCuLlja5WGNm/U53HyJwZ2b6XP1AeeXs0VexEyrK3leak+nofEC8sMaJk725Z7eKA
7j6g8QEWuLnWw2vLG3jxF6ozK1N5E5M4rrBBa+8CUGbXgxxeHb57N8CDsk6IWO37fd0Gy50qwYVJ
kUn5YDUMjH5DdKwNR8a9bqaI47Mvq3rRTcAnFMBAnW1B1kvw18BtqxF+Yu2t15o3qzYrNw5WtWO4
KV7BSjD7fDYvdI/ueDuzfwwkhXperhapRBCNm13gzPC6Xcb3IZj/K3HI06sZ8KzsTS0lesOeTo3j
ckaEcUeBzmgUEDkVGvq9hE2aYp4ktbDB+DlwnwDlmVZCXITcYYqMCChzlMf1hJDtnoW04SVgCgSN
hGxxl34lM630fTN43YC8kpKTY7vKSymbf+pXQOLdc7BxFkkohVHzkkyaiZkyKljSf9qk+zqgsknQ
JAmaSkICLmUwxhvqGpoAZMcKWcoxAmkTSb2hImFYc/8lZR/ncmBSILNCppdRMWJoQuR8GM4k4faw
hB/JfKje/uPt1IxTD0nrDADX97jH0xGiC2iXLKt9KIOI6phFy7DRpXWYVRh9wCdRiBktZg+sH5XW
jO//rsulGGlSmEDP9JWG9Ws31HMgz7VUuynDuGdDVis7iXI03tCSCpwgvuaR9dSc463TRFUtt1aj
lJ4rjkx8x+PC0R94DPAsgjUmOrj2fta91uQXlAeyE10+rUzYTXQYUfBdO/eU5t5VDW7J+ZybFjmy
7Lq/7Ki+CECJYzmEVMNvSGdEkvMOfAbpLbpv3gvzMs0n6tAHI9qDYeX4Kla5w70EVUmlP1MVRkqW
X2Z1SsqmvOvhx7TKO9bta/9efAMHnrWvHghuHePH3rIwwGymoj+Xcy+Rql3KNG37kYBB5iEhcqca
YYYaJoM5vXMLCxWb97W9lqZARM9L/TaZQWGxiQ2EVD2khi3BqSdd/cFeYcy4jlga+1CDUIRYjTCF
7uNrRAtq48zjtfvxbsW/G+qxz2Lh5vcP8KTOBEWvlJRuLWwGljrz+yusnvTW3hXDre/Cht9HCt/7
7Wq959ftL1P3wBdnfQGJAjuwuAoqLNg0lmSsetZCTtIGCcxxnDJoX08CdTwogoUraRNK1RU6zK8e
M1npUxedeGfG5pOfMSXuQdZiAa8k+LHM6Wm7RfVxcVbC+wXfos2bBeJC+yvLXMBloz21+6Pyrwve
xIivnveKkAvOUppvjLKzoB0WLobUDY6Sdfh4I1EewBCFlWYvOLEoPo3szFGjUGBE568mnXYISsFf
4zBn/0oN7qHWRM6loJ3cuAX6uPgTMx5vPM//HW7g2XU6zaQw+GrN3N1W0PfcqSjHA01eAUeQ1pDf
DyqTWseaTZTE9dEb57JIqTT3JVQcrSVhBrOefh1RxJ0hriMn6eLTTvVORtqyQa3ijqubHc15tkQL
KL6UflWP8GIqZp64qGpCKQ/wfdo7xu7J/UNTbRLydG+hHLfYJPsSHmL/ZMA/G+Azd27gLHoMXPNB
36R63zAAeEbSpj8ZbcwTOMmrMlHbm6avQhvI6sfto9sjow5B8l0rsT+tLvRwOcx8eZq0OHYB+/Y3
PYIbLCQyhJaFhaBLyCHknByqDkUa8GXycsRempDlk6cXR9rryvCr247Gjf72750fp1Xw/qn4qEle
8tdH3ldOMglpZidXMIL0O1XdS+n/v0Xu/FkzezKlVNRqzC1DTJOcTXQuY7I7mmtlTQ9qA3hKhwlg
8r0OX9t43FOwBRdFZAz9/YCZpyQeB51nv+bDi5Mmib7UT/l/NdwiwFROnxQzVDHNpE5EZtcbsgVL
8Rq5+OxvsVdG6R21zUgKSDHqdFu+eujL3puNidSqsMOv7q3Y9RH6pKysfAbOaOTlpAfzjFtzNDy+
mVhWZjn64Vdhe9FaA/v2aPsk00VhbhI+qRld1miKRZXB4cgGegIlj78h2MD3kIix6QL8u4cuIa6W
UdXTG8oauWDs2v3tBsxlMVOzrSQ3C6ADUv7KvLzRA7g7vEh8HYqAZ4m0FWHIU66PpBqrPK8pLWed
RYPjS4/PV9Ek3xKGWquizciSUrXFAUCpajblSd5i46KS7YW1FwZY236n8E5nPRgoNoH6Ic+Ay+Rm
SzQABprYV4zwdW9lVRyr6L3pqCx4DqTdBNwTn0F3haUZYpAwccKU6lT5W+JpNstdQWqKjPPawQFI
B4hvPyPJ5ov+Y/8T/+PSbewtZTC2CTPNVEhA40brtcTdkLpH7rKDtT6YWygEa3prpWsL3EmSM1+o
hiw14nWg3s3mOAtJUXB/SphC05mf/tkKSy7pwZe8+DyItpUDIXr1RTglsY7DoCHnDKHqCBPPa7IY
wmwzfw2NyNcdfc16EnVw7AQuwjQcGxxZnkpJx/jNf41f57fP5yK8MXTM+D0GJYGESXFrXOd9kbW4
oyHhZ04G4Oad/Ny5pJbJaZoCazE7Pqzdo9CmWvSvMA8PyWo6n17QnKGFTb1a2p20xBu9QoSyS8ZV
Enmqbe8dOhTBADuGXxXIBfgxh+oWupiguQ/GNPnnO/CRLbC2JK1wOJrz6aEBYzbZbnttnnVsLl3V
QO78SsstEcV/CbAen2+Sl1GoodjPeO3dL6JGsUNg6EUanF/VFp4gcxdrLztCb27zocoWWdxlvcHa
7flC/KoVcZNxkVo1lMK9Pt3faR1lFkLAtBucTBPv4gVjIk5aq1fI+UTZDEMvv1VMidEd7HBmo+4c
B2lKlBNiHTH3QPfL4IhN3ERdA8WH2uneKzj2mWDFFQHYRtqU7pEEYgXJyXaJnYz0z8shpGK/2xCA
4QdwFy+TiU+lCcjjeb1lx/YKfMcoOaACs02pzfFDolH4QE+KTy6O5DTp1i911kcrxxJ4jcaKTM8h
veq1zPUOKLYbij/vEvz1PWsfmv2FGFt3qLvjYz8cL10j8pQ686prLIyBP40FXYVKi1q7R2s2k6gE
GD/coRQ0VenAbeKRVwuVzhmS3ouM6FZd+txksVj1PLGTAE65BCpNuHPv4OUADuQR1v0F66aiz+jq
43E8T0jDj4yE7FD0NG7bAGp5YUjnwPFewikytaD1Vk+xol46AdsQWangty0pUXMnoeCmOHdNHafY
lZB6Fj/HgRoGhVAeH5EY0vTGlA8TduKj+2c8SQvnnxYjY2Nj54W5t+Y7RDXypktq8Zd5o8sewc0+
WTXXsG853J5/m+XNR5I8gSY7Q5iNOjIS4rmlTnhGr/ycAxO8jpYzE8+Q98lqoMcr7rvHxTAD4Be1
FCW+HKWFE7W7GwVWFyD3Zk5TveyzxDxVKh2tboCJBvGwd19dy2gYwN1B94nQo1+xekMQ8zO6MX3G
O5H7sh8uGj/fBYeTiGCvRDiBKiuX16uf5BxLkmDtvHcwUn05ejPRtZBmO1F/gz+F28Stleb7uJ8t
iWLCSAGi7WCTcjK9WKxRbYUuIlSnECi8qrn9xXVzy9xBTy7tisn5D57r2GSH+ApURjXks1SrDVtw
/I+moG8SEX0gAU3oE2wjMrKDQmzSROMa6T41YYjjcvihwVP8HIRX2tLNujWWL7yW8OzutDBi9T/s
StDgFHoeQ49pSCIQCNfHylndBHwofYWIL3LdwfeJuVRyzO191LKpWPdip7ryJrgEbm1VyLk9Mhov
rs2MMWpit5o6MTixVBUh/UEtzKv8jTLbasG2rdi58QJ9HgOewbSepvEuAL1gdb2JdQ6zHwpPIThr
Q1b/Xb/hzEEW0RTbqBvPHa/RWnbXSTEI82vPZKAsGS57qAp5u1ZGN6KBDmt/g1nFhdgiN6tCFlp9
6CwsOM58PQyR1Ib8tQlsYpwjjY+mPA1ajX8JJPzYEwqP5GqkwF1VyHQUclkAeKlwQCshcDepYf5Y
lXqkiJoDTv6jmj/qREwRNwL3s8r0BweQykMagkYbQrrf3eVx5AEe4b22g9xJtM4RqSKacHFzNR6W
bh4PSj/fBXlZs/8/XfoqgauFBAr0oBllSwM269kPuttx2k+KNwqw5XWqAOXU88T9fXqrR/dhfZ+L
jYHF9f+zGOwR6YI22ZsjWLy0qMTkIjcEbbdBMij1T8KHEcfd3g41edxAxEFpEsO4OwYGlCY4iBCJ
BeJ31hsZRlgqPP2fGxjcUvFt+N4bUpRgDrSMlKEHIXKNHE21nxiYg0kSkKnW5tLCTt8Q7owE60QO
zF8Eys9EXc/SijJMWlF7vwa84LElNzWEMff+gyEkgXHEES2nYU1g28G4H9bFWeceXZRaXQND+0Ko
RAY905vF7uWIb52fKIepsKX7MGHL5k6ogqbVk6IpNjan4fBKVRE1Z9+BRTodjV81uNhmFa49TwIT
B4JIPx4f7wCvA0Pb6w5GXCyNpmfnbd3deT0Rl9tvmSL/r0gW45FLfQ2ASxPCY2CVh6gWBeJYFDJK
w/8HpoInxRk5+1zO/OfTPvdsayBbKR3PnqRyw0Pue5XXI3QRMIxhn0kUgpu/JepwaJeidnyScsjN
W7W5HGcdKIUYOs33foRI8yI8//yDSWKab5p/Me7VDm3gBY/lwF9BVKI0HMqLUfwwBlKjfkmQ+ONE
xFdC8RSINbE7I3B4GsCRujDqM2I64zrLtolKWxRoGIDawkMIK7o2/9yid4ioRa6kOSEZfqt06/mL
As+q0JRek2APtc1Wsz2bAc4hKHngi1UV5fV8cpB2P5Mc0fko/BfLnIrdFezIiRlKWE+DGV+upfQK
vlmH6gc4/LcjsOo6HpJozJRj399SH5rbTFKZCb3qj4b8CYXV98FbtBy2S53DOoPttzsTueaXlwiW
WDfW+LIGqFPhQVw+Sk+0EL4OoUv50exnh63RdSsD/BZwuE5UuUYGpi3EXk4LFO3vsIIc9cRQxVYY
VUqCGWKnvDDnIsYEkIh9hsfItpm8CNfR+aTefHw+EyhC3jGZmWCuZdA0Ayw1F/KWWWSSMSDv+8sv
unQIu/LG1U9JpunFgJuBHrUh9sITILLuYWADoUQm6uFPty1bvOyNsyO0CxES5u5/trKYmks7iLPZ
VVY4uSUZ1ielz0gDHthLxc5cK5t+tlhQP7uxomZQDm8EM1qR9bpLkOXX5qIzEwWR2IsTpGIkDryu
oDlv/HF9nyIoxHepiJ9ctr/bGUoc/XHHa39GHQUuwgYDSSZgH7g1xMHXkYLV2Lw2WWz+ewOwKcb1
Pa7q9lhZb1jHiVb4nLhLu/SKMWV4yV/exRLWLMZflhWmo40drvzN+yDrj7+36EQMM/eu5mdlorVK
IOMuqBQHGCeYhKG9SP1RqIhZIoSP2xmK3DsMkaEaE04TiN7yFNL8ZsoHqJ5gUkdWjNUGI+Vr3IG6
W5mXxDakx8x/MbhHsK0FfmakxRAdZXdKww6hJnF8TjQgKMKrlnPA9CtyXXQmlc4aGDLWpyiLPrVb
AdreddaqPovPguqwBtSB0IIeClPeO+WKhQWy/r/8Je2c0KdYouFSZi8a4LqUayP5DOMOAlsZVb8Z
EJmBDQ8tavyvhTeSkknC92YUGf2AX17rKQwMebV7kaLHy/At9wLgLPaeVLEDY+bfmrzHj+9mBTC5
WNYRkyJrKAESF6S+5//eNVKBc4uvh0e6CM5Yuay8AhjAfZf4LqID4TMrS8wNoxtNd6AWjQjXQRB/
pQ+jmob6XrDfnjB08tIjZh/TBZQLNVCgIPQPTYppHb92AErUFJOXat3JIU7HhfQyYYskIvZx0XAm
jTx0WQqHQgR13iNHUhbH2vUeRJ5rJBMigKWc3XAbiF2kmVDtZc9jSgqsdJzEQzE99in26xy71Ixb
KmauF7oF1WzSkNIdT1Ibo07DNqYgHOltBKN/wUIAwJG/ReT12/4du33QO0Txf+aGjEntpkj0sMKY
eTJYrbLErnIr6scPqnH+/EJQGmahr7ek7KHgZkShLowcZKGkG4Kbq9ZWzdsaVF12fZqFLPIzzS0p
QqWtbCMlP8JsBrwN2xdrbpDV8pLWxumoSB62eP30l1qzV+cGhA073qEjDMPM9X2upS4S1EsIx3bn
bhHbs7h7LsjcTH38opmZhs3shNcyhaYm3t0pS2ImYFBHr4Dg/aJa5WiP6kiAbNR0x3qy333TFUl7
Sr70zyyUEXuDqU1okjkX49ZB8TNQtL6GZp+oOmwhv3V56xQbZVeJXf5VQXWZo/qrVx4eR01Z6tMU
5llZc4hXKsVlk9hrTLo7oSP6qHba4NnMAelgUHpvC5ul3UBwIHypGmto8vnALAUgm51cBXDyr0bN
hitgPm3L/3n6fajiVZ8TrR27X04qrcuB+xsbedA20GtyCiJO3kxvl60uvl6lZ4wp0DeuO9M/rdfx
lIKx6AFLBcNBHYD6M689TQ7RnGFBEeZ+SGOGjCIllV9oOH6gb7ET8F4Kx/JCTIAWMuPgnlwcbAHX
wZaziayOXC2PP561xRsTuLiinJXQZm/BYL1kaCWsLxrkNKMPd7MD0peAjih0TBvB9EyJSt6cxOqU
C+8iXNsaz4wRpBwDlZr2SAERpfF1AGbn70mDZpktYF2G8XNxYhHQrU3TpggxySCGyG2Pf0TaD2Pz
k3ZFHICXnzPuf23BXW4Z+D07tjQr1jpnRVAxe84Z7F7ACvflATKC/qoaOIeaYqGjRCpiqMH4Vrem
kWFlvs4biP4Gc6S46TTwuvnKEjtLxr/NfCsY5qRIcK2wjNEw8KaeCLCt9K2gzRgJtRxlmyQNxReR
FeRrLot0QxPLihQZUcs00ntJIA8TrV2nXXffsMc6X3Q2czFFsii/1nn7j+s5Hkkq7GkoYBe9lmvG
a6UbzddMwrF6KUm9wTyViD9tAsSCAzoo2lD7HFSM2/pA+0XpwPJzrNVNjsx0PkB4hok8sdZC1a3e
0R357C9ty3pI/SsimjjKqFTLmaqZEo+7VO96UxaN4qZ5tOeCTUrbcp/9lsUw7OdzG1sywOSpwNx5
mztqkai2HUdG6BSAmWjxbHRSq/1KbC44rlGYtyDQOF+6VE11KBKRsYTGHgqgSZuA7MjJmV2AoUN8
4McVZnpRvSfxUoslVJMlpZd9E+hcDSwTYYljPgCGEFoOem/A/dxEiQb0qqdZ8NKyyYa06aWsxqRa
hTJWikxbvxB4v1jFHQOY8jXrpkmHjzRwKXcJWhSaY3Gf1VzcUwmBYP6Ql9/TL899fUXehu82QYPq
aZ+5KVQXrt1ipef2E4QYaO9KKFOFR1Ogl8LNwVcUORqokBjtqu1WCO6IEVB3i+lkgTW/lnt8jKRo
33dbyed8k8AFLtBeQEW2LhxvQefUoYIhOB2x94oLq3odDGTBTq+30HwsYd1vrCCh/rOt+G36X7/4
5LclQ0LC6rlcsx85ua7JfdjdggzOztDj7XyGkIyFuqKhsmdCMiz2T/iFs1TUTbiaV7iFySbq7Xyx
XWwGy6KyIS6CWW66Hm+cmtyihh0ZqX8Xz0Ca8z/lEU2caWbjx4ksj9KtMMv8woTY3xIjgYdMSra6
iroXGJJm29GDvwYNqxNoiv2Rc/cwYcjyyQdX8ne5CTe4XV//C2QQBH8rSP0YZb6jCqqJf8bx8igB
DBODUPL9YHsRmsVnpV/2HKolfu6SwAQp9LlSfWQnj1Q51mg7NyEdUHhF17ggD0D9/3hPjO/7imLe
4loVOU2Hrom+gglNo8D1rje++B4BYrMiPvq4Jde1K9NWwqxGXTFtu0eeyCVuu5WkzS68VCA7MNBb
WCo0B9FLHZIM6U/9ePEkoszIGFIVkip86y5qCaBlb4q+m0SJBFUqnzEG4pk5Mz2R2sISLcr7h6p7
LUyI2bAqQuX/a6XCAI7p0UOW7b3EpWuUSK1fKYVp1YnKRyC/CDaS9fYYQmmIV66OgqURB/w2jfa5
7MqLbfYbT/ggsJjcdpH0ShjPQOD5l9IlKxAIR0ukOowrl+XsjnTKotQnwck24iGPy+SLlt4imzgx
ET4CrMxCYak5q0+yy/X9MmouDJF1w3ywUe2+kznN50C4KzAiSwktUoqFzPMrf+Cx95ySwYJxOOCH
8YgPrwjDlfFjc6An6XdOVyoj2au7icvrz8Sf32gLQICSQbviUmphdNaEkP1uIY3vwpa4qo9sQNga
41O/CRiSYi9Dlc3zwu0rGfvL20jeDYI55tiJ9qELoXEN3P3qh9tDnUtkT9gXqPxGVTMj/4LDsZln
ZxczdpCT/P+v+Hiab2mwJLJNSyvPOBAe9CEnOt5+qgQnkQVNzvDlZkPuJNKNn71zgrsvJurjCGtu
qiDRWvnkAUvw9WVBWhTW3S2aZfYIzci0ZWEFqTpLfRhNvrWRyBlByanD7gyfj1b4C8/7RXjVgDPa
psP+Tt9X1mi/AqwOKIQswSJG0eOoE4QiqkKPgrH5HUoDolMhylkp8R5l7ZJyTXs+h5EE/HNjVNpK
TDm0heGMmgQJ7S3VqP08ncnhLA3LUbi02uYnFwsDJ4CzNScbh8SQOTWf5lUiEzW0XDz7kCpItGaY
R8EFNb2R5XEXuRbXIr/rlj1iVLYV4U88FsFELaU34n7MsZMiksIZPGEuAgb8Y8MQJDrDi6o10umJ
T+8RK9Mh+fS0Q47GQSj/CAjkTgIPwVRZx4ZYjFjCvA4HW4UJ955sqy+MvuovEkLY6q+bTeBjjJyp
InNR1r7BQfIHjEt4FzTE9jEekRJPrgiY94T57gz0uC+0ydUcfv0EWWcO5MZU6U1NJhGJtISEloBR
7Wei+S9QAvpDGKfm0CwhNb/ykxJqIUFS3pl9OZi/0K5Tuxa5E+awAn4ME4HUxWdrdtnl/q1dO7zA
ZOET0/PkBezv1DJZBY0trkpCZtWDMtUcVtnrpToSl5HyhqGgXdtmvJCk4R38P8n8yy36jo/SUx5a
0bmYbzMPOyXU64vEHJ3dU8f9LvJYoeU4sKp8ZTQGD4Xu/svtGaL0m0y+t+JnzCx9PUncdaepgqwH
jPT9s3LRnsYoswHpvna6Hg5NfqFLY9q41OeybLH4onGurzch0bflBYPwxWkXk5IjtDpm14C9V2ZB
JL08iytCga0Imrlog67MQHXY08v0NEjSwvgtnMymqangMLVd9Iz1XPHEYWsQt4iuVadztvOGSDpG
S+ZN5VoDzw1fz1B1jGSavH7GiVqX4xZfkUKKlpZXiXWOQnD/kzR5oub6/ssMG9QHk3/eSgBBhb7Y
wUT78RJ6VGMp7XOx7SBazVZfwuzW0QXu7YsnO80XiLMqP2oKRQ85AFr4DzCwbu010LawQToklHpm
9dN9kzBInJ3Vr0EwL/4Swk2fub3jhbVL5C1jjnIX5WBW9nTmeltwPmRprCer5ZP85JCyVGfoSlAK
en6dwouBQ/LHpT0J8j6Ghyd/2bAbdASMEZlQMwAmNLwkp0k7vhe0KrDRtzNF0IgUP9w7GlMK2zM7
X3arh00mZG/AVK2BnZ3eStX+eeUmr4iVpnpcyC2NFD2sV4KxGNkQD8H0JJGn2P3BOfnrcI8WoRpa
TLCeUS+3WFutpWjy3DHeymvkZRfEuDG0UyckGEeYsa8ipYIHIJ5RrlHsWdnYVUwK8evapCD+3nJc
r6qmFXPMdn7TSR4XvZPGpOsC3UEmr+aFfxkfds4HfQXrmDDM1zwHdNI4WMh0ONOVa8SQErczVf8u
aZ4yc4EogffKvN7ybFN6FI2YNALtpUtogvSXRvCd3QNrcmvprCCkPvi+fCdb0FgZFF6+NFIAAAt9
DaTtzYTd5k/CzRuST4CH/Gt0dIvI7zHvCBLhGVsZybNFil3cSFB+eeYK4Kmi0QP1Wldow1FTXlpJ
ji8zJj7nzEl/pfuvm+llkNid9617N4csnxx4WhWFogsXC1rYeyHs5nRKjHQFa1qJnge7Gt7IY9PR
ILELa0XzZL2i3K6XJYVjcOFHoE0i4OYM3uzKljOImB+EnPI3c3WT9ML0Egeduo6849sQ+fWuocjA
IFU60HW2EsQ+OsGckqL9/T6gRhZQszzHNmwuAEfAa9hfrKEVAfQvn3JZI/UK2b6+OtJfPG+t+YCV
HcnGK2CQbD0f0bUaokbKybH2d95zIqrCuSd0NnhjGnAc9VdsXycIEI41iL9C/dzv9Poz+YKICKaP
kAnKwyQfDjGfh520GkY/PCF+2VjTQ4IHptA8syJr9nl+ETqZzYX9w59065ru2G15E/HihQOejgDo
QUukYTpMIWz8MLI3Fiqfymseua4Mg/I+T2djrC71ZBxHfPjuO/jh4EJ9FaT3nsCOrilEukEJSbre
QLrDlqNJ6hAu1hK9w/e1XOZXTbh9ATM5IE8zXriR/viXnVua5CnwcT17ZVTGfBOP24AdUhYSrMh1
2bwIoxtdAQ7GB+sHhHL3uBVJlP+RD7FHw1tcdAUfrf0/9Fv0A+xIzA5GwG5sC2YsgZuedC4OMGsP
I3ZnKNYfgQNJujhIYNPuthLm+3wavYfysQmbtV4ynbJyQJCUKlRwIJUtRp6wM71vC7UWCbRjbK/G
FZwEs4W8w1WfRDbQOIElW/4+f6gC3ns5BwIO62sDgZ8yb9q3SQXGzqZZfdqCQ/7SCpIsz1Iu+dUs
1OIQkBIeDbsAWgm5iSade7ZNUdLe884WyaC62RmiWBwW3v+tSE7GcvvPtbVuE4zQSFXxv7DiDzqT
rqmZ05LgETG6n/Utp4Hl2Rtiyc7bmk8Ndodm/vMUHK0xJK9u8Qnp4s/6G0pzU+sP7Jv5hGdbb1B8
rhvDcZImE5/IrSgcd/a/dQ0uGlvX/oD8YGi63EE31b9hAHel646q3RG8Kf6nzUAzUMZrjmSYuesf
9w1fK0+jJKCKPG7+0V5qcfOkPtD13RuQo9EBk/dCEFbv/OL0PsQmlB1DVN0pRuq5WlpnMYN45lqY
XaFapHEJNmOgFl8CUw19SHzmUbFa/WE+9h95RiTg+ZCipmfXKdNrw71xb5WwdQzxh4ZGocd4/N5H
jGdWm//vIFHxdZ2tfAzq7PgWtdZiqBoH/q9sVdld7tJANYxSeF+wBpaKXPIQwG4AxJD00FVcvQBF
dxO6/CSILSyHiNIONQWu/AjY7Bae1oT/z9+X46bB8XsW/miTOkOUmCPq5YCaDjdG6Ei5cDvG7EMR
j+nt1hqbOX+LWBRnX5zVBMgqEQM/a1otXXwJ7zzHNPt0QCwtLdv10HLWVi4B3LefoCixqe0aD4mT
Udb9QoGb+KWSiHd/Ju+DjnZoe44ZT47Js3gM/lY3T69GrGvM57O91vxg4N+qIDnJSm2MSSqmxXqc
S/4YaO5gmlorKWsS+AVsP1/9n17nWnQtAeu0fVvV81M0Z0Uo7gRwMcSINW5LBL6c7iE4xpLdIfGP
PuHmWCrsV8caVfHMGJVdQFA6lApVc+moMiUZic80BIl/XhG1SY5tVbg0QB3KWp9R6Vb3lNomDC3R
lSSAt1CBPkO6wpl6BE2QJBnazwBPYcScxzn8KA7TplXpOIFg4eZjA4aDiDLpWgYD/ZKMgbrFKJS7
X2cuyyrcTXlSEvEozPyHo+fDLDEprOIJ3Ao1sJ2v3QrKYOmxEZW/n+umFJElHtdlYGhT5n8Fu3Ag
/UmyETV++mK+rZojEcHzOjfg7v1wctxq5/Evjbh0FGtjTOnj94hTCBWbSUTWHyZLRQ7U5zKOeJNC
I5gVtNGDiO7bIk507tEWorXqYBLoC+IWdYm/ougwyS9mgDDTA5CVCu+8RZwo/PeljN1ttklu0WL8
JVmAVxVFaWWKvgIE/2ZNfAnBqMpmCd4I7bOUpkIf5FfMip8TxPaLPX4TKs5EGCVN4eWjAFBlfs4+
tkeKPBoB9aQeoL0JvuYAaise/Tiy0o+R7ziGfvIVSuLT6/P1GuBu/iPdnhziJO8u33qV8+ra1JsO
Fj/bIZoVqJlO0JtkazwPboqm8bhLm90W1Lb5H5S0s8Mg8Wi0CwvBlUldzvl2MN/+e/8LRqzp7UEz
1FxOMinrc0ygp+HjOAe4Yv50Myivpsywkhl0/kQOuJCBcO9FGWJFN0DNXD8C/5zsTcOg/A47vUpF
HH3uemO8HNF9QiuTJE9hS4PAjL3nxlosxdySvIZv1afQOSGMU3sqxmmHql1zrhCNmEbjuOexZ0JG
N4MY+nnxATk7k3Jr0Fz220NyU/8DyFPYqssIlrvnhDCwIvFA1XHcsLeUXiqj0BbPqC6gNGP+IT5u
Z0VN0bbrRvXOTV1PneIQ0IgjuzwjSYXtHPiIHodCem+zQRoBLF61HydL8tboaBC9aulZ0TdwILPG
4WeyWUVr1I7wve1OFrPfk7OtbeQ9zdDjzBZWlpnlkOJ6dSXdni8UUl2zhiPIWq8uCiBewl18rnos
cM6Tib6Nk1sInrc3sqIgsDUoXFZtM3XqlJbbVjUwhPGjoinjjZLBY4bAliwBg8FZ2BfI2YFtrCDv
UdtCnX+0Br3v8Rb9DzfJPmyQ5hzD5t9psbsmnbYtdXUGmFxoj7FPB3+TjRYw+u5nb9GsQX4RUPrP
w6NOovvEg5o/8xP2iP3pQRjs7DhQQnyKpQVMyOKYXS7vYTPdQGZwjROLCAQSfLnQ+IZQQ0+Zao8L
4LVmyDs6lQ5NhR6O3tZjlyeoduFxyHgRE9kb+rlYEFetE0ltMqEasL6p6oNKbIhHeUU1F0OnCryN
NdTx/4PmJOj/Iylh3J8J4ptldkwndI2xxcsjRcZubSS6x4KGiExbWStH+4EtOt2Lg23szERRGEVE
qaqR3ejMWmxwJ836Tqww5uXxrwd3gdU+ametIgF6IE8gfzRww5UWZ5Z3M1BlyyFf1GiLRBHmDqqq
hABmvyOl6bFxFFn6FdXo2SMkVSp4ZiCljk5mUvoKUHIIVMYlPR0AuOQHu/IBEkKiHglIDSegw85/
zJdPMSG/1+hrof+tFew9o0WfUkT2y7XQC0zfYc9/75ATW4NhyO3J8G8+v8h2Gx43vgxpDC1PTDDK
6rx3RfjCQNMD1BMWoxfmeLWn3ecaWHLLtt85JOcAwqixGh17GM9PudrWtUSMOfIG9SEkqJudpzg6
gqrENmIHNa/Te/bIIPul/UY2DHQefa5GMtaf1Eo/GvUvahf5oRoU4WyOYItQRQhBBNGUatVeOtuI
LfAiC319TXhH+iOBCl7qS4KIPGrjoZLr9pFV48AY81YXMIrNFVr3TpGBDPyChgIwMCHUuIAk/9gw
eByUkSY+1ThHU5NNmmXvMbs30Q/UyDpr8rD0/UPDn/Wr1c9eUnIxL75hr9i61Sjd3CpxVoLQKDGL
+WRp67TeBAqHYwIeiHO6Vn3ipKPh665zHlvapVO93RCWOlWndu/oQI16ugUmVbu7PsX9TvP6C2a9
5FqkrDJJCXPkyVbqVUvzWYh+oPtX4zQnDf5DtuPurGnro8viJJ8ED/wy+W/ij8Hg229HTPbN2y/h
+mSbFX4yTaxP1ayRbzxiLBYC8p4mDlk1ND4aTUNNl6XZYcTMPZtc/yzuerIWtCGRx+amQ/vxEjBw
tJWha45ZctL3p8hBBYkvQEmz4T1X3iMiHOIjI/O3uFK7ZtHr68k9hObWT9O9Ip/z+hRPwTa5aGhD
0jcOvbBBCvyjP8XoHzSvrtjTiaTNOUAVsYOy2H9yrTiQwfAB5EnXk/f5TRjgbY/eJjGu+8Ffe1tM
4uXSd03aF+MKrY5EnwPxW+EPIPHzxNz4+fAHMhvC5ReUejFonTs2GjEnhNye/oO4uDVouF9mtHpI
yzQr0OtQSQKialEOM6Jf4mY7ZzqhXY5HQkQi9Dh7HYZX95TUkLYVShDnYqq8tfaxVwOrw7Kv1bBF
dv97gpeXk/ExP8rCD0tHNo7HK12+HhoHAJhX0khNDq4J3aOnIiUCta7pW/HQ0JjPem43kZF/dKb5
n2+nOKWRld0IlMZBccwPiRX4eDhKh1r1pfDWBKeuWnCeBGD8nMYkysirxKarwROZVwybjLSVXbD3
VkRX6YHWIYqz2qf9fcHI+9x3Vh/wlK6LhLdnrfCb/6P+RlgFKZV5iBJv6YjShGe5T3Xee0f0xF6a
ImAeC/UgrHreHO1RthJEZYtdpTa5tLQc0zjF/4C8c5p3/PrbksedCoC6F1t7IJ/G5+98Qi+7gRJh
y/wT3FyAY/zZlWGQTrHc3IF1lTqtOWwrDLmowOpchXUXARuOxDijK10OpjMkRSKw4zGNfbdeX5TE
luq+9Nqb+bVl2ifk7WRE1f1rUHkzYL9c89uLghG03cOyjI2a4e+JCxWLVlLeZpL9StGSyphaN6kE
0gSh4cksJ/nRZE0YDD50xyer9QrWxespqjnImcLXE7rkLVYawAcYQsWeMcbMf1USCH8kmRSfQroi
WvSHEMWgVMIz5cgkr7Qc3gwl2JOV+kYDlP7J0eGv/2BcFzRLwvlqi2WxL1E41lQDBur/pJxfdhtw
4GQ4dZ0EsGi5S/sSu1+BxjHfpgySDOYeLu7TzWgQZIEOLs89XjdaNcaCeMlBdSRkNrvGYrGFRGWX
H066mYpdfuNZJjPxNoCZaiMxVExFpjgSwb8i5pCBVFOa3JVrtkg5cEybMC5P97o2KucExQJsSsYI
mGB8GRO55Uc5w55DdLLOB56cTTX1MSUzJssSvG3nZBUqFK3vxzaAxLwvxtXYoSBjuFIxfnDZCc6P
12C5/lwBqOL0P4iByhPVjUPBWb5Y/J0fdp3LstoUrP4JW0Hxauwap1gTMH6xSTk41W9Ljti5fNR/
yeZ4Fr/MZd6Ii0o3PBwHqV13b9l8Sg4LQPKdn+1mJv+E6cEf68zY9h9ryi3ITc4sa0hOcvDUJobt
MzwOxAokcrxEtb5JeFQ0fpOvYVgD5MMaJ4hNF6r4VsQnvck0zxovwCipuu+dlNMy2AM1LTCBfwmr
MsYu4ZQWVd0BbnB979oYb/AebRB1jdHh9KQgoY7+RHztgXjswCxDBDZqoRuNQemLoWBhqNR2YKMw
+FAjhxYP6ffzIRy/Ook+HRDm1AgqAfpdsciYlqqNrBjLCngy8Ce7PrsqXE5HWbbUAmOLm2RIO8/U
P6ehiFX3yVKC5cx9xtU2+mDI5v0fEkvcZxRlac15gRDacxe1rfEI+jr7vpvIDoqKQrcAw4HVqOnu
5Fht8BNch8MFzUxa3kbByoWfh9s5ca4AilW38qPgmlIqiam0r+0tTAPHol5BSrbBImetnnEEYbd/
E09FUXxBMOMFo1iqbx6qggR72ht9DjYVWbF4UB4ontmwRAvgAc42IT4bav3vGKGu5jKJLMw9Nmdm
M30X5gXozTbUOLVbWKWlgS6bqkeX7K/TtIMgmlvyhGcqOECkQ4IJC9NC/X+P+tJ3rS88fxaDO62d
DmZ7kbmBCXAbyvasnP4hz8678htjK7Jd/3JpVeME8ThUy6BBmXABdRtcsBqQvjeAxUeYFuN3j8yi
slmm7cOguzuiBz8Qba7HGuEbtHQjQvfVFnumISqff0LJii4kU2ekCJu0tKHZHQEbQo32G9dftJju
vCfIpL6hmL4Gg1K7lA6FNogTiTm9xr1TX3/TN0dJ1ewFnlvfTfpdtZwBWnnTs81fUdjHvTgdxGNz
FwUTCka96HS4hp5wxOg2jA7HVgYgo3s2pLEPEPctN+F9J8yZAwdyrti2LiLmN9NxaArlfplmJZ0q
ud75825tlfmkSzTHzFm3R9Iz9gfiy7/p8qH01zsyYUhSwjxSVEdBYsjXmKdlefBFQEBgk9h2gUE2
8w8wxE0EaZMe+I8XR96H8JBFjys/MHmEWl8/ZL4s0sgN8z9oW0dvnDDsek6h82D04RxVgW165A9i
EIZAk13kP0gZDE7zb9oQd/Q+ZvrJu5VeL0IzrC4oFc6CJKIdzLxmJXwLB3xgcgvqVuFYZVYMktFp
I2Lkdf54D48JCads5XfeSzOT7cRxNSSkKc6O864LfMx76+LjPcdmZ0x4L5C1O/QCE3htUXmWJgtx
VigRzgjBDCwPrw+1kHgMjkx4d28G69+GNcX0LCAzPySFUlY4kc5g0FsYz/oknKd/BPOhCuPwXPhj
uFfYe+sUAjKrJuGOWN0q/T8D63ZRZ3HxykQaV3Wvh5J3GXAWT9+GFsnWROD0ysI1Gd/ZBiysb0S8
cYvneokcL4nRs44PBQ5/M8l/Ju12Hzz7QZDTjEIqc4kuMJj60YEYdQbHQnKbqyaKKV8y+Mfz/Pts
rdIYi1H/kM8taW6niQRX/oj8Nf/KycqDcVJxseag/tE9MtJRLiIduFyOyEMrycW1cg3sT++rckfJ
NCyXS0ByTvoygGtCPzsN6G11GLwmJwPzYYw81TSvDCzVGnmg5B2NTp99TMQBT3+LNtpII1FL+lZP
oUPpnEt3ziKI4GoyK7iCZm/czeEJBRlMZNdQzCQiag/Rkg6E2SBz0cBTIbHFxo6o+C5FtL51hB0E
yPlEQCF7ybSJyHAnWNnBVuO4Q7ND2TCmc7/8p4xOv7joYNjxvtKHb+/w5pNOWSC6D0fW7g12Kp1E
ejJ2Onf97YdVbrtQ/60cazMS0TfSYB6w1iiWo6TU3Y3hgTpBHpm/rrjn3+lL1Qrh1NexKGUZYmSy
VlKw1JEkktv1HIdQ1wqnAn1R/2J1gcbH0EXyPzsJMxGvLV3o7MoAqYvtDyy9/bvad20zAlHtqZ3j
tpHVi9e/anONdDFjolTZ3buVL8Peett3zaTp0o8qIsLTARedbVcaLUmvinaca+EsuCUg2Cum9vAE
489afRn4cNCOO5TNrpysj0eUDEEqradlI0AWhFD8yzl0z7Pcv69Sb/mUqQi6GZtk8rLw5xf8M3mB
w5p9vUsbk/jypR+P3Zt4b0SIhkGTbMeuAhcul9dD0jM1/S1Gke0MY+XPuuv8aUcXbal/e88JOzsS
d3DGRUohwckrt7VwGWM1i5lb3H1cF7zthjxys7QuqBORvyexlhfRwaJ4ZKZ1TqT/QApvvP8ZPGG+
3Yw57e4FXkYP2otq9Mja9BUAZ4fWJ2vnyws4VxQd3TfvKek50y/nXrl34LX/cyw5MrgzhBnTixO3
oUDo5juHxjBmjYIthWw7o8IeSMjKJ9DMnM5NgRYMkE6JqDvlH4GfBz/n8dntfKtePHWmsEgkaMU0
jHqZOxxYkfTJwIBLxeEO9K29OwK0Z5xHgbp0ecBzRTfTucRtJi7CO1ovYE9AoTIRZu33u7dTASCz
/11cPzqe4EBkXskSu2tP5+MO8N1wrEYKmeCv/sXltm5DoK7b6EPhVVHjElHnr89LSSCRtpNofQP9
6ZTQn98Oqp2JvoInTTWspCdmv0KCkDcyX+Q52XFrk9yzb6QZ5vFPlrRiG1Oy60SIGkJcu4wPDoqK
nshCWRibAOUr2bWWR+aXNN1MSooGeGCU9M+bJSj1jQJ88p2sBBKV1lFU9kNQpqCWcCSaX1Y4bluH
1IoUSXo6FutlvGrUrjU4o8pm9QigQZYfOjaoZ1kfOjW3NlukFPBuCk7WDxve05bMzZCf+Fq3AzwR
H9Ipci+8Et7ebhIqKQ9fmpHY4fYnOLBMZD19ryCGYj2gWHrMv+dt/q5MSlVNA3Fj22KfrG/sicJl
ZqAgjJXfuxGXuz5rbVx06zo5534g7uNDGxfmmFfqPeWpMLfq7X85m2HwQYgrT8CTh73051jDUGZj
/lvp7Xm35BjLT1lQMWhA4ZWyNVrJf5nIduEVg8C4jrdvtDvFrUQnS/4rPL7JSK736NoNwT8ERuTp
RHtdeqEr66QPgDmONiy0l6RAnnIbnOMooCBU+229R/0cv5rSGMbutoT3bP6pWEXBfzpnQNK7dZfa
AAwXw29PNduNK7sJvYit4zwp8KDHrzQSgVXuMZKW1XZXttLiPPYSqHSITm+X6DyEPDxAbMzKz3db
LAqXC7lw33ttnSBiEmFPx1uUpzNG2ZMQm1eJs4UKhCNHtKCIT2htzEpPsNNthiP1ejOCJSTUvghm
VxvY4/FYNOIbe+yU9HdFheMVP0HD9YkEuIg00NWvYH+R32zMJGSxZmNI30wjWbFKi23F7ClFQZhG
jPTWewG9pJ1lA7lnifhlagw7ZEscBzwH+F8HbnxJMaw78nnLy4mhkoyYj58VBHsotY4q0dOwlIhZ
x8OYP2YBbWnMIocMKqyrYdyavtwLSao/VByzE00OayhxDFpLmSV88yscidoZdkUvFUKuCU3h5wt4
xqFlUBPCl/JVVsyy6RBF14Bl6JkbtB+s7dgnI3qAzVJK1hBp5ZM9Eyh/MnSgJTca2W2uemZCIXYz
Bj+6pjDzgFXoh3/TXx4e3JqJxpXAh7MAkv9Vo9rytgM4ITmJ/40QZGP3u0kOXkqTxL9JixhGEYkE
nXxH84WQs6zmzwKozYwg+yX0+wHhNobq4NXNzJB3/UtMXZ9Y78o/VKqAzc7AR6ncUNkcWpOStc+u
zXyidSkMoKR0DfHhU5XpTuRYkPDYbpsd5QVBgq1ijIAPcsyScEJjROC39mUbwOrO7/A4vAuLJKAL
Xi5rddjneD5WKlLi0AR1ZmUyfhqCJx0tJg1EfekH0z8cLZLCxtpQvLj7sa3XsWvV0w91Q2ZNJHKm
aY2PfxtC8Eh9qaK0Rw9xv4Q386mICOYKwWjIJC8Rdn47NkENCao4X3Q9Eq7QRaIQBx1F/4ZaxulC
dZgPFtDbwt+eYNQ1qkalndbF6TgS29OmC2EmDCu5v01D5eV3fjjT4JM5K5obG16kO3aDJmbivVW+
6Ag0/L0V3CI2Hap0aKZoi1iGsKoftHTmhYEriw5LSCDONN+XTn8VHcGHU/CUTUzXMtSREKlzHCK8
5oaM5bowv9uHQlnBAFDcxikEgZGFvrXlQmyYC/FZ/pKgMepjW/U2Cs6CNboddyUM8ernjRw6jorn
Xcp6bjJK1vOhPjbLuBxqz97iRwMZ0468+o5KbXRFWSo8O3cOUmsqeYaYUn+pWh9vkIoks2LaunEZ
Clbx6tW6HmcabU3+FAifOM4FWg8jWh0PgFAGSUUZj5AFhJtMlpETEURBDGedtu71kyU72APzH6yI
3iUf5Bxonytpx1bXH+T2RlOxirf27jVhybQ2Gg6feOFv7X+f5F9VOCNh4IDePbMYVBJa4zsayTG/
eeDHfpsaqV/ikE8SqLeA7CMh2sBfp3qm2rYCbdywKSoOQAwfBL75RQ0B3thD6PiEBT8GJtFCKXhL
1T9ssFFWLoPHizehElq0WjRfaD8ChoLb8t7EsLoWHvuE9gcwuvqYdVIgjjzJiEpcuKWnYIMkyqWs
CHKpmg+c8NVEm+NJ9f/M6+6E2Ci1M5Okh5w0LnZvdb/JI5LfbbSD5RPerc66wViF/FgYvxVuAFrR
ic0yyLmS9bb+iVEHknJIAmJUguhhSF2cpEF1jMcPZ32pjIw5fxTeLyHYe1P2HK3/qZpEyfHE4LQZ
N9CEOkU1UjQvgAnG8H80KcHTy9TvwZVH7kDDx7pUDeInB+x3s9LVo0wvMmburjDJ3UYKSZLH6AAp
NmIICVyw7VAO8eUG7OWiVhM5+mtnPXT0/yw3FvSSn5+FTAK2jxQ5EAQwZ7azk3Ag4dVocuhKpftU
MuGCcfBNSS5h+TiZvzblho/IfvsVTn2IM1YoEMl0Fo1fjyo/5SnOaMe5iAVLJdWCrI1O9W+CwvMI
LMUKpeGRUKVUU52hmXs+TlnX6InKaBdnh/TkIRNYA0TTxjlhWEB5VnwoMgfloNwGJa4I9Nw2hUzQ
vUtIMkYSRLMozwtaMdB6E/Y8NiyDdFCH2DOs6rG0MYkfsPfWAc5m2DQiDmp5Y03Cj/U6+hVwNg0l
6JPV294R3MTSQG0/rvYpoOF922Q0+nerb3eAFX5BO86QrkBHmndFcrXOrzUQHZBVQHgISNs76BjT
kP3gVnz2THPPCYACe1Cv8mUWTenQeYqE6ee/8Z//7KLlaLd8YKf0mR1KaX1myXXOogae2jh1riHB
8k4rex6AY1NEDCIayP/1NSEgBWUM+nnh8EH7qpuB8HKia2tx0Uh7a4eX1u9oqfOGkCVkh8TTQwSw
s/mB15uN7WC6F10o4LuklYp9NM0BtODJhKgQ7gpoNYPIbv5yMqVYW1eLQ5ZLlkRyUK2MN8v6LiVi
IARtQZ91fq1bPxraVUhjUxB6gpIwbPjWsntM3f+ICtdZTFlqzqHF50vRom+VZE2+nsIzw1fwM5HS
k8rXZAMB+P0fV4qJ7I28z9OzRJqJtpCd65pVEyDeODKeBA591deBFFYmSHlTmGNy6LHoHdIv3M1T
yw9mJbxw8GmzfING77sM0YjYk9froyASJc3QI8CHy574ypezofaA+okN8ow0chuLIGAaY0/aFgXQ
wsPHGSCirAC9hGCigwkBWeeG3tL1axL+VX/hVHmZVYEua+IhhNLtDH1UUNvjJdi2N9vORlIMTV+Q
KC2RXldDkDHhTtNOoxEOnEGvx3CiqSQWsv/FqvY0H4BEZDHT1zNICXFCVIQFRm+rRgJPqo/eJ++3
HnBIQTn2XPf7MX2enCzKgrO7RfqpLb/ZsMM0uO5D8j1QaNaiGu9uuWu7LzvEHWsAsNR6qUvRDyOQ
BK1wrW09tdVmCWgpX7YVQoRo7KtAVn2gzvCYZ+nAL0g49unOAh8NRxAREba4ibT/4KASbGzWuCAq
XJ4+rN+ge4+VycEC4ETKkkqEXet6hvn2KUJC5hFk3lSU5ZoTOH38C8YPvCXNVPKVKVu+RfT1S9GS
ShMyxyzxHWp6PhnoDlkhpst8lZJp9Rl9GS4JxBZy3eH5XEwhkOCIBDSddAw6N/Vt6DqRJe+dpuJ4
pQJ/wHitjix2PsyC9ZcxjXPYxSxjykqbdUXLvVYJl6PU7nax+VkS8+ZxsBu/8UzxuHK38vfpimSa
560tudAdHi6qaZMQ6on1OBsMtuz/2Wuw8+HqmhCIGqlDCr7pcXdPetnkWCHoPeuqHD90U6Rk0oFm
xfL+gwChUNRLMXhJ0fpJ8hTMtl5dS9Gu1imaH5Ri3PbXtXLUwm9vj/U9NnBL9FVEPrGAxvaeD0S6
2l4ZsPAK3Hxr2l07vWNViaGUIyIEY1hZdacJg5lnSXlBvfBpSj7cANsRiQCNwMgBAGfAQbUKJsHg
PU4m2ySy4Fg425VcIDxMuwJNCzkwa9emb10B8P/+HgybQ8bTMCOsymFAGi2vmbyFOeqSmyZkAxIy
SG1dqGVeEQhQrWSABnSw1RSnEVdpHQDPQnbsh9IySUMfi/z8CS4p4jACIjRpJKmoBVzqWhhQPZCL
y2hNJQ4BgDccCahdUmfi3XigJBLnIbTV7YcKHLi+wm2NvNKGQk99kAhNMT//L4uysV5KEDwlq57K
T7Se+GnTbhlvaqt5byNa11yyn7dhxvcxpPIEF9UORkOOthBFW432KM9yWlWqjoVYFSoShJHmW99q
9+omrr6udv5HTEP0ofMVhqlA5y7HFVBmSwp6XdMQ9gRLLi1XK1OtdP3Gjlb6mIf2qCT3zGa1SHJW
tkCh8JtA7qC1AbvjBf2mlTdkjM0dPmWtuDDRD/CFa4vKKd+hPTlgd9fsQN5sX7e9hCWTqzxwvr3R
lFV6hLBb2KLZxMYLLm4UsWobGOZzXrJVvVWCyhaaiF9tgu2/EjpES12gY70YP/PpByT6tvSoHakM
iFrkymHbNmcnchZii8zleHvE1F5XRKEIowUXCfP67HLnsxZPWXXoMJHRPYe77JiHFhyhG2g8PCm8
Ysk3A8JxGLcvYoXj6Bd35n9oPreJ/nXSh5ESpKK7M+2eQ+ggNGkTD3F4sVkSCZlN+8DVQ1bYrde9
jjHFOKiQ5NGVkUoWizqioan+zKscNmUU4m9OcrDEV+QXX+FWsvagcbk7e2bXlbfwolQXCT4Fr5QL
05poQBZbZVYY5sVVaceQ9O0rPaCiGkf3IN1efWtqLnP+MKDT+uOEHsD+QS7f1IX7ErM5VpieGsSF
xxxVYkqVhVdNltC0xaYq4H3HSdP7frw/wiyMJj61fZVbKzXI76m6b8ywbRr1NoRdPugLk+w6TG/B
x6VtSHuzgzbfIWkJQX1Mg2mPiDwkRcsY1yAj5wcYuAlhLZwxVKap3C9kBr8Dng8npoSmGQ6zm2zR
vAJl2gLAC+e6+R6cbj5AICr+Kbsr1B/AaEofcuLmajRvJ523AUYnY2bXF+wmxZBnaXL/n0POU8bZ
hqAbntlrp0W8DC4zNqnOq3LtVQlMxC3ZZ6pxsFq2yCJw+Mjaci+9CVI0FP22wPAYfUCyIF89vxla
GtBvA3jYzcBoLQIw5Z/qE2I01EykGkMzx6a8F6KnPid+sla36mQaLjAXAhyalUhnZkLS69GjLa1P
Gx49bu63HXiKG1VdIQd65rlpQ29VI4loY+Ln7vG5/RGf6qnOXc9HmRHOFi0ClOzYq/bg5+N5UcKN
cVScbDoftoh3RiZQnXyANir8eRG2IKREIPM55Ft4IF+1CTCJ3cHPpvdCiMgR4rI9XEAZ9xdgQGBA
AGporFEKcHBddWdpMWqXqFCI7AWaIbV4x/dLhXGWrPQQ1rNMuLfokCMFvtpA+fhVge7NvW5nSkfd
mx6s2RdnTplBrWNJE6auQKZ0+i16aAusLxj1wJ4gUMZWOXVTsWFK3nvjceWFFxhJnlYXa2khrs18
8saGfzrMCIfEDl0Kop08hxZV6LHdlirwuyWD+BydumyGMXUXyfRuXLgkSdxLaxPsktF6K7Sl6J23
CRvlaVm73cDIXmlHTwqtNVBFTa46Zw7FF5vD2v3+ozmPWip/6HtHWtbbuu6vFCqaSqAssuSPkxFp
ZSRr7qGRs3FDs0nJ786HSadrKu25vk78lwzyoOM2xvByzwTcOeB88Kd4PqjH9E4iISnrgNa+Kjrv
hZACEDjPoAYaz15A1sP1uPYAOzTLlX14bo367MIeSWf6CiwA69Lik+pSusKoztaenIJnPe0ZMTF1
Uvzx48ID3PUtztXtFYM/N27FU61Vh+THMdiwEX48PrISkuLz08n0VS9Q2/rREJt1O9Fj2dhZ0Aao
LMBZnCwhipYCoVtb5SFrQ0lTFw58BoPw0Xz7nm3YhLdeXoQfHdcnvmTp7r0+FnDygsBLSe+YLRO+
7KygyYPIeZRfC83kpDyMPZUEKDkwr8ofA+p11Mo6V9Pk0YQss6P8uYwN4STuuRgXNQVHyHDdITkG
5p+Z03SzinYy73YqM0g6SQjxjYsSs2F1ggnWGmhiTWgkfeK0PI/GaCynMiBGbPK2jExt8BVDibf6
Sj18RTL98nPiUjHmZubm/Pn7eV/LzbKx0t0wpP951Ja5MptE0GPVgaKF0fiLpjrxkeouoRf0v4i+
8fFVio8CPveD5wopWGncj35lTdNfDcSixVTqWC85irPJDBYAHqO/d5+ZVsbbW9GoJxRRguRkJXXP
/Vjw9NT4FGRMhZWIean5QTFuROEOmGnn/hFSitJ1HPVAxnl998vyDJJ+LLQq4qplaJL7Wx/qa+cr
GKIQcNlRaFSUvjpywS694DOV6+vdn/92GJ8zuzKKXuS5G2Pi9RKNFDyGVrxGH/dulASzcfZvAuVX
FeAv/Mx4cFw5a+BBetk6VCMksGMpxMIKm9I9nrx1iHjGfqjoj2O2KnfZsv5KECe0fND0/Uc0WFQU
BmgjeJiaSwso5Hy1/S+dE6U3yfTGF4CGNc180XYJnaIepJl1h0mHCzflrw952olhsVewTSHWRYeM
0gdo7sIJrywKSQRKcO0BV69UhgDm/NnAeP+YVaIM9SBpngRs6uvI5chl9LWLCS5SxU94WbbUIhFj
BoTyHRyI90wSc317vLqECcD7dqk/qnyKOcA956nRhQg3ET6L3sx9a6eb6qACWkN3luGHHCYpkLFs
q6UPpzXjOJ5sg3klklBqjAlVUYqYG3Etk53xn760L+tfy8GSwN8U+t9PERCOs+HXhIs/4pFek0ud
yxPoepkZf4ZBQ2qMs7xdRdnbTWA9z/X9hQKVjPA+JbSYaCARwjejfCDAvo1ghjkeZDqaiH9qGthB
drb3rHlu19zDST9+4vgk6gyz/pj9Wm/YHX0acR8Li4hETW0d0hDYgbF/ePUVUvb4Cog4dXHabZR4
C8IHxrhy6IdqZ4vWDwWzcDjUE3WrnyMLADhKPzW9fj86fm/+BJdUyDN5gHao4OjxtKJDkWn3bZlB
Cv9vkKR0dJOUuFvhSlAYhvBp0lDCugaeRgzC6jjAwT/Q56ZPqiShJJJG8R+QNALdWzmy+91KMT4M
kGojaXoBs9vWyIftmcUoPkBkdH+b5tXCy/4+zpCdShrDIZC8PEwvn9EhzWuqL+fFsxFcusPWtKoW
8Zy5CZBqOskptaTJtl7Z+Sftug/H+6i3a9j962onsXroUTEnL/5eo7VQKSu8+fC2FVwYw34k3+ZW
VrMwJy6toK793F36qp0G1i065N6KJ7Iz00UJfm055qmBEXubDaP/V3Nq9sV528sugaPfbBUUX567
xZr/zIq2E3h8gSMTt9FbrjFEt6uf5W2OTiUpWoqqszB1m9rJZ6ehmBtCB2SYRgycC3TogSFCNaaA
HqKVsupbLAnF6JMvE06Eade1Za9y/Maihm1LP2a+TPQamckuyYm5ZAqNl/Aipd7CvC8Rhrj0CAzn
xuEgWaP+mzofV+edcT16bW/ow0LZ1cONaM6aa6xLeQmx+3xYk+JUDDgNor2kiMqqy4QG8Sa9g4GD
GpdGpbFSuNT4YVOUGf648yEUXv5whm4xpETfu6GAx+ndVEVCd4dxPp6bAiux7ntGChsBOUMWJ+E1
sl0o6/BWJ1kHoz8B6Jxiu5IdX+MJREKj+J4Du839WpJnUNBudBd7S15invW6oWtEFe4XL3CmtCrQ
n5Zqj05F2h5144AXZCy3+mO8TSjhcFc5IhGeTR8x3+0Wt3qpPao/duOvbAUxRScv1WWTk2Y/iapx
v9ZDLCofGRy2hBF8QQ8vCDHHIVDFVBwvRzDnciArHr0dZvMbslZnMw17quhtzlhZiOQkoW1myarJ
mqB7orT+FRDW3MfyB2FByCnZUnm3fTn3J5nluJRfGXdMyUuCRCyO5G1KXZj+UXOMsFKLx5LgumUO
GF+q0hdECRpMRCRRb8I9c1YjuDntaTeTWjw/MUmUFPJa6sjCsK4J/GNa4yx209LAPu9Lfy7Rh4x4
3LVVtp7RIMl5idTZBfp6b85//H1G+zAbTZnneXIsfvp5JCL9WSAtewQ/Hif6wJ4XA5F504ugKVYN
mcVbNa8kJE66W1MllpGoUOdJ5G/b2r+L0ycGaOWgKgu0B4eqrCIsdJZW5p9QvfUc16T1U4i7YVcl
hKuTiEdfuLP2K40nNSoKAektC4kmtxDf30ALrPR4OPT/vi4VYIENE7dTTy87O0CKErDG/rUx2Fba
5G9eqbVyw6l350AVyGPKAPFt7I/sdtYbIuafsy7rupccjUzM7SzrctLd+vMoNkS04njp/3CR5jbL
k00m212pUpZc1zVVXcmI43SU+rUp/8369ggnokCs4ukr0w3o/f2kdUpSZaOZk3jSJCInq0XQA6d7
oum8dGm4VpYF6guEdvWfjelu+uXuoHZmAY040NS40CmFsS0FalTeetMNOAGqRjN3OFbIqI8axaNK
1nlTTmk7L5MIF1bOHhJJelOFjp6G3wdOYT35JtGXWGL//RfxmgzPZ612ClD3HYLn3t1ifbkxc+Vz
0OPxqL3pfWhU6Fka21yN9hGrO00LWA7LtbXDTu4CSdeYAJqwsDNIdv4csJHcOAWFH2w/ePR+anaM
wlEj3bQ8Ix+JQbLQbM/R88ozEXbqeABgxe+DYB0z6VgrQQ/japAxsBzw2eEWu4NSx+Ik86awPldY
1fE7bFRTcIoZYORb2yhDEHt4Pw1VqOi3LkHPTKgDcTvczyjjT+YJMqHuANXqFsHbLYjUoT8J6+aL
oerR3IxTVp1/0LoAhf+4SRCqxxKDPh4vNDMSDDMOC7duFxuBOD9VUm3rH4HilvwD6WenLeHiX4Jl
l1GSmwI7WT8Ev3GuU87w0sTuSRVJqJfI3SM82XfYN3kH/YuggDseARlttMSj4T5VmXquMYDQ9C/J
0coyZzQg23yRDj+g6EACq2N9g6u8ojhFi+oaC8KFpXxEDzXhpNsa9Swo28XOyUXW/s5fqk7p3U4R
vDceWV1ReYPMv/r5qakc1SVndrkKNSI+rzFKt2QUSNuUiHtf5rQn7nifSG+QXryo4rIxLKJA9hCD
XTkPMpSObfwV4lvmBdUcPqEP96F4McI38KHTL2IjtxQAWOmbt6olao+hNFT+4nEgiPEF7ZiwhBgL
MgwukGSyNLrI8nIlwF3vU8HbV+GQgL81DBpjdgnmD+bhwsM509Fze1CwfsDJvX2cmuw9qnoUfILG
csDhLafsA3GsgXUC4ldJpV8IykHCeKc14aqd9WH7mNkRBOr8+lJAY+Uoyfy4UUv5+nyOKgekJ9M9
kCek1VYVjHGpgjJbvq3tw3psGFVAHsExdci5D6OUW+/Q/ai8z5PGy2LnpDExil17YChPZ6AyDFg6
vrf2y3OrNtqybw/mKhEjU3Xok8ZSCj7mqwW6bmotwMPTNrDaaxFD/DrzpYkIw6FD4nKXvTIVVEZI
E/OuDSrz/kSSEj2yLKz0LTXdDVq4aAazyP9z/F16EGO2pmjOy4Xqtm/GRLEKayo+7GwltscJRRWn
/VxdXRsrWu4GvegJ6gIu4Zyb3mab8GaULiMrURJZLFAJrf9XVzeP15GJnP9zZKs7o8cEtTeE1qdX
90puwFS2haZZbZDmavJyvpPDfIRMy3kxnJIWXF80Ik8xr5B+oJqBsGuiLJ0Nvvrm0fyQLT21ZmgM
DSfLBqnt3BTC9vJmDMUtsvMsJVl7AceZN/T0W6qF/0rWu312gGftItxObUSCRlezoypFzeDB4zgR
v6q3rEXHZyTgd7r89QXKSs3/2N1v+W99wE8LuHlNoAul+HgHwKqAU1jWxctO10ilPo3l5tW3fw+y
7IYIY+EWIuqzrQdgWxq0f1foYcALnI2jJXj05wMOLsTeECvDz4ix6BarYMwE3qDAom6Zh930NL/O
QU7n5LcvAHY137ipW0NcVZZDiWm1y8EJ6uLtuBWWoX+MuHpOP8HWcPACCLbF+Raj9IqiaPVaiOVJ
10GENgRdICIuP447tS44xyi3RvqcWyeIMtzXcEStfQPg0KqWdFEND8MHDgrjrozoG2NOG1zv1Mc+
iuUyKvLf6XRWb2/Pr/krJsK6a5DGVaVqGSU7X7dn1riQ6uYb1EwDHHACvJmno17OG2yo07TOu9Ow
HQZlQ8bqgC22AXr7zD+/EnGh1iFJDAcKZjDvLTjLh44KnPaLWY7jb1NsDXCgNeZeDQ+RORqh/E+Q
wZgOj2SMkEXW01bYo5FM3w+Kj6094+WuwY+iAUWvsPAS8aekZ02kTxbyzoIyyePH284aAHqo1xaF
i2ahy/F3GgSmYRwdn91b2Lh/fh4YDTrjnxy1mK3CmSRG1Wxa7S5MoHO5M06jpOJXZGeqS/G5q3Px
h7rm/I8TWGTyfsrp5qkWfrkSa2BG83GqGSBtsfffhNCvEW8p32XVnHbaX9hR3ufKIjfeyIVBOomv
485tco//87GNNbrwWiaTBJMfdeRcmbq98kWIBRUImSKMnt2OdBS4PpFCTWndg/ntniS/cDU53Gce
+yFc5qSutEp8sOgRB//whxfbXN8W5uNgyBJy5GZP8MgbR7dk2LX1BBIG9Soq89hP/GP9nu0lM4b2
URhT9dLMopfrY+8/q8wt7aqpXV1Ey4fr8BLvo8f2ziM7DmXUApfhPdMx+Us7wnO2R9CdGuPBheUz
Kh4rxaZlBNmbanNhVXx253boMUhD4RAwfWJ7NLMeiQPlmH6AlljaP+iJa4SqVOErJCujZRLdJCG/
ebAY45lglXSDlM1xACuA+FN//Raz4L1RUM1+B3c3Px9cY7aJFoheYOJz/FDgB1QgjfkJDlZpqzWU
MT1ly7ZXhziErLDxaCCWquiXYSI/panZ/poJnGHEcNqL5RRWmWLUvJjUoaBVIzpvrGgsLo4hyYrL
wAPbahqm6g0AEOEN91jp0N2ynn1AIbVdBpTwugA/akXOEYnatbE9TV6zklVUWqCdiqob+JVZS/k3
XBu8t9SuBheCVWrij3oUK/J1X9Ti5fcP5YBTFwng6XRVWovlEXT4RzY2W6wvxbvOelvLysfKMhxz
AlECuvueXFDIp6GhVK1zrDBIGJcoP3ezsmgl+9W6mbq75jJrmsZG85ngegJ9RxEeQghxaybxVq1Z
No6elnpJUWVVbNfONmBZqj1eCS7uLO+MTva/F6A/mnDXbtFgDXt+6bGcorW9UrbXhRT77XaXK2Uk
45WxjFeT67tiJyoEha+sk2ne/axOnU7fRnkQlfh8shPA/ZL/sNkO9/rqvfPx21VRdNrJWhUyVbMu
9J3ceg5QsUnUdFuBxqk5ntJuTN+16VyUyUee0O12yLn0kd4hC1jqr2UTwg8WeG1oLnRx7/KnwTpi
iw57othUwZGUEe33yIRy64bxUFa5SAU5V22QNVWLVBXeJ7xtpeThkn4Eht1hc0J3m4AiQ085CTKf
aW/c2wV8TXFmwhwQxCKLrUCKR9zDZMa5wCQJVCPxoUU+bjh8t6eqohdOMXusHrQzIogdQPtSc4mx
hCkugAaKDyCeB/m0voNgoN2C2FxS99tVxtdcCl3uELhZcczvrF+/cFOZ5rt/+yQL6Y1tt9h4KcCz
Ftd4rP5Xpvg8C/qe+/FZiJ6SKRCVR7nU0MxmC3VsVF5TMmnljERCL++0VkciCdT09pyhogQ0zzXH
3H1t04dQrqG5lMYAfieefsGBS2ttJ4vVCloL+eADdCd9wJ8aqmv2QVK+WzJVSnfDGGpSJcEkCbeH
2wHsjq4FIpnsz/tNyNXFsHrB9SnFF1TWN93l40ux3CzAWg9xhYvFgOE90oEKNf6N4miaRgDApoKl
6oW2Wf/5gGYrioKUjCM/bev0JMupA1dlJbUUhSKPWJhuGl8hDlp9CzE7ZEutgGTlUi0XLQ5kaecS
rF5yikarLiSrKYC7rWjmtyPkv6IcO1FNp34BDLOQlcDt+yYK6T9+ZXaC0SFblra8xwgZft9rqenv
52uqXhjvqucbWPjNYivMb+ZLItx57+KZRIeRC8ZlydPO7S7dXH1CRp7kRc7QldCVkJ6OeJPjFEXu
KaGqUkdchh7kUCliYzlviWHkPy/jYa5LnilmZVF49YAPcFxuZxFs5O+PdKv2j5ymk8K55D8jHeh4
MKSkCBHXwkzYPDnIRVa3SqYAqG11YfEL7vApH0z91VUj2LC8eQ1wRktfw4Dxn4nIpd8ErRJeQYxD
ekDNTcWCxLLxkDvUIbUkQ1vVFWZ+2qdjV0kV96cRxwPy/4NpZNSDEYuSlvPyr2edVgo38isK+Dwp
hvqaKLY20jubAdevha5L3SvDGLzBumd99e7/tNzzjF+Tpjk22p72pKcDovfUwNJwHxlDUNeCPYeV
pCFUALDZ+3lRC1dyWA/vFh50ivYt9TsutPl7ZEbR6t4cjO7jilDywC/DS1/dKt3/njYR4UpY/l5Z
amdy9ZUFkdn40BxPHGd56waRROpMdf0wmhyCE6ZmJOB0JavPlIXLlHTIfk9ECIZ5H3cl+4HzfZyq
v4MDCRoJSqMwdsBLhyAsKYBmgi4cmsHrFns4LtJnY7TIMBqXd2rX/e+sxgac7e3wqZhmdyu0xW6E
PijLxJ8EGoLWDfb5pu8clYgxjeJ8gl5tnQnyFEnNPpzt4V/Wrty+1ESwpxKMzU0w3mPQjGvp7d/D
GpD5X3epnyBXR/4iupDIXyywuFmtrJ7s4GSbs74MK1eJHeykkUSsXtTLJaET0TTPIxKXc0EHt+mu
tlWYbaMUdKXfzAsd1/AeY907Xzhn1BEG82/Y5g16SeiFUbZQRpGnRoJM/joX8T5VMXh4KX/LDs38
1Y2LdzMIGF6Hnc5v8fTWOuLBWW5GrcFUvz5s28ItlC90cJaIBFIFEHtT9QMNgASlFQ5ffoWUnZyN
67rzjD9ZX6gxaPOiSLD8Ko+hoHEahyBJNW3vaAvFk/xvxAemIqE/wyp7pR5bVByh7roTOcVqfFnO
QJZD/0f+mZQYm9N4ImdmWZbyzq1Jphe3h+ZOnc5DpTBO7KVIr0Z4KEMpYCFTlmnT6kTLpqmss45b
aN/ekUucbz8QXGjUaCaUheOsOVdgPI9KoZk6ZXbfyrLtub21xcGSE4jlB0FTvuoIwylur9vvLFCV
OJRNTHO+nNjQNMzfvkp3MeRVXZb+tgqIrp7S0YRnSzm3hfESYspPueFgzi/MSJeUJ24GzpKQffu0
h9V4Va9T1XT0KE/5cElEC+TGpsH3ln2R0f8Sok+mXmwcLaSAhF4EYi9wnWwYxam2G438ZewOVej7
P8nIow2xu8ywDMjTwV65Z8D8P9Ui6HX/V2W4QsaagDMVVGMxmgIePSFn2I0QtBIzIUnl52zJNx3J
DIqgxBPthJmOB+2AqpAEUuzPIg+XqYAHS6Ba3PJdCYyO+QImezSZ49E2+wDVK2QU0s6W1EhvC5rt
6Tkw5WFCot60/CF4M70hLAnqE1zaYsWQVneIRpHd1kwX+n/CEddSi51nx6UVeTML5DoOGtqGvXkO
0b6Ic6pN+6yxQ7ybsC7ZOaClJQOugvYTH4RcElAshAzGzv3NPjAuvtOFAFeKleA052iIMK0NC4ms
AFgIJrkDh8g2vs9ZP9HBgZY2ER810ZzuTtA2Wvz+Ys8U3KFKzd3xSAuOQ9EZnJtW4l9FmQEy6UZO
9hUugMSKgPhMRCZkR8T4kaVvo9Ul251bnGIxSH2F8XA78mBpsanP3fliRQys737dyuPNGP1mmHq6
PIU5ppruL0NS8lwmpJQYLkyEBRt+1gDYmpZ9t776LJQJyb7vnQSyUOvxAicxM15wa1AiVbK77n1D
W4cnD+S3tJAKpFVpja7nIwwgRaz8FxRELFGuV6Tuyw/2fVv0kMc0dALXwN2eXGyq+r+s9WGxdfDB
8pFSMkbyF+CIPtXGGN8zpI8xTEHjF5IIq1fKSH/qpMUI8BdMzAQ4k5gj4rskYLk1op7npyQf75pY
W0gmgzU0w8GoBucKg1wxPRbmu2XPDfMsCdWS/oQaBpSEfiMJqxsNEZaQbN1YMBGYxIXZy2HlnBLV
rbUCuKUTaqWu1akf49SGNsiF1RHFFAOQAmVBg/218TsySsIM6KjqidhKo8CdSBy663lXWKAIUwOa
XgxNXm2Q9Lcn8krAGK3hIN0kzUHwtSs+6BaVR7E+BMD7R5cqCvT+YGKoWrcFe45XSAQlZ+M/OybU
xdG5nocdZzD8Jgv0FnJn/CDPrqxDq9a3z4f87cMKkEX9rYgkwGCByt3OXsGGLj/d3D6bLGV/xcb4
EE0rIYLOQWOvYtsp9OJv5aVMu+eADvroJTis0DsqC9JtsoP08ieUz9Lvj57fawJ4Z48dQOx/uCyl
3j4Pm9tuoImJN+O2k+EpIZRqDQ/m7JCFp+nSiEETgHHxgQDlYoMMlwszykkupvxT5rXAzRj61rw1
1Py2nxUUBw+MSEwEqI9xPTRs/H5CuQx+bratlELotVD5CGnxXk1V9k/ATPG2cn6uwWxiWJP+fM49
MnSjH5EPejb2Or/scKzpLD3RK8Lql7mwMJLsJ4dtnDn4SJt0IkXARtwgrQxiB8KZjnF0wNMpsQxk
f/tbqspL26pHd2Fj/QqB8HmxarEBnLpjN/Ppwp6jzrtXygXc1xIXpMILwuOfWl2h6uyfG21jzkOC
v51KlzD991nKgYqMXV0HDZfL2YfTGxCvN7Dv2sBS/mTbquHS3Igj5JsZebnKhcxg00XSqhat/Hff
QxpAF0xXPQeLlubln/T824p2KASD2d6KAfo7yIPl3B9TEK96V50XyaMDcSiSEX7VussD4o0pRlBW
PPWBbSL4jGzoYUPsOBKreIohOUcXh9ZNlsUhmUnszqVtSNGtS7mwgCGM7FrqSxJ9SNVjbi/ij4LD
/b7Z7D4a4wAum6UYYVM+yh+2QOIPSdTAInV9FcOZA9qNV/sOlT1pBg2USvEOeb0oK4B0wQrry21L
gEa9HSe5UFDZDAqgpNuMmELmyuh7xxD0MWV2xlKm3Ot71qLCrCE8Q1CM4XwutDpiTbqqTBOAam6v
iT9irNTdAw0E0QTjIYNoY90NkGnw2wzU6CnJDLDm0qSkTHi0RH7ONxV+4MdYBa8uHKTtbHazMKUm
vAfTrdFQ54X4F6SKHi1JuJFcBJn+8TzPKoCNgMVqRQDaH2QLxsS/E61Yc7MaZST82/DjxYAP1tHs
21a6WOO+UpRc48b/mkcRABM/GyA1uxFEFBFas2hvE9q2ZvV+Ude9L4g1ZwVFuAFr0ASPX/SocXAa
oNZJJguhiuYsAVFJDI4T6UqbydgmaKfYTaywcasYSdr6P+9kX7rHcCKBiCZiZ6p9s0aeYrSzm6l2
Xv9rGwgrZnWOzD2IHzi6trwkUIcdFmfieNr2YT6tdRueZP41yzmWUGtRQdc6jfh/SqGchPjqIz2w
qOMulP5vAKkfJ1Y8gonmiYoz+of4MAq/mt4hFgeDYNDjc1p2WQJ7BWUUZOUSNLB4jwoI5RZBM92R
Jq8Fp/iwBJ94Yuxyho8xqe4+eVX2R+rppWZ6pnvJ33yPagwhqvEczZVUJo78A36lC2CXu4f/38po
3AE265aCIxsaNHezzDtVQrJk5FSqut+CWpsCA+4YNkYmc8HugvVAcIlHl/4ccCg7AqS7HvVnjxwz
OZPWeOqoN9Nwk6JeK92l7OEXwWkhEtLE5/xR1c16VRIdouMJ26TRbRDXQbSOq5QtxqtsaBIz2ZZK
sUP+0ohJ2zWVGpMvCHhFZeAh5BhEfZj5lMjx3/bwjTRMf70I42qyzRyJ2hWAvwjt8DbD47/oV8Op
4aMgEUQLyYEtOjYej60pgyomVQDDO66EYbhhjiMMWqlikB9QubWiRdl8YhPrshTtLF3tnEgRROpA
6hBiezzpHgC24ChTWc+00QmkruKe316WLoAz4EDIvyIU1LrHJee9UJVTLTqjxvoUciZvfA/gJKd/
CSACgp44AOMs04jTxXhKHRECFmGqfOu5KtZlYBiOyt0Tynpp5dKKUj1lBkuQeFeGMZiVrQ3t5ePn
tyCgaN/YsEHaDo6QY8sAdnloHcsF+d8l2d2It9QNgxCy9LqCMTRyQaOJzQX03SAiCcqUnEmipRth
10Cay0qBuzyE9Bs9XuIreGYCr0IZCqJwVqr1IuaIFucKyD8FJsiT9A6AtnVFlPWy0iNF05a/0FqY
ObmetcMqMj8NA87GNjGls7fWoENXi9VOj64B9iJqit6TaiRHgud+4YebdKEd3dBXYD85RMMeAEHy
KhdcfO5x2doJd4TKlExC1Y039rKHBJgfhLWTTZA4efztL0UBzwZ6Z4Yr593KYWDBdHBm+OflFPIu
FTqel5SQzNE8XfbF2+VPCfF2DVEnwgkAVWP0HzsavFFiTt7w0gHwcKjVMQY02+lck1ZIyO5GtkOW
9pv3Q3VjIhGocmngxJpIdNck0X4r60f2TPKFUXddY/kp1YMvPPGbFpdJdJ1CxgvCXWHPD/3H9iix
h300yJdi2sxUCBJ7gzIuuPE0S4VQsog+X5l0tBWBpjRg1C3EgZlD4NtBa3VgkqXM+JIGGVsKkOZr
vkk3O7DGKItreG44hI6aRFpWOYA4yNSuL2ls/JGT1XlF2SSz/90P857rEUhy7jnHE/fu1O3D2R5X
RDXyIBTm1MQH4/uXkZcb9Qw/ORYmvqUwWhN3jhGt2ZXJNTBAE4TOlmj5ad7VjPKeVo4zt0adrilr
OH/x03HHCH2G2U0F0fbMPmMxNSdrj2mwy8DgwJjDafcCf3qXXFQZOIvmFWf7CshgV/UDThv4ZrIl
Q/rOgrIvCYhnoHAg3c4hQg4lslF98JkWqsziIwSda+OYvfaztaIp59kKaqyGhhj5d80+m+WHTr9u
55NsioAWt6Upf9JLxFg2uISYGPxdZEwJEOix3cEJakAzB7j8VPcnwCZRl+jYOzcjvcXyVusLyIz1
ncY/FwQL66qEHGv65iVa4oH+sarN+GrZwOZXXVPbjxcaNgloiCe+0gO/uqPRzBPZzxvRz8qh116t
pLNkolHCGhp73i5uNerwBSjlfzPqklh8t3NAkXhMQKltUZ0jz1ADABtMeiPs1Mhamb3ZrM8vpIeh
A+oGn9OuXCtrbiBBKnLiBGr6wsnEhVLFRZ0tdtC9lYXhdrLR6iuCl0Ogyl4tARQcH6FOAQZdhbqy
lUzssYz/HwLxtcfiK/brxOn6ZnvzWg/n6v+e1FGm2xuUCKx61ERGNiB/XP/boVykquXs3T/GNGPV
USskXaMyFpWKRNagltfbIbuqZjf5192gIm2UNQfidAjIQhNHNPI56VIqVKIQ5NuEfx7TQPy301Lb
V4z0n5kK11B/GBaKoeIsAX9z9HHsXlYkNIlD00d1fectepGFF6Wk4VpjbL5nsXJv2SCTwPxjfRTQ
4TJpEgZMsqXmblRN8fxr8DG3y3NwbTrq5B/yDkJR6XJq0T3KDBzk6Yd4ocFRG2ynFa6h0TZQpRWW
OSdOvjbQ48nbNzZe1UXmA8nWk2u8xkOknHKlxEJ8IBK0DIGPvuidGgv1/+Wabq8xcGY2IqcVLST6
+bl7uvxIj/B2ibJI+nhn6cgeSe0tupVZakfToW7FuNLC5IAKOihbiBj4R5/4vdwF76qG03STV3GU
Hr4PpuRQPogne6BK9lh7HkVsd1szFGujFKZbV/IRlKwbE23NaI3YnAmw42jSbc+Hpg7er8lmSpP7
KF1ow3ZChoj5fRIb3re2uu8fSvFHq9I7sHmzWjbIWx81VXuwrPRbUSnGc6NqzfM297etXs4kRME4
c6fbGosJUDDhu2yYSLAeJ7790hTL3M25TOFqo561Vs46wEUHtmzPX0kBlK3x5QDHUEZkZBIRCPhH
N3F24+2Ki/XqZ8UsgP4+exPGAfoxlFt9ztRyTyPkB0Q1PnNmf5bvAf0Kt0Z4o2y7U4/XxkiiCKif
+PqEF8Rr3sh8eXC/46B2pZ9Ux0Av4fdJQIwR1THJzTdaUj3VLjsL0XIgFibkmrOsPTbhw1MgbreC
0DXWtdMnBt7JyawQSaIV51j57bV2dS5SeLjVN/ThYfp+vAlez33z9eUEaNmUum0uPNTBz3yZHUvQ
zBr+tzQe/ihzHmqoBxohGbxja9V8CXhj0qKWuHGqQnywSINWo1tTywYi3fcCX+KdMWzUTy1Tg+8q
KLpNFrNqkpWA7QpzBwcmHsOFSgOhejwJyRUR/vQSbd5Pm8suu1ZSqWh2K2DQ5P6PIHcai4pXOiQH
dFKLDJLRnCnBQSHNfYdWyvtTRMJ19owpWpaNWTwr2cjAvz//hq5XiC8M0Egytqdky0sGPNp4VLu7
tuePAR1Hi130x2o7KNGRK9Qrm4OSEO4o8/tERo1uQk9dN+y26uDk9aNz1N9vK5UtxVhsI029W7yd
vfSudXewCeQUMlf1Y0172GBFQ/w0ymOeAikTv1xyMNDyNTU5wy+Nawe/RnrFYtnSBKGS08G4IzQ/
1SBTUYlPuAANS+/5FCGrnOEAlSM0k1zPuAe5xzZwrTKn4/upgyAAb4FcVf0ifGmksl/BdEIIdyio
cRDaFNwouhGkmQLsQBMYr6OmTQGOukoVkx47ULkihh204YVCzLvB0siQ38jTAmKbX7CRBduFa9gB
pjSDFYrURvKhGGAU+uRRW7y3E5+qDWNOtRZYClNsfdczzZrC238J4xJwYlx6d/Vg2FZEqeJyc3uN
CLOQNy34odt4cptSmmD11MTtisocg3ehplPK/8YcuUiO8cFPTLFp24BNU3NgW1TR8qebHQLBNyTd
iGQQM6mOc3CX8Ych12bUNk+V6beVdkydKCn12Rln8KGGgn3XGCUI8mC2oUmu1dX8g4wXfZGMjp7h
jyTlbZwAY6Czuc8Jr+k5GBCoEvhrvS3pfqJgD/BIDrprSo6J4ryIYwPtRVL7IMcQm0BKXj5miLCg
m4ZFrIWEm+UmdMWvf7m89K/6Qwcffnss24YvK7iSVL0vJ9u9xe2uFJ7EdB0fBkwdxiK8qR6RHSBU
oo2fI0t/Xj73fc4kGY1WgLj+cZsZd6UkhU7NNjJhSQHAevZIzuTRT7LB1pqgxMZCc3gXJmSBAfnU
eB4m6YKxbN3X2rncZVds0l44qDBxQhrsHp7NhNW9VVth+FIuw11wlVoGS6zMGs9TFLXrufk+BjHJ
zcIpmfjj4NEJQrXQUN2upMRzFP4J6UXqjp0w+3gxvf/FKLq3gM922NRcbRv0SWKamvuI6pZ786r+
5Vtht1IV4r9X9XUFjsZXSuJk83uXbq7zlUmcKI9GaR6xadktomVQkKd1L2CEkJyukUaoG3GEANpx
23jNioYBeKGs9v9naaUR1yaBZFTltVZ6UsNm7Jz1cO2Wr3P7LL2oThxE0+Dbn1KqMlNkITW2U7Dw
1I3EYSXDURfITOIJx4IY07tq+NxRbHwvKpg2N0+JjdZAD+rVbz3j18D2sVZzbimjLYKtzqMQ/QHo
M27b0terdqP7kWhG6/JlQfVp9tVhTtX1F5cQPG+9PzxPKAEKChP9iTNrrFpyBuMpY6dl+P2Yo3XA
w5OQhyYvwQYv2RWSzE53m4qI98t/C6Z+NSClh5DZKeHMReZN9GueNoyurG5sAY6LHIVTBOT2iFHx
y91qI+sTHle8bdyGU7gj2ymZfLiXSLle1iEr56rD/0sfJx2HvMeIU8IZDbyMUVUtmvkrYxdoLviB
klgVHuKOEpMn/zuBg24ZKLEhL4KJiBtwmycOK0JCw+6sSFDEFpYT1yUo+DsjpOdid5ovgP1hRL3Z
UPY/yp1yq9S+Yz5jsA5PRd8mjaIF1ruOaRzf8/xRKtiRYen1lLJiYcbWbYfmX9zptfdRlCFMGYhS
UdUEENrlInjsHT1icuuW7cF161gyZghGlIWPaMAUpmCpYSJYk5FOrAV+y84+x3mOKsB2cjn/I4Fu
gsj1d7lGmN2NitSVJOhGa+cwqHKViy6ja4Nk0RCyKrrIJSJUplc4WOt3+TrKHULi4b013pDO1T/x
6ssMK3ErccoY73Agxf+1QDGf0Yoz7aFpYFIAXvMPjpxQSCEyN/QLKSumJuW1bK49QcKelJxmeJkQ
sNPIKZG2vI5cbF0LVePwoKkIBimGQT0NcKPcjOVigLnZfWeQsSYewCZQ6GR5Hns6v7vhQZcVCZUE
oqXKgiDwOa1DhYI0En4kGy+x0M5ac7ahuB3GEWYkfT+yIxJ0yekodlstjES5urqVZtGcFZG0H952
XnBluAhX0Z/f/xZtCVGk0B1tkjQC2cXyLFdNFDmS27xZRwXiFjnPgwXZkUZnV9QjeRV5vQMSIv+7
+lVEbc3DTpOlpPzVqlNfgUPe1N+dttnMojVRPGxGBn8EFovlHQURQ2XkWDbR9m0Jv/ehlupLAS6v
be2RZ9rZzi9MQgNkkExNbSyyvsilHRPTzyd+4non91UBrPrqAV5ib5jMHfSj1UtlACRBtnIxrqXo
Afct8Xcrc2WBRC4RKynYFCdtcycopMskxinFkZpXVd+K4mr6PhTe21xNarl3ZusjccG/1uGStVoU
tM6D2Y9WFWLhnnUrW//v/m3SOCMnYpFC6SAWz2i1dftZQR4tqyU1++JBZiZP5RS6NAnmnCKrPRWW
NcZs5HzW3GpMREj4Tu8VrJEI1rI7SGAB88Yy6e1oVy8WuUeUTAOwxtry5F3+sFLCnHHhgZjBGV/2
CYNW/W2QXzlz8mzacH735yng+RQqB+Pt64ZRC+ipqEnh61HXc4iWJjf8QDrfc1abOqE8C9hnFcr9
vHyV9A01N0jnVd2ZuOaaSynKZcLynkhPUr2Dki4p7kbBqR4n2hRNx2YU+t4yXdIxgTwLWdjDz9Uq
5RK+k1XFaieuETByx+QJC8GF4kBj6ruTYKiiglofJVQZeoV15SNk/dVDUp1xu6+1+XQq6CDACrb6
UXw6/8FeWse+A/jr7aO9d9gDgjxLN4C6l2vaKnn/tbRWt8y9pCX/qe82Y8vPsN/2YhuY8TnTWi+Z
yYeYGV94g+YY4Ud26nCjvAHaby4YvJqebkzcKJkRukGog9Cj9iTaAzAdtFPBHgO2hXMfP9cSOygk
fkr4EbTvFwc1OnVO5QwlWu2fJQpQOl8Pdme+1wXy/PnIMorl3NaOcc/dWDl4kn31pKnsnFLrVsgC
t2Wy4m8uX11V2DeiNDLtQKCjidlDoNnQBJgClR1/Sz1qCKym+eS1XyA+HpY0fhGJj0bz+vqSbf7C
InFetR2fbZKWO93mi5b6olJVzGvQ+EZnQGw3UdDILm79ULzVvnTHNXwdBiUEWiy+OymCy5jFyy6W
3ikS8771gmCktGYGpjSqTpYH81IZTkCp6DV0EMnUvTkvCkS0iID9Hg/heySH6ZHXMGUpv8UOkSzb
QGSzbfKaCR0VIuK3h41xozjZ6obRazjb77q9BBtKWl4wpzH8LPLMguo69xIk1M64xj42L1vqu0qV
nXDH8xEnNvKF27WnxdsSo/e/rvDQ5Z3ZTpJKV8VErbnJUfdDbCwBd3V3ic4Z52P9rAcR6LRrXX+k
sz2pkt2rV+e6iDRQ6fAOXlldwXF1v1sVoSey7i2CY/782N4sfVmgROcVG2LinAr5sNdLvDeDsyEZ
SyaEhvLF4jDNEw4zYH+nK7dUfWtt9JmFCJ4rWQQv81Uhnqb/zSJlUvm6sKBv4go106Xmb+3PlpOD
5Um3wGFV1/YuxuyX0fzvgNhFYdYBuBqO2JEJRP2y+DlkLW7vf61pqxaj/FovCFHUPa9Og3LNvqZH
1qk7CJr0Z9TTGFzFuRu4hKOQMjUjw1IkTlMXzVRS1XbTUz1aIGRG9B87MHVlNwdpuq49yxYnCw5T
lgZJUNi8mljrwfuPV+7rrseHt+2mx6KnYZfm/U33c1D+fCXkIDRgV/K/XphO8bncERJdjVqOjrnb
B8cCyy+onKDl/h5AnvowTk95vPBa0HLC2yAL+P/AGwFvEPGeF+LCgTbG7HGCt4KZ0g+MdrwkL7g1
BtBNhKR9E3wF5DTCoghrRRKBaJIe+yfIIsiLOtefEe6GsVqu8qkXvVyz3NBjlAZ16xvmSWHqrquw
ng2Vs5Bx+IIGnUvC20SWMlLWEULs9R1ycm+DyCOAJu7qco1ssOPZUAhIkMW4kXeehkXLZ+nL8NC6
s1Fk0ewH9aPGTBIh0vlKDmZeBXDCS4Qa6zVyPnsQQVNQ74Pg4M7viFwZY17+HcA0RJbDILRYvME0
oN/dMwif0vhQ19VpYI1KMVFsJc+/OE53cYi53uzWSZAIArkrxrLmNVfbAFWdAWekiO/GzQnhXlWU
HlIwKhMJBM0H4jH9sU9iTsBgWiL6JRUY9AMOxfEeXotcPf2nkcrgeutqJJHSLvXRXvfT3xWT224X
wkbX6XmgXDh1BETtCoLpykKIm/lYwGkd3FDxpLnsXmxoOEMWqnWdS84BNs77DaRJC5I5vVvLsVvJ
RJHcUUnR3Tu/vqpg9KngCCtIN8Q1gppULIhplLrSmONtC4bYTphxyvcqz8clq/PD5mmR2weIZCqN
iZGK17F7OWUExyOV8sol3VAyMny5NKRGBqfMKNVF40A8SqogTwY/ivdoFcGU7BCEt6eSMG8RwsE/
scLI4q8Bb1dRI0TbQNtTHJpnw85+Gz1i6D3xEEP1kX1HgzKKiFKT1R35SOEARSLNQFrID2o/TNDe
YXbc+s+7n18Q3mHY+uUTDcY36Gua5i5nP73IETf49NRPtDi/TPZ4CVe82LWY2WP2jqawO1N9BKKm
Q0vKLMozvPNG+bgCbhiev4fyHOeOeFlt+4Xkg5uERM3j/mII6ef544cd+fL/XYKPOz8r6WnlY8Bg
zAbDzyjny6c9tfdnVBXVOdFoyowMRrkCKwZEhTSChJOcT7EJncOZGkgulJxnXeZpEHV2IZe3PmH1
0n3ayxmNA4XqYJSt1/E5+OSITqfzt2fzIYn3O9Q8IZljZIGGHtw9GSo/FRBktka9IkLzag2P/Yww
pbO/Zep3C5YFPYdPBb43Bc/bk3CMPk2QF84oAORoss5yGXW7kRH1VIDAvff//GfKXwec+vXm3FXl
xkcptGz15QwERE8927cHe02C12bELhlcmbDqPZZDvVZLFgdPxSzz6V1Z4/p8TL4utLfas2E8x62S
msXzbIk7Z3p7R5RC8yXP6Chics8VvT22clfDnZCpNDuOP8BV9EZMjlrLK2uiXcQPIKqcTuYtdSWL
GHXLIavrA9ClwktQd7XEDlp7+OJwPXN24nTUpNHfF4ZWA0jH6ymBs2Pyt2wgFRinvEsm0CPfYVGE
EZuuroZZqeDUuhiOZfG6onDdCg0sr9Upb6e86JbgyrlQUS2bZ7JyGW3ppZeaJacemdX2IUGMaYms
eboBUptZQlz9Dz3ef7iHbcGHiwVtmr+wJfAOFV8sIQgHEWoqHWAslbwcjGkBKY5Go23QNQ5utAfh
f9c5xoJtRvIG6FLGjNJ1t6aKJwtnD0WoXhawcJXJLrZfAAgPuwyPhDATWNAIJRFMIte1cg4MhTOl
JQTo9sni737Q7/rgyGTJi9yakv1/uq/5AZp4nE1k9yYPjQ3IQmG2iYC+bnHt9hUjltv8MJ8mOn9t
fCnvgNFl6WkAZmAjDEqg0UMQKFgkDbPD0e5DTPl4ilVTZrmF+ciNDh6YYgEpI7J0ay6FN7fta8Qv
oA1nN4yHw7a1Or/+Du6RrVO2D4sF7pdSImhZVUxKxpfEnmJvHe8OESEvr33MG3ooqBLiAwdkVJZg
T8jEIWijZdHWJsPD7k4alodGNl19KUoopaDGkA3BiOY4Hcne0kGNxRVlDZnlPUC8hM0RZDk9DuSX
11z6HphLxtC3SsZqMV6Ce9mvqQ80qb/J1FfcC81UWFbAXIwMoj4YILpLJJ4gmGr6M0NdKQaZC89y
1/dvA9LM+4L6oe1sGCPs3AYrdZYw0hPhFQYS6o6CzV7oMscac3sfeaE1Nng3frQ1GRPUuhsJrqDh
kF3OMGssu8Ktqvr23k7/Z7NGR/P4mXA8wQRzDH8EztE5a5n8r6zu5xTvdpiCKkO/mEaT2lN5njnK
RMDsw4IhyvWL3XMv+lZZ1lnIOiasAtknWxn3I15yRgeCpDkS4HSkkOYL88jZ9Tv1cxWmYLpvnFjj
CDSF6Vbk2VknlpQcFqfUnuwOcXVOhWOR/wIDSvjHylif56SZ1KfPseu22pH1QcAyeJEYbmkP9+qZ
GDyj8AgxQy4U8nxisxkvSE7xkQIFbNDCxxwwnmEedDeb3iYchibc2dBq5FRASUgxAEweKm+bPySu
CiUL5Yy2s9dbmK0VvAoN79f870N+bt5afKg03RhuZ1DjakX20MeGenj2JRwhg17l7PTYgBUtELgY
QOLPWQdqeJVGwe+NaXAhMXeFsCqgEp9cSzh3DCR7SR7Dwfl6bRJOk363HENQvx6gd6p2DXvkk0Q5
RNqhvZdspqOohvlcGnAgMJAq1RitMUZW8oC5ZN994v86YAOarFwdDAPn/NWdDF5vhg4dgTipoU1B
B3S1mX3wgx0lxYic9bGb/QwgKIbGONjF2tSnP9o3a1PPZTFbIFiJG3n7MneOkW+5HZyk6mVPEKV9
07Ev6A5De+z/WoJtIwaOHZFCfrODe+fAGQDDuF+uxaoRRt3VpUS9W60dniVf/Ya+0MDF+HPHfHEx
LKxb10bLn5dtEzTWeAKT1Bv8TR+8oTkglKhyUX46zmUlyDEgRZOJp/wWqom6Axlvuk0bwWbSpZAx
RfxuNMYjoIoInu/mIgzAD5YLkNkFjSEKU6cfNi7wEpr4HsFZiCNFZS2UcTyL+YC8FCmxefjJq94n
SjSqJqj1btm7jnkCvuyHQZpiTB1yLdY9aP9a6jBVitEpZNpNzRpbVKKOYCEZDPxwo6mFdgwAkRO+
yH/Li0GN+2nxhMboEJ42vrTFN8keesWW6AdhQ4/xdD/iANetZcvxlE0Em2EJWnzNzTlt3XI2AhV/
aylTv2fqlrGF3uHf0tJh+2Io43jSCI3uMz+h5jSsRuvXfJvOnvQ2+GFrInschGSJj0/z7g6uiuby
sdWkVyALFeZL5oa10n4m2v8g+fAWyAn3GfHO/+JFZPRDZoiYI2YQ9QIYKmOCzI+eDA0XREvx+QY1
ixfEDnVfIsEpgj1jeCiRFHEkbEQz7D5BN64kV78ZvOi43KHqtN/QCwgCpjgGvi13kS2rUi5W/3pp
egRyBBSFb6RBwFcdQEF5R3e2j6xZCUVL/nXKCrt5f3KDkIoNCka8m73chVF0jZJ6rf2NHBhzqiGA
p8+4NJgD6Yemu0BKkJdB5R+gnGCZn3o0zwVeRu2CIv2s/l9Hen2Ba1/sNy8+T5R0HjQtE3zX5nMM
ZIOcwRExCkp8Nail40H4ZauUQvffmw9m/1FKhkyrpU1RYoNYkW1ZiSTMk43vTILgX7wQdS4hXyyn
JwenLYAnRgXMfRY4MGckOR8SdoH8FhBO7IZt4B3M3NrfQxnuXcxoEcLVx8jSv6KzIBf/ykiY2YlY
OQ9Cq2zQ8aEIcEMXqpMkFSWbWNrJkPUu5hfMeQFyNLgZ2CMPOANVyKQW1cwxPMlYW04Eprd4c0bx
CDD7EsJ3Os3/lVXbZNQkXIMfwKhLbxSFa6sAM1LQ7pPZD2LRY3FzobJm+NcpPY5aPxttcRyxd7vZ
iL8ZyS+isnWoWhCpSe+K/YFkaxJsZE0HmCpJKuiNWkvwyOnoAl5Fn9O50+fZAQ4CHch1qeqMhapu
8L/u6HFAvoIN5e365gTD5EH7kj0ab8eY0fyEmwE/GxbjcdkhktsD8Ai9bmd8P5BzhLYBA+Cv4u1q
T8ffvDe5RxCKPF1Ek+6q8KaMUwSZwbbley0YEbjzRj+doN/I7AzMGoyfTPADAa8GeSLj9VYCjsfV
AABcK8qqX2a2BYHQI23VyVaoKLK+KQXygTmGgPUSRsmsvP5vnMzoulZzBa0ySXilrT9szBsWOQSS
YVo5HTcW6Ai7+TlpqObBoqs77plQFb7Oax6gl5PooL5hdET7mPV0Lavw5r9kVjA1CjdGdDm5Ixk4
OIjx2ib6yHKOQ2J7UBQmT0LHAytyra5rNrGBjic+OUQQbhTtZlMe4Tbvb2D1a64xz8sEzLvtY5Pr
YAvWHtuJwZpGdtqa00+4svNBY68VBz/Puy2d5eIHhXUdA5u28CqDTf6soTRCAAfFhBRXNs9/mRhW
WgOsLF4o48zi8jNgGlHFPImuUSu4lSdNH7n2WZmYLN2dJIqqT7AHl7opz7fbFQ8l7yCO1MQP3jB3
df3Hp8CDQfbsX0f7gTaukwJG6VEi4OmKiDVgCjt5CFudSugKL0g21qApFRz/mlk3ED7h2tYh20RH
IRzusTQUfYT5qtYb97Wb9e4Y4RoaC9u42aMpgxIzNPQI3TQYkC6gXnVtw9AwbUpTNOKoQOCK8cYl
cPLdYJ3FrY+5BhS2R1xwgH9CkqqI3t9Ndx1jbO+pIyoRZTqRO7n21NFRn93gs51X/VIxzGkIuyE1
pRmpEUZWFi3X09JApb6gXwvgAGgh9wQvTJlBHfCKUdYtT0RPL92sOaNDZjplBh5HoIGFwt7qCp+w
J9AXZ4NsEJloGIXSiP6cvYh2xT9PWIcyCDpbngWxbwILu4C3cw2PUul8IVHsH3PnyZ4RKLjjgHtY
ZWSb74JurRsyvQojT9QEMrJ+sqSLmqm2IbEkWLgLDCwBS51aTjdynT1BxadEOFYyS/DOCSEHJqRR
eZDyJQAqHkL+TfmFBsvtk5Ej/PzWZYsJXTKfRJ5l3DBIWLgBwclIXtB1D3rJoND71vWqbgVF0tv4
bfBQW0cw1PNwTwZ2EwGl9Q6p82qmjUCc4UMZ2oPQvJTfPEsFzyzFqlgz8SvwEisNN1NGkjRNB3Fb
75PCfWF/qmIaI9iq07qZ2zLfHElzlHriLImqjWdKmpgwtqAwV1fApGPYVxIARkiZD6W6YOVJzZlK
OvTmEySKzxo44NdDhGjEjlkNV6Mcgsi7pw7IL59lXmRjoZYxgGGU0PI0IgL0of08WfHjdJ6Gsn7g
MNcCOsNTked95gLCfCDyvbZDK0gQRWhZfN4UpbX4pE72lL2r7a9bIKv85YA4sDQDHzibuV0Ufcsc
s72DuZNhPQlyQ90RnY1a23ridtxlk7kOIWjtHTJNKPRQtl1kyXltw+YryM+PebL32cv3KyGDN/qg
XlikMXqMvAa18svmSubcDM5oor+P7kEtRsCP9MVP1vlhoEVYVtqA/f//XiXCJPvU4LEhl7tuvrQ9
vpvTPjgjAyDu8MEkfpHRqn+myNdSsPjF16QlOXLDdz0gcuGbVfYgcdq9hl/7ROzjqFMtnPah4j1x
jfZs/E9JdjgO8hVpCNJ4TzJFl5esBYiAfMKVvogHvogK1wqLnVzmDUxoEk0F+talhOYUgWTYInoM
eHj2DQSxGTbZXsSb1Ugt/J4BwswWWmpCRFvaEL/SUOeLtoRPMoiS+9MiCwAQQ+10fG/KvhdqSaa4
MSi/yiKQIrg0V3gBhMqhPiveiD7OhFr8Rsa7YlXBeaDFecmLRbC0hYcqRTcL5n7ewzTrggn+M5zf
3gY/5RROrqasbqty6jZ+wjOe3Dlx9OX0NOEaxG+xeckmth4XLPcpksm10HMx5VK8M1Dlr9dmauv/
C/eDcFuqVrJ/GOFpHek5crC4nJKi1+15sRQKe62+4janm6E/IUn3OrIdauIQJ+tTC341tGgx0iP5
nIMfkylbksxLcfuCi2gCYfVIMWfaN9QcN+GgE6GqYNqE7jdbamobU9aJeFrZ6DOOraMu2kQeMU7A
HTiDb3ZPGWnG5wGJs9dbWJMUxpeNVxp27+zyUfVpL/Y19nD98yNCTrEltZvWZzPty0mWfpxZE7kK
/QmJODqnPrIKP2dPQZxxcfPkruh2Rc/HLT6O2pVnDc/AtZDbfXxVF4LaqIlKqrZpjr84u1sggsxx
HU1GlBRjYdLQGZLKIq8S5TfMO0Cp5KfJcvU/5QqXjwwgKA9F9wwRsFApWSOiyRjPoqolHXcLdkLG
AYiE6NPiw2TGxaV0E1ZEPL1zE2WHLtbBVPQrZV8uZ40eu1QrSN3L4DLbBkboQTjUUAEv7GeQhEMZ
FmC9wR8tbTpzWXvIgKIPC0QT7IEZMIE/XfngRPB53wOnbsRa4+5tKjOxmj4YfY4n6R4gjTr4TYHL
7m8J3tUD6vp9CfWPHefujYdmbvqpNkmUxnzx85Dz9gQ36dIzUC2LBWN+dk/vsADAzN2hxKT0ZlIS
8+f+TfcDwy/fzqBlrvVaVXbn2ACQeEkEEq6+2nmRLKfmv++7tYmB7tacYgJ9xfv+NfPqt3YtPz+9
4gdJS+qIixaAe3JFVeN6pDu76X1G+owSfc+p9xEyk644F7Hb57eUDxk62yhRzL+3aCFV+98KwkFq
02OH50vbyLO+qkO9WwaN2O9QQVoN8yhqiZaK10KagHMB+USXXAYLOrY6aIAUGX6VRuzxi6aX3WZ6
D0tECZnxiMLqs3dZ5H7Hs7rjlF1G3Cizm7B0qx9fwLjnk3e23a3gpPB+TfFzGPebEVTgasgwzh1S
jN1TEigkc2RvL4dsNpNgHwPa6dKWzgqsy9GQ2G63mnKitVHPP6La3BPjnMavplQot8mvEqXelbGW
GtgZ3utQWNm9XeEaoV7BCZAxX0eEGWI8cSen/V/Ikumf4D4bdZcqRa0/EeO90ZGCUi2WXyO8jvGe
2pbNX8lNG390P2NvBlBDGN4MnypZejkTKzePOY9b2AQkxXiV79iNJ+nL/LCopBLX/2U4aSU6+G8C
eOMUJpSTbDKhnrPlhXOVh1Z4UuSKnpmowvrFXMlSIyn6Xp2B/4U1tDY/yz2iPDKokOM7aug87OsO
txc2vPHQBSgt2mLHIki2k1K8CgyAINz4Kcf5btcghw5kNFwsfYzKIkh0T5zHkHg/yui8S991Z4Z/
v0vVrq4HPhkyicSp2QGB8G9rA+i6sjt+d1DL4FHwJhrst4DsvuR1FL6OcVfdcw3b7pRK1VJrlpud
dOtWT/FnQ2LB5+y6v79kzxoFrFemjqKS8otc6dMJw7YZMz8+vhnBNHO6aV8nkUPL7RKoxoJrWGqt
BjibcmSjbhdACJ2ybzUx34Xly68CCwYADzRGGpUiUWaS+L9SiLbalfkoZ1lSC23HLMFjuq7T+QLr
WtbR8O8fmrcKjX8BriQeSKt56WLohZILDvRVmQQoOFnfbxk5vHTncq/31AMECx3Qkm/2oqO/jAEP
ZVqQGCfvAwO+zDRt3KVfwRGP55tuuNaJFKNLvU+eXQYCZeswduJVTzXB94pcAKIXu2dri50+SbQ3
tV4dvNGnKCNE/0uZ53Vu8nE1Yy7GKZah02mBGD7SZ3aJ7TTbzdklioPqXClsGpH6AAE8eX7prGYH
dYlJExV9/UVJn5KLbM5mvuECuZH0SFcIuBrmbDkfJ78EfyoBvAXz0DHNNtATH/D1ZD6u0SPWa2sx
L4//C6xtG2Wf8YB0FQiXXIuc0jiktQgbljymcOHkl9EX0DlhG7dImNfiMt7yiE2qPzhK5SoKvwnU
4mzQpDo+lmM6mK2sFBAO1ohjRbv/WGzDnuNH0wpUe+1tWZITFpxStFul/cK/2tCER9sa5XemhTBL
echx5eaAEjgqBxnAgwhp4PWldv+t+aOCxgG0HGDbDmrY9exklCWCvCUEMtj7yDxz+aJ0qu+gaq9n
7SpKNSrNwzBxmUK/xGeIBPZL/uAWh37KGmiPsisJ6LCxu5JwrU3Q1cEOazVeJ6dhHHGgjVCGIi2M
TXrk64r2iHmUFEIOTfG/NfbyWed6z1LKA57Sqs3yPN8PMt6zwn0uutf4i9RwFe1T5cBzOEAN2VqZ
zcetUnhCR3puhMyaWAbrhzVFw3R+FjKd3htIjvrIhzXTsSILDXjUULgrHEfWPjRQBtor4KZ28FTL
o/WUkqEU0EfKoqby+L0OO6puVuq6W9SfWTrQhBuIyfTY8DGYZDv9TMPkE/s5rQ7iuWbhmLvZ2O4I
Ftg/8UM8VWI20XPax3j8+XDqveSZ0Q5iWXUsopv16zhURHDiuHlS/vHGePnEvsXDO64bTGqNQI0v
mSXhkEuS/P/nv6tYAhRU5I8QIedvYZmaQ6N9qhpvPL0tyMJTWQ0KSU69i2YkThiaO6eIuscM8Cyc
KG2X3NlnO31Ej9u/7kck285vL9Ozn5yzQfnWK0xKet9ln6YuFFOpo5OnYdPurflxTP+DqVNK3n07
/BNBPt4Ig7rB8H1aQAYFAzTBq280dsNDmeXOMpy9zPMCvn0p6L6qT3Vb7yoBYNHPDnDKPA8nUY7/
SyhH6GJP57vWrISOcAmrwzgwc3dB2hEpftZ/9lQeu+SM+r7vHjRpaGSbMW2Nc9woMxdLb/7ymtaH
iMRWT8lQv//3Z4fn4SuZgQl10zAxuoZMNIeSTOwXl1A5wuF7Ay3dteEypaNE5zNyGL+Uxp7RyLO4
ownqKTmcXyU7ySsR2Ug2kGcCNHa/IlUsR0SjbgR07RfZWPZEKh+g+oPNZmUfroEvujlI04eElul4
es9GsJY8qEH0rpg9FpCk8dG89e16GmPhmeEVUd4YyCE1QC1bc12mMt4n1g4agWhOvL0I+VmdiGZr
Q6JcvIW4Xz1pE8gv7TjuDp85wCb3HvelnJ/jMQE5dgjQicBV/29xtbUxfNZuSS4FuyvpQ9+NwpxU
ptAMO6Tck1SSjeaM1XNIa/ga2IUGqozrCMGCjSkVvgz5Z7A4kmSXF5AKU1OMGkBoQOLk2xVC2Zcb
zTpJFKgABECAwnH3VUTn5p/q98vCqYb6W5rW4Gk+vuPvFJ89jLxAacLZU3Gw7rpkCM4sjkAqIvYK
g9EsdPpmKmFsQ+WUZkQJG5uNVw1opOIh2YQM51DWNaOGrOL2HadYy6M3mKPw9TaGNTYjT+o9NgJw
IgHutF/t3wCSALq/hw5XQdIavjjaTyE+acXZipKHPgbggPS69ho3M9gB4zpxAEVFN9LMb9IYW4lP
dD1wEs1r054HFoMkWaPGw5eS1AX1kfBHFrzzT01UB5CVlNkGH9xyRBdqPyxa17oBbXC9Dpa8nV1C
cZKAKgyEZppVqUdDu44Xwf/0hPL6z+9BVlJviTCTLBrTNKCuXcidXN3DzHSQLr0GB/yam1xc2D78
OPGEy5HRyN9FQrDGGZTVNVOQ4Ivtk9QwlWXeVztd62dazx2IcjiSZcuUa4rOZp7SLA7eDF2WwXA3
alL87vUwk0DOtA7J44vShu1mf72Q4nhcOC+2N3/X6nx4IgBg7ZOqlVtbJF+/PP7hFs1Nm9XdawdG
N/FTtfdsbl221wt5k8k3+dCTDTutitCaonNJKxf4dtiaEzQNiKgWTo4ViPeCezyOF4tRCoTMOg2N
MixlWbX+UOmHsU4wrQjP7eW/RlGvjXMgCZ8O2IhimJiiE1s9JUGfGJRcA1cp1eeTu82PzEYkJ50F
r44AzILi1Tw1gCUJdu9X4/14/9sycJ0Q+4Boqv14Y5PzuoXf+XjVjRLR2wpJtTpmwKrAoamw7JwP
Xph0YXvSr21r2rcd5+AjPDa7Fn2znVOvogijw66zaSEbk5nXxeGRdr0lIA+44Fr/YjlmJOKacW3H
HlTde23zX5KG5SaUTBVcQ0we6VUzJyCRt0eTHVckcPOtNToPtAFHMB9dxWvOT6QP7eAtkzk+LN93
6YOzKjHP5MIt/nZ/KYPu0IBRnRuO8XeTokGPiHyRmAtCzxW4p8LdUNlXiqSn7MFdznCaZ0gDdD+G
NXmiUoCN0/V9hYmJTFgf5b07XQAY/VJsHq1mhxNkmfF0LAJRGx5NpHBOM7GLk6icAP8+ut7QmNPw
+RNrz3eMVpfR9nqslhRDveURDIa4EFjWwO01Ht7pZWaaG9Z3jG1OIOt8wnIrFODa3dK9qm+oQQXH
Kg60G+WysAeUMkfe+NQ7EotO2kkKCue39p8fK8AKgCOcz+4vOZY2cGaShTOLwsaimNJ+U3FJBrH2
ESYUbyRTmuwHSbmI6o/mOibeQWy7k58ENU33Giyofqc258dRS0zoFD5wwto/4gvTwH2pinjAQPpT
+RWE0GN5btfs5452NbVsFGR6U0QhiuH08xpLbJgOeAisRuZHy5cumF2apXojK4hnhMpOfgJeoKmP
rJZ1xAdiCde74TTJZHKPJPogxDvuEr9LOGAb0TaF50KSEPwcGW4ks2Qzd68kpZrF4MYdBcyfsa+S
TzHzi1nAJHCA9MjjHajXU7z/+Sp9dBnd6SIpX202ePQWjT2Ex4QugqoP5QIg+ykokhF/rY7giNfU
dE5RF0hN+LC6k4sumnGWcthfdjiBDorApcVoKVbAB+E3+W5ylixlL5TS4EFTAnZAEJG0PxI71o0z
TPPwoLmOs+Nq/IjvuOLcGmEed+upuqvdr1vi+PPge6pSCmOfdn0xV0Rar1FnCilIlVNa1opj9aoK
yKSDm/DDOC2vNuH641CK77bwcbZMDQaPuIO12NVBwSsXMcx+64E9D3yarZCeG+b5pVEEk9mYimxn
0Rn2hXHWu56ONZvptIYkLk/x07IehoRDRnDRIs++HVXJcJYY1ZBztQfMK++pZ8v+JoUp/5XNUDp+
Mtd3jUxQl1bboGCeAAjlqiPn0c6CrNnTB5Wg7uEheZl0cGnbBLFASSpj3saD6ivSLjpghZDB9wlG
EWSw1EpNg125GfPQkMoHLevziVPaTumGOmpnYhkVKAWI3VyODPDRAquUyUrzS+AFJ2R8ztruQHwn
Ly2puB4L0/AIBjSUB8q5NZlWaiLH4oVy2je82ahnFsDbSrZ708n2KfpqfrMwBu790ZXjkUdH4Wd+
KU+lQo3j16mmhMegdc6VDekobNh4TPV+jJ0+KKjC9Fb4AaZEw1NmIwPxhj3x6++YANI5oXmxkB40
Bui+L9eMe8UDru8Bngb+H5zmLqdVbVHw1ffSptWxeRvCPaL+B8TZF6ADXPAo21YIl074uU0RdpJF
oiCupVim3ynb+iFu9v4+YzR00z5tJ1ityt1G3MEvOqTNnnesofvys+B89h+KFDZ98pDh2rILO1S+
CBolN6TW4EV1VL/aBdraMylipoutdKFQfl5I1pgGiOFSUWItsq/Vu6d6iktxxmRlT1+JmnTxYlq2
6JycN0rsvFWctCy75U6IkPeanXV7/SwsCSCXz9knlkUTg8pNtbcpY+30izybAcjtRoGWQQylgx32
Gf+uvZa8rI6cjE+4jJetYgDka4F8KRLmFO+eDFhEuzryCZRIwPCv4GGRTm0BaxmEkOVfbtFYgbTX
nUrBm4BSeQrmvbBTb4qoDIzidgN62phwtQZBhmLNf/45RCTsZcG6s332UNggD3y6GULABr2V5TW+
lHLJiqI6HZ75/MSmdI9QpjvF+OVameGeHx3T/44tel2FSu0H2HQoHT0KSLMWbKZMfqkbpF9p/i8c
9ScKGTKxW6qmHvjUAMaz07+edJA4gwighZtIQBzGPvwA6RZ+bWz5i330Kq3kAhCQHZFgHNKfHmkJ
DCtoJ83DgpqqeubqiFav0iyTxO6Wveu6azu3o/V/xDpI7WgSKrvVZa4lB/ah1kPDsuIPSG5NX+XF
VKnSxh/k8hbr5JYuEU45KbcjDt7fmX+0Cy/UTTvS1y0rge+Q5Crnigt+atnVKFcauXIpusrsV/gp
sCg005tWJW8SUMVMt2tWA0zjVhYtX4bXgJ6KZRY6wg0znQo27WCE8kGqW+g1mZoa8fpmeku1AyqQ
JsZGS29h5mr1VeQ74kdRMUPeXk1+V2Enbs5C5HfEi+uvJTbfcExprI8ZMyVtAhaMcLbu/9RXJ85X
GWEjgOt54ubzzcGcjf2tButx7+6BkkvIn4RPagjFVusXiQ8q6i6N/kc8+oubMdpjVqxTKrQDJhen
PRkxK2oklownTKJjaXP6Y1IdS6xENOHHzZtzXou+G3IYwcrO/9+48yFfVQkRSBZa11LKB11zckMj
5JfP5U1C1+3FQ/yksfYb1fmTazHIsfKJkYtjRg6gfiOdu687VO30duvvO0T9fE0AWBvTWQBhGsmV
KnaBeNjYViYKJ2iuMiT5vnLSq964Slt92XnlmNijSm7oTgUWOrcrk+FXPTDs5FwrMInX3qg+VwK3
FVmjMwt97HJikJLzypHs88jNuVr2BUSlD8E8bILO7JRYMInG5izrdkT33h8g+RqoAMWePAW6RTKJ
+zHtxEInzxxI7c+YN4F3Y6HgSDQh0mmamRS5zPevDVGyfNt+4lGBnI6S1dvFtC4YzFxAsC4yFMhH
niEvs7nsOFcZRYYe8LcfCvyrB1FI/BchSfNc4VdbpkQgpXTjZmScilAM5RlfOUvDjDvNvOy+1z5d
KPCgnW1qN3I4zbxZ88lKDmdV0naiUwfvF+KathJQLl6znZA+JfifNERMW8chUFdk8FWeQgJwgCP9
ElrwI7mESqvjtZYo0yh62nIY0GlFhnn3EdOHfZcv+YinevKr9FnI+1G+ahpfONdoO0ueXGY9Fjud
JG77OecO4ZvCWFs2ZwUs1WI+WfGjGS9rIlNd3iBPxyaYwbt0B8ilg1s1Nqe8LQB4jGvQMoNaLtkW
52SDRSEVzUOSRcDyq+E5+wmGjKYviEmgLY6CVp9CmoDFt+dvhbc4olQ/+jRLdclrNPKx/yo+kUho
3oPgkUeV5COiXM8QqKF/z8Fa45W1Jq4padZEgFAmC9qZj/T9pMVMfgC/Nya9yCklTDp7+gxlNJYh
93dkXZ7sJaPDjhQyIquq8ebvtdGvC+TGIswlzmqVl3TMmIvOvCgnS32FIOSLWQfJvrfnVOG3Pin8
JDyrMzdoANqmwT2TkBNtJv9odELI+4qhOFvdp6SS2JQ3842SSurA+RQ10137WeCfI/wvGZmYaqG2
xISNUPXIKEuV3ZhLALkz0RtdxhE2VMITvA4+31wjqvv0sE25O81/+4wl5pmxr+CL2IwvKZcjw1pz
zaI9uTr0rAdGxZvUOixGfCQ4VttT+Xopq4Kpz4w4k3eWuoSy9n0aH4ALr7ZJB+m6RDP4R/CBeg6L
NFewK7kRfVh47TZwv7HjyymPZ9sweOMMYvAjmgD05Yc+4W+AsVtmtb3wxshOKkNQ9qxl1vxeDTci
E9gEZnlPQwhyAnjH6Bhi4E53pPbrPUjghoAVzvT/yLnP0oxvlehslkV3V8YQMht/63bFS2gxIbSg
VnX0nFjprE1KEzhHbyb7KeyCrtkQJYtnXfyzvPWNTMT9nnxXL9Acg/xQ+RY6y+30umeaVtOA9qjW
lI5Z9Hh4KFgPbUJ0rHpa98fZl1RoKZTxhlU5Ji6r5pfQPC0KVXfvlzryqVEmQrZvNH0Zq+DNGAYa
pVt24CT6uxV2xRjI/yrKDmDImmH4SImwMczWFL/virVQtT/nbr8e1fxGm5ioYvfUh4eUYjfXUBb8
rlkfwwuHzSCOJg9QiaQk24YoMjCx3ssBfxUcYqOl8Qm2/VIAGapAk6NsQyosvGJkbM6hcKIg/awg
CEUAhdo0y5kF4mes4LY4aD+YQWnKbZ/AQ1kA9rZAxeojmZP4O+Ygg047SQABUsAl64mf0tDYZHYV
aXQq9J8jc+QFGVoGFJQlO2P51S7rC/xcFsueCSgswI6+kRjiVYGXJwzR8ljr6Xf4Yx2b3viWlsem
W2VpdDs/o1vjwc5lMiJQXyMBhbxsyY8dS3fmTgiidP3FiiL3YQBKeVjqbzx+uVW7AG3SCFolXrGe
8mVCCc5S2DQ+FlJU1DAyh/xIK3fdADeh+CdyB71ByYp0FjOCAQxaqmEmWewM5DHNOG3l+Kq0zjfe
aqvmtJYmv3cgLIFZ3fEnX45tEcwdsPYB7T7BmW+b2Qrp75Di6ww5WLOU8x8qnhX+OzgZV7N4tNrC
bIJXB17JbLv9CDCXAJdAWc6N1iOasmufniko8WGEwiTIPZr1dj+MWDwOSTMNVORwDTFo3ovabFPv
wPA4bS/C4CEa6GyQLPMQEPu96MeI2viyk5QGevUbAQ03BbjdWDihf9L1oPM6Q5lGHXbafYA1C8br
u8Tl8Kx+lycosOYb6OMsGZUHXnvn7/fSTF4YWF8ybZze8eerTdS4VKQDgvGm118QaulC70eCrnzI
rdfSNf4fF6NwxPsAIQ7TQzKo62LCqWlvXPmDHHStcM6SV0FZPuK7JVGgm4Sw8gFyCmius3YNZ+cd
wN+5UUeCP/D0Vp06CdNTIkUw0x1JcfRUVJMpkqQ4XmYHuYcaKo3WNas8KrwRh99I9+RcuItKew02
yoCo87aHjc/IMJ/D5MUSW/Oy3HVtZvUsK2yC+8EMTdGcJgX9qWkhH8CLmk0c9v2F1lCiw7fuvS6Z
K0AUsVZe+AyMSFaKIcDYw3tgXRiM1DDX6Fp5oCijPo9X8O+jyR6YKNOcBQ3udUEBuW+paS2XPdA3
lhE4/I0K96MYpls+9+QO1xMEFVPzF6pawHRnzoFS1m3sCQ7QUwPx5bYt6r/bq7h0x307OtneJHut
QTwYIPNNKdXsNlxaSbOXUjmhpiflMjSV9klWfcQ4tcqtGpmNz+qQcU5hwR6wONwnqRGnnClQQNyr
pKrAQgP1BwE2YgbcMq3H7LOHF7ULXpA9aRj3AvCNa5Yo+Amnd94ugxpbl1N6QT1WbQaNS9leKkYn
4U8LK+NVW1AWhbzRcnypYL1yY3v/UKZCrJPMxPwQtoIIJvF8ymaRnp4+H5MpmMpgv+wrrq7TMvwE
YwmQP5XUWV4r8ydcHzaGBgqNw6/t2+1+l8vQj89pgwYw8qAWy8W8DLDU7+OBV8YS5qtC6npiCT7N
XAhMz84TQsfOEes1glSx0cMNIZXCedp637EKBAi8NGB6t6oohMkesqAt9i+EkcFWse7Ahsw1HW/y
3AVUT8HNiQ5rP9lq1Nip317Lch6zaG/KsHAEtJPUbRFo4QHv1HldtCNEPUpGpS3knRWnsP+QVmUA
VriJMeVZtdes5MW1d517wWDbhQpYRueaJVOwVZ+NRPAsHSc4DNASB9CL8SifPj+29CoXX3/B0COx
dctik/1FLtvC3dxEYFNXj+PUOjqI/2by6djvmTmxfX8Yafr6Su9Wh3wzXAjpnRhd9+Uj4MFFb5XJ
uBNKKbrB4mBZV8pgMcps+OzohOvpSCbRWo44Y/eHed+UrIUBDjSZ3tlAytLNj+FOnAV9jadyUjJQ
nN5iWqp32Jcv7GLR81HtAWZR9S6WYPV/KA8iFU3D33hVcWTQdA8YBxPLB0M+uwTC/ppldo4yHOkY
M8y7X1P/0UiGsb/HLdqaVCjez7x2WpKyyzEcsO511QVDNtaZqs7WiU5dbZPMDxpEP8QhxgAr177M
nU8kml11a5ty/+ue8crxMJl0oxQ0AEUmI1F0IDQoCO7fZbMtLJou3jKI2EMk9ORDs265Pflaj1IA
23Y+8qsZV5EL9BR+G78rKPf7bD5FVtKNqYeYUbqsNX9M/HGQhnJqZBtt6OR1Oft/Wf1H2J11xRIf
HwNMQsbMDzDRCTleIpFAeuz0mnJzXZGOVA2duYgekSEyq+OWY9ED/ePuawoD4FygZVM0wfS1kfuX
nYaIXnryQE+nxenBq74uwUvP8LYx9q/8SzlZaV0qIoZdefhXg0J/nd6Smc/8vw0P2TO1PvfKjovg
uBnyvTkT7tVMYz3nH9LhmiSFPsyEjoRHGuIm+GD7GFlULWi+TOkAnlo4HzJwsBm/PbZg+affLUx3
M6o7ETMdzWstsPwAaaiFXPnze53Y/xH4FjFEi4hGd+XR16vTYgX6+azNq6ulIo8gHlKVq2lvyPHm
GH3S7hGTGxZqy10CiSAQHSiCViVh1QFEoDs1B+AoYVnr8CJdHHybXZUSqL8r/9whkbZm8nAmBBZp
yYzpwO5PrCD23dGERTCSvDex7VYKu0NKyJu8YxFPmXqBPgdsEGSuO0aR1oIiLGcfUdGBH92i65UT
N+xuaYNZG2MxxDpOhV5cJ69MX2appGG1PnVfs9k3NTvVJWMbXUOvOwDTxeZh3ExYNhfpSfw1OYug
jM13On5l6CwsK3/OnqwjfAqAQu15sO+u4V6Td12saaiJ8tZge/k7HjhngI4WgWa7UFlkck2CmyOl
Bi7PFujrNCDQryna6WAh57tzqQi7nvI5Yd546OsfHiV4eL9HyUwQffLftXfvJbm+5OG+mxCkZzZL
87q8BMzZxwyxRTBk8oWpOStMT1ZlEQ3YO7mQHD4N8E2dKJj4azaR/HGYoP6WF1F6syM/M6JwUhCP
a5dFMlGi3re/t6hgQyF1cWL4WCNPecP/tpZMVGEDDIJSELsTj4YdjwqCmXd0vCTl+wbg5LR7/zeb
yrxJdieSYwsEcpvXXUw+7lNyTecNSjerOusqeECdsdxPi87rNpuZLXghdVDT+WfnKs/Z5ZVSSSwO
XYa45JXMOjRihztf+dp5F1bsvIBYnzPVB1H96SHMf4BwpnzgYp8ArB2ki9bgoa8292CvhtS31RPG
MEoFxdzAPkdUp6ePTC5XP8SKImX2cOAUG8a07At5V4SBQZmGFctXjO/+rebCW4gUh4MDpNMoAJKj
c8hGTkixHn3IKtIL007Iwp6utJGnQIsnqP8QL1vxVaGObNzQhJWUUwguY3pbWVor3SPiT/LSRMDz
zk3kdxxeKEI5U2s+vCIZBg/eNlZ3V18dg5AUyHcLCZCvTv5hYdXIMsGxy6kk6MyqZuXr1zDiXPa9
mPqxJ0lX92lkCGeh5b000INZXJr3/XwqHhNyuJW8npxPJapaj/CEUbl8KT0bYjQyhppVGiZnvMoe
agFuGeWtuXx7h1BkJ779yV2uJv3tT/qhTOjMGi5nuk6S9gprQZtz7N43rEDGD14+l9mROc2KP9/y
9h77gejBQZR6Bc3cwCWXcHeBd63vlvAQNhYdlVntDLATHnBa/Q2wWU27yxYgrKwcSiDhV/6UrdNL
5ig7ypfRD8A+AJUWoGqXtuv5w4ME42SRaWdVlrUDspEjiDNic1nC+Y26p3oOQSr687xEH0n2kYgX
7Nbrh+8tBb5Glg0/lhnoqwjzflzPUhbuWrS6hcyI/Z7E8mxh/BJ8g+h7ycBWGgZTiFiJo/xNKTTT
LpG+GhvaG8+841v8wMepNSu5OfAf3qVT+nBzV8Ena6Op2kBfAuh1AR+ENijZ1vl9vTMGRmU2DoTe
9rRxAMtGXOTfoIu/IqKTaZowGAsFXFsVVNg55F/Bo1ZrSbpb6cXyxgxUaNif+i1bO9PM3rSZ9N1B
xb9+x/Kz5bU7n7pj4+j8dAneKBgZWfBAW5TW9lLwYycjsbeoWsCr0h8JtUAiaTVq4zHYKrc8ah30
ngVCjW+SRTMfJINhh7U0ZRbXKcJFoc+3qyUI+liAVbKneOo2uU+XekjJ+lOs6FSV7YQBW8DB7Qdb
leCZVM18DLDkxiT26TrODbYwqP0YbgzSTy2251Jw5hiyfzofaThsO7tBANcavjE8w+DaC8MsYCnH
J1Te9GYkh1BVCwmueo4ODHssbFQGr1Xl7F97fGUUDGD4KGn2cbfaaRJEMglcwcYJJ/Ow8VpAJplU
4TpZWnl2i1g7j4pj47G94Ei5Hz3x7XlfzPMCM7bv4MV6X9jfLAu3F1YsWQ0rBE6VpxcETfwC9OHz
WX96jqL+XfVbCDSupA3U17SIyW6GWYLc1svm+r9Ke/T7NAN0AcnpWNvWrxhZCVJYyjuoCjs5NjRa
sjurgHGaJRzFqBQtBzg+RXz59nOrfUzraR6PI7NBeD8bkgMKmTmywojrYBbpnSY1paTW21eH6wxu
n2ytibX20KZV5a06UFk1cdHUHEJpnaG6Y391H4LoHA6A48RdBegsJqoDjU7TNmoMtQTwz+zDxWB5
qyGPkIL1INIBZyhB2qqSgCBr+prW9QnF8+O8zpgxKrz85fi75RHSkTI24D4xFQ50e3xYezDhlhdU
+ZY6sydHl4xp2aD/vsb83snbeCMlN+/PEjXW/yF1FeXWNIoMxGShJtWpFIeakUbElguzEzEEon+3
4ROrcvqJ53PaPunloHrW/wZysLvW3IJl+CUbUIKAJKnH0wK+YdWPS0K1J4jzqMpujwUl9R7tOJXH
H6/6j3kV00w+FbpXzv9inQvcKwOOQwYz+BrJQux1jK3FHintInFeQfxqokLS/Es9c570UUf+FsTm
3WYIfh8H3LdrcC7HpMq3/LyDasIWs1JLgWH9FoDMqCbCG28S8mBek+j1swIPriMolD2de8+CcKA0
kicA/Ila2fyTRdsODzdXCAQPX37elOnyJuHQjr9GSkwkgTOZBQwqUQfP+PUv/hFl+STMcYA55Plv
IXgWJpU+H62RcqkygidtuqcvvITtnrYV7/8zwjP6IgqGh7mUZ8YuupRN0LzsO/IfilmdhQVOMBKN
vt+SrZkio21fJ/8znVyFTokvLF+btyuhvJSQxR6mHpI9N8XSueqBlx9aLQOzsh37wMuil7DJmGhX
BT0t9QEAAVQTp66nBGMRBGnyNoFYQ7ed6ijef6cSjLin2xuq4ngYD2UGyvyTZLFqDBje83iLD+bg
eDu0d+PNGibCaE8XDCOVUQl0G2Ipfy1jYOYPs+E1hT5ZdXmqLXPd4dcfGqxUSBlPB/cZKTHQcrb8
HJLXkr1eMgzuKs2BURlalxF45vBsoH89EgZ/X1Vpkz+Ea/jeqO2wGKyBvY2MxmBQNPED5OBXaDyc
xOCGbjv8KsGiNXCqzUidHmOlHkCnDHWMSMStcpoJVWQ+VIzNAH+PAGkxx5Tz3HnUtwkY3Bupzkwg
wKwf3qLay8PvJpwcJyiL+2ghOLkVejcHVhHXKO4aRHDZIude2bIdF7Zs2hUUw2WxQdSnF0qg9in6
71sy0092pRUoggZZ4rtfEpNSrHk7RIjuDIszoTZU4H+5T59VAaK0cqrv6fSr01uBd94Hn2SI5Jpv
oEyqTC9yBeCADoisunJnv/FlTlseGRwBx5K8aU/3Xf/Vk3WDuvTjdcry7faQDMoozXj/7z7BXf7f
+YRwRF7vpSn6PlMbu2saarjvcpfEyiDi//k3UiBct9XqusbvdH1uHvyHvV8tp+D3Epcf6FQ1BM8W
opQ0OG4ubbXgdW9KO2IJqewUBqsXgdnmeg18l7d3OEY5o4BkB3DbPejMJR3LtI6maksI7jZ2zWt3
kza8J74Lm1cVhFspI2juowQ9HxEgNecqquujWtITZ0HgSmVnxXlOwRmvk5o5lTXb5erGkQROvfsh
BQSOcMY8EUpX/+5GFW+7oxintzwiPzcSzTzffgMWiMhZY5BPfOhJRsFxhjbv9irNmQmllNNFv9bZ
giwG2SvKmrc6618i+C1Sza8i+ByHae/L6oMpeam5yxZZWCzEoSS4Zy61TVl8RuAnCrcrR1rMKRD9
xlZgax+kgwOwtVrEkNQyLnppA2FwpAsM+mLfsr0tO5wAI0vFizN8T0mGNWBXR73H7+ZWyAh3C7h1
3bVvK5DPGwt+kA7/NiQRJtiLT5i/ZmsBsr98SNfcp6MCKqH5kd276jsBjqAJqEWJkBkt9qu9r+L3
qxQiyNHMhBgOOnM+zrjiK98C2A7Cc64knNMmEGs10XytNtX1Ib52Ef2q8W7PkIGynU8xybgxt7Hi
ixI3kYX3FhduY6a1gMNA6+s7N/1GTlrb7tzVNC+Hq9JO+UksOb9Pz5QL2+LDpvL46vc2y4IMlDEY
1OzLe86uY8bUO4LWAwSfL50IQvfi403h1E8v4V98venIZDqcWHFji1TZMgEl8B+xvRalmWzrwboW
gEWuijrx8D8mjy3hbLQQ9wOZFk5/KCrTUyyOg3/8MrZysovdG6GBkpipatZmEE8mNF8jxlz4CdPk
XdqvXpA3BaUuzKEZhxU+eAVj4kWtfcN90bteN6eCQburemKOlg2a6E7Ped2YSmJ2tRheb6srbZZs
xOGMAbTmTXMRffG9A38Ct1jisdc0V0+dn+IAiPNvvIzVSPxcm8UjIFhAPiztzPIlcomdQq6REfj/
r1hgp6Z/ngdqqoj5AkY1Grwg0wM0govxJwARGd6NaLYsAf83q40/JcU9IuG0rHLw9VumCzplObAa
qhrvjs8n4zkso0Wllv39jUw/dzaNo8Qqxie/d6PeyW4d1SUmiS15ECqeX63xwAPzjCYoW37se8eI
zkCxbOVTRu+7v+5YrkDNaU/znGpIQhGhTG1xuL4CA/rbiuj8tmXzRdW/anap0U8kPtg1uqdmXT/Y
XE6k7o/+EXZv2rKWwq/BPoLd0VRyBspArj/+lnwvDgxJDtLaGqP7p4WknThvMSIOgL/IT+jvVISj
LfDrh/mTVF4z6lLunS6Z2VjOAycAG2efNvSdCaLQFVlCrlE1Lg9pnEffu9WnM1JhuctgQcQijqgE
aYOuvolmgKQvkQY3U3Ds/L+smMqHwpImqaL3E7QrtiTGwXod1gkHtM4MjALO5KBjbwI20V2D4q2i
woPieizbL9DnOK0Dh06JFzWVydx/nxc0q2CeS811gLWi0j8DP74QA66/hxbIMRT96U4XUtyAPeIo
jfT9TDU4X7HaARFAi0dAlvOfOK/V+P6pigAh+guzenF8VNkfSNH5ICjXv7V0fjTBJXBGGRdil6yi
aK1byt2qEhW/gFUultDrkRdZEZlJVE1hMEsiNebrTcpw/aXQhHfviJg3m7w0iHmDkYJedqUrmzZO
U/vG4XhmGNvCTJIXR6RS1yXjaS3dbuaezZXbR8KN24RUraSHX1QtncMcd/qN+/FaVX+An3iYmmUO
/my4jkhXsrFE904ex/3k5TLY8/+0PyA74GzMvdGLdBHlloH8Iq7/8FcbfsnYIW+jcA4Z++ASPltM
QJXAUnIvYWZ+1wAEgx2xkU5gDM//YgR5OMBqK5WCMtGXgUShMrH6EZgjXG5Ci27h1TiBJZX5TPY1
rD844w7g9qQ2Twj5f+j4C0fYMcHOzsE9GlOFHo2xtNsJU+l8/s4pylAoCdfpENr95vlq12CRMOC0
AQa+kIU1ZXth8BR7lqfaDi8x5ydD6zqYy/CCVRkauk7eYpmEZ1Y4MP+aJfOuInLT4PNRi98GFXKi
hvgzTxjDK+FBty9rwnocU2Lgnhnd8De6a/XdXzCudrqU91rGDuFrkZhOCfrW88Cv6lfhXyumhgMv
15RZi3PEgdsc07heyIE5Aw/YfoB7exJZdF9l4N5XynelCivvt9o67W8Wkm6VHVr1zuXJw4VjPYUT
Z5LIOfozWU8swoNVR6nYAls1su/XtRLRzbo7IbuLi6iCqqPIeLseKEIYwk5Uf00YkFZSCDQFmRqR
sFbQ+lf0cgKiHnGBs4Ptw/tRcwL51GATjZBgNxoDL6X+vPRd0sIzu2cDFKGkYK8x+mORuNgIhyPO
zKnIP5VBIS9s3Vt+VChm+lDWqJsx3CM0DQzmnrKK7lbQlSSF8U1Z0U8e+SZQWM7vtdnuwo1U2VEx
vw/+ecdy/C2t4TmfZjTUzztug4NlEPV4RBQlsgpH3nkfWXOHJZj/ajKjA+WDd6OUykHPtrvYMv22
CED8Q2V6pNeskNm2YvpeTDqFIlNv/xRQVQ7N142E2A5tU5y9UOPq1mqY54yACiqdOmj5Izk6ZqzY
K/ozBzBjawrUcPIfUqBLMsLvJ0is2W9wdzJxCVw6XQ2ASY/eX4Q67aYVYrg0J6m0XVlP1uPxkGai
z1HBGB0jIRpKX0Nap9Meaym3/icYaVJlXEWB+uCoycNYVhj/53ITk5gqoebfPmWDU9pUB70TeoK/
YUnoALxeKZk0R2/F5P6AeAbZ+8gLbt74S8rgv9J2IDVToZFIggqShAiw10k5qP3mbHFwcQ9yDSgW
sQOyq24MSJrYfvBPduRInP78Hz1dTStiMg3B+lwwHPPRmUFXItJLVUByJGZp6McbvQ/c4p8Lq4xq
1ZYaWP/c/a30+7XuOd4HCyA4l4zPHOw6+Sgvqj9nEw3VRKsTZ8c85mEEMByasJ+pL+9wMCvEvWjf
Ys/Yh2irBYHl6t8B6RlNRDPFzzwiOU1oqNBGcL9BqPx5ZI4FwVg7ZUbIPWBMR0kns51/W5nc4NUl
Md+5F005ySA3CeV2gN7qZSQArqOV7J8gfTyVjI1LqyHksb0VnNOyEmHczPEtQ3nVVOMZDu596g2U
I2dW4/rciPh0vYlwuGvXLP/uvw7RGg5Limdr2JzxGnbi7565HenXeNEbVVkwtrPObI1rvJdZtUyG
sCDrqvduCAN+D+/XVyvZQAbvhuVTXC/bgpRUNEATSsnJJxDDfg0tqJE1HJ0YhohENI1bcMwe5/jW
vA+7fGRFn+N2fhRTB/RngAxzC/WUuWr1szBN+QDm+2D4vpfn9SHIoS/BbVSTE+72PLU5nmFbcDTU
J66qqgPWOUtxFMZ0n8Gv1LUprBUAZ0YuEzgfifulqj6Wasx6NEyjYadvXydUvZWikgZCf9v+BRA6
yz4ehp+y5FekYog8uplP2VYEQqDLV7a1/IQGkGfi/1Olw4Mw/MfJh8pG3xDc/B0kdtx/vR/HUj46
7iM0ssXIkU2I2ejifhb/cR07/8h/+G/W0lwLQDXNmUN3R3PRfGF2ZOZLsVVcv2fhjLsUV7IzNMVg
0+I01FEKXkvOqFNlPLjj3KhkOVuUFiTFmIRvOTp2TgVMB+UgygPd651whtZQQmxHY4wquCVyfCCf
PvHMqx5X63QDdvErD6fxbIYhF09nizSq/dME7rno32ulkpl8fNB8mgr7edJFVcYOKvH2aDPOQl1W
buJIzYDvChOSaRtvE083lRJsWSHZRtr5yNu4HEbngmWTbz82PtVQQkcioph+RyCbWJcSdbaLTeho
Zz+jkSGnlIVJdGI0dErjuzKJkM9NcJz410Yx86/qXJg2LXZR52dmX36vMhm0rtxEiECiVE1CSA8P
wzLyMbxRmO+8kbqrFw5luufE/t5dsgsjRcB9PH8b9ZRUyGJFx2KgA33NY6exEhld2z/CJztLzb89
XLTlwGy8LRVyylHx8MGLel8vpLvPvQpTwC1UeHaHnmRmUA+hSLCHPAygJDxJcfbmKdrjJDMeRjUR
jR8BF9jc6EqfnPk4emv2qdPnW8+w6vjnZMZDOLP8w4KHrzA+pveUmX9eAtJssnFqOc3Mwtnh619b
EUWln5I0L7uA8u9wRGMfRga78N6Xv9vRyu5c3TGWheAC0WafIIr4wc7n+edeFW6ZtzuIqqffGRew
EAw807zwgMTdL7vfiPTIKRrQrVJJh40F5wN/EZWlnqT4OibyMgIhKjiso6lLxv89IWFt7njz8tfo
cSSF9Ym1dKxOJZlg35+vheCt9un4zlKiHMCn/zujSsCgsa5QPOfkl2Np0KMMu6nd1OATFAgU605k
adf0ZC7hKPAu9uVYfWc5/uo6IEQYeiYTtvMzG7lUwryS+UV9+Z49Ghe2uY67B0Ux61JoZ2fiYV52
QwCAfSSle9kDI2X9GadzT1CVdUJsfkT6VuKcEH31SKWnLMrYHeI8IpbQzA4FCRE8X7y5eYy2GEpi
4Mei1Es0KFJ0GHFn5o7tH72DK2rmVLHh4+Nbvwux4ykTL5toPTcFf8yreyA8WtKbCza8Ty40aPHm
ARL61sLvDo9QMuBaVI0Wj6Ky/MZg8xt8s83NfFpkfI2rJI2RyX4eyeQfQxVS5BijE02MWyh3BHU5
g/L64gsCjvGniHC5iftaucFJdybZk0e+SSf/9YiYnNe0kg+PH/kikgdQfDTT9tiP0X0nS1hWJ8/7
ZnRk02UKN4NJkF9gVfu744GzigYIo8DpKJdxMjD2aiyBHNtreRZQss7+x1f+JR4oYPsp6It7cMSA
GmG0CdJ+1PBDKz7pUgJ3V+qRxS8lPEAgy0YwK6kzXggL9zfbpgVhZySKUnqd09chfVvQGB5gnr3h
cvzk2e5coK1FFeiqdx2KnKxPuUJpngtqTF7l9NEveoBREBzCezdsCSzCu0+wTIUzWyhgynYFRdwB
Qb+0tDmagd5sf5q8Kg3t6DHaq6PO8so8UtR/lV+oHTI44tlPVdJ0f5EWOYLpl8l6zwL/MHfNw/li
WGSI5/FmdudrAN+wiEDJRdbfS5PlWMFcfJEoIVqnwm21nzldSFMsFXn8gGFv3pWhIEPpp0GJ+Lvn
MpPCFymFcJh+xeISDLS8AJIhMKan8G1S/Rpur/hEYy8cB6tFRTgPrNGml/066Qq2gZvyzUuOK49j
x9L7AXxkVIHg1IHBuGOE05YWnidNeDgaoPEnZjZjZNVWOyYqQEIOtOz0NSHlSDE+6qZz6Z3pdOc1
sMt52xjZ+tA01r2KyAq/20/YyfPQnyypq1vBe3k8TOCCRKOsTW4Uhs1OKp6tzpyvJSwVCbC3GL4Y
ULth3NRZm/qZsQ+hqKAywa1N0ZRSAZgeEfs2+3YgWAkWkZrjPo/1JYlwUSBx8bbumCQ5aJXaOE7X
5QBQ0gNC0JPHzlZp2138lQ+iEjhJ/qAYipOwOP61CyKf0lVBUywJ9FJeFChhYOajLWP7b4FX1PLj
gRAhdFmB6nAAutK0+GBDdkurOOqeF4tKeR4Q0dBd2FMcA7ZuMRdjXdjxuC3uqrtjGsKKnXJ40blz
7o96i+dYT6oC3KBqjYYtc/AAEoTx1oSIZWcGry8RKVq04Q+BBzryp6qgmJGGRvWs9tROhegzBpQY
Sl8K858WgxUcIGn3ZeDTc0DyIzWKRh4gUIbBM0EXAEQJcohRmiqfxJZHrAE5B6+UY/OgvjxSyzpF
Uwyz9WDK1xW8o/E2i40WVrrW7Phq9+xcDgXP02CaEOFeTS3bbz8oMKGl+/L3syGigvOcZVBhYM/7
xrXqbY5ngYEkd++IpCo0IzFZOSNx6ENW43/eON5jAK42rtVhgCI81rhJdjGq5G7GIYeUtw1EpVOl
byqhrvJ6mVxnOXipmqFkV1GyC3Cx0hKN1u30VKDDbUydECTBI/yXPKR+Wk+F0iRS/InlSAFwTuZH
TKGW6tAg31sPlGJ+t0kJYWe03dUHc1MPeW1F4HkcUjTE+HFuq3ZQVs1QdA4qRqB1P7TcCu36AS6u
/JN77j3k+bXwnEfC1Jyrwjr0/P8yQzTImINj2BZelXOB5REaqI+RxNs31nmOLl9u8gk0sNMgLP0s
fP80CI0zCK9QQ+N7CM7RBJZxaiXdHqQv1uWw6PFJf2bp0Ag301wVhC74XplurOnlhQ6vgbhocn2n
rSIir3WaYtTELQd6RsNbNo7AE8I7gRM0hfIDGL3WHirIbJidaKQmKnt9rDLy3NZgXNgPek/M2iQI
9L3pwzEr1bq8WwwhyLOaHSvLqNKPyI/9Va7JqGrv+gpG2e0bwrGX5Ro1EPyiFSF40coC4zksCM3D
/FHkYOHI6U9gesuipwQSdTwNqeryo1xBS1ZJ5sVwlWGd/vQpyEWER2IRHNLoiJytLXzrwUnjOn+S
9Xg1C9Tsm+UXjj8jyNrBsasYXriafq8aAjMcv8iHHwQRr920H0QUTswbY379hFkrh7B8bkldHJtz
9r8IHmtiAkmTytsoqDh0hTJGSc+bUMibJnu24JQOVerkApXrmqh7mGKJS1k68tR9V6GEfio2muXs
W73oq+EXWH6XDB9UP5SknqLlwvygfGRCxl7xLXpwPSCEa8O/53mu2HWpDk7Nql0SIegGRMD85iDu
RVlN8T9tLTt2b+mdVazcFYhrH+Ai/nyb0SmyogrpgW43KSmflMdBpCH2QjMyslo4rUUHWDjQFZkH
TWxh5IXA0eqveQAUG8SqL8+vbyPZv/2T0HA1gUAWbaJBHCDy5m4UTKk7gcFCM6OOV4/WcNS5iw2r
RKAYjNhmpgSdwOa7rqfh7Jyy/OuhzYNyeurPKrN8qo8OlvazicdqicpBqFnWJxbXn1CLSMusHHFU
tg93YHBpTK/VpPm5zbmKtUvNVGou3ghZEtyp/aRiDeYM1NLAWJC+zBrJ+aEzNed/fnNrr3QZXb7J
8A4BbHkrhtU/WhU9X+u77ZxbjMgbCSWY0A02l0oIRPAEajeXPQHfsd8ujkxIMLZtisPRWtBlelVK
a+TEjQiVyrWzskuzD2AmTbf6LqNYGri6iQRD2WSy/8V0UyfkL9mX/8xwJ9+kPYb0jpVk16/Nr/0B
/YpKtwEHRyAC2J2Maj9u5tLFRgvItb1YilsTKf0kJFpCuwiVGBz0UOg0c7BdsTGzabtcEvNlqmgI
LloAt1HIB5R7L+7PT6v62LZseZnO8+GBOLeDrXtR70Ywspd+OkxQIUZepwMfxYgf+hdMYn16jmmG
J1sijlmFDo1JNyScdJT4KGoAO7Lub/eFOKyGnraprtr6aA9s+CgnEjT69D1KLfnGuDueTeI4Zus1
zGQ1wSGEU32S0RUjcluM5HasGcG9SpgOfCeD5qY4dLuRtKMFEtYbj5SnJ92BChKxxM/7zJYVT66u
ULPdyJPT8TDIL07w4tdCEgQEfwXwAQwdgVjg6L2zp+vbjPqR0TgfNweEBDDZettdYsfxVrOA3piN
a8LE386VJsB9QxnIysK3eM5jWozmPklyDkMRv4AFsmBqjjU1CotEBvAZRPVzxnmio21VzcpsfnEM
Pf5HU0TrQjxc44Du+M0iDKVDWAMxY8ctLqAN8UvRcSsTo9VTBs3nL75B1HS0LfhtddY0w+RECi+e
PqIwcVhyLQAB7v7OvGVwhx30bs1coy/KsqG8ls2e685+ipqVD8zbsRXYb3prIX2hINv6vNwCxK8N
7SMVInXsXt3h07sGCH6lcjMNmwjwbpulzIaG7RH1WugjH0qnaEW6nF+ezyDeoDX+HzQB3aN1DBGo
BNT8qu4/jVg4iqY41Z6YS7Isl0Oe9ArGAJmVX+QXeS9dIWMhQgBjAO5HuM4PKSW+MXL5tai1DxHa
1/O61rOQ58o+SD4UOzL1t5n9+ka+bHD6ZBFfLxBzLRLJMz5A1sIkQtlwe7iPpVUXTC5jYM2jIBEn
OblT3GsVEJtkPN4WEVhcEz4i41gKlkKfQ8ZouZg2T7hv4dTxlMmzwmKXHL0QINFWi+h2bjdDeJFG
hfi77j6kHprAxHEO+miTw+tk3a7/zKUNejoHxaI+cKt/x0Vk0NNutc5tN3T0+RupphIbRuxWIGb4
l1evEXtJYZh3MFYJt4335zmW9iSSqg5VLPXdqCw31riLv6Gu5K/+uLDrxNbnGHQXssd0UCmtWmu0
yu2dFZgaVewC4sR59yIMMq6jTsUpXhZn+DR5W5XoZLYUXIJDhS3ZbxRx8Sof1sedAHa8uhJ45ME2
A93EhdHHVum3UAM7A/gYS76hbZ6p8vSGGn3KfhghDuJUS/8acPHMZ3nsRibWwO5wrIzEPBtsTwpr
lOdCw3b4KPkj8Jo9X3lIST7NjGokPXj5WXRHWy4MJKP9FyYz7Mp7oYrIITsQfi021LALmSZgmpD7
4Qo8FN55A0qN7loGr/pOvMrrbHBUfqAwI8+4zS3Nw6PX7OeEML9Nk9BxH7qNQjv2I1jNRN/biRj0
vKt1a3MQphyFrhG+C2d3UxXY7jVcgY22A2eM6JoWNMABlNnsx9hrVu2o0dzXxZh9FDXIMwcen8t5
OnR1CUa+4YkFKTv/Uz/5KavrBBrbbIGYqjwreJnOfKFcXtFs4oXOsUVBFH1cwfXRnEAvSEWMW9KF
iclfbqMTurR5G1k7XuI6Z6rNtFmnweJwF4sAigyBi8wHWvtAkc5sSj6QvggfcScUf3Pafp3FL47f
DvE2FMIePH7lWQ8/ThKEMZnHpwrT2rtoKNpQCEd6YcLoYX/UFHd/ahlc/4mAl2m1CKhQ9Y+PBFB2
m4IWQfav7EXq+mTcUjZrjjE+n0hoYmqMFn813XAQvYjisPat4UhGIw0YjNUetnwkVYRnf1N+YD22
DoF/Lj/o7/MWAqBao3SzbwtoSfW/3nDoNdrSWHXqxrj4dvoqH/VcMbXzvyDrcBdxWnNdIw491QV/
r+BXk27+fjIpQ9vB6X425GdYhdL/yy+2LUpbk477RqOQIEfQJwdblz7m8fonG+vrC6pmzhcfiiwk
BjqpgkrNXkgBmvTuD7JrilKFNiP4StPOLwxL7Gg7EU3zGHCiP46xmhrWF1THRogCdPQBwXRHFLn4
9TsY0IbMcZY1TuHxm9JEpxVJRLm9kPUyscvCE4mzt5oa9UUnvlrV480CCnR28ETNsyV8BZspfYm2
VCYtB2I+nOwtna56SDgj4HdQrUWbMVZZp7TH0VBTwHdalVihYrM+hA8yN7kdoJqDZwNCRiEFt0nE
O3B/YLBHDMuYdAyAUAss7WLQ60ePn//MN4SCWQ9Oco93AtmxwmW2chqoRcKN82ChPILSKL27kDZB
7H4rN4QEKAM1DDNiWYJ6t/t8iqcr8x+8fhxCEc/5HpBgIu5eAfACsWHPFevUfrOupvI2ydVZHHmR
AgdnwdPNJJH+TRu2Ia0ospErMQ/Ra0GMDQt/YMbirfT1W5p9YXK2077+UXUP7Ay99J5YYk6GZcB+
n2KdlxQTF8gRowI+R1F/6PCCTAzT5Gg83pEqTqz8qhnJeUoAHDH0sYxgs/UfAd7yXynwcMpNRVCe
zalCU9qgjmTsQCf1esInwuFB9lm8NfafPq4HxWVQSRWZW/+1ljuu7iyg3BjVOIFjO9IP7r1j4ESX
pZlGqWbFVQ0jYleJeeUkszJGBRy2QhzzzqvkEPw3GavQ4VjPyY+JTN1dfwi2sQ6SIs5vGiBtV1k4
Xie8WUW6u2yV2oWE5X8ajA10zbMZoRGJZpO9Ol21yHDA7O0RhmSvshMXR7ikTERflHPz+TTC1/Pe
Qmjcweco2xuN8FKpIcavycoiNI6cmQtGsbwRlyFsw6QdQQBEZ4whk50cXDewhaEm0KWNm3Chv/Y/
T0Q7QoXNz+eZDdfcqq4GhzRJMMSnx8cBUQi6f4cY/P0pSrMhJB/jOxSWoSaogBP4TYTsGUQVbv24
iLy5OiZCLrUCOzDH86B5o77VdNOnTwgpRUMuqbbgelAWzjfwldtoCF3eh/p5eKRleAT1jFxM6OHK
IpllbPfBLIxBEDrdDGxXZDMTsu9azm9PWhbZM5Xyib32ao1ur1TUvtCiuZZcO6j95P1O/CKMGNyW
G5J39dfgKFPLwcgXHW0Nug0b0ddRv/Cxp18z2faP9S9sfLvR+SxjcWnGYjOtyeWGwIl6sbeHR4pq
+4Rx2IF9a1g7uELWnBwH0xeW8tVlYVqvMDuiyTPvfJ+aHDIHQY9bWG5kOdQWXipEx0DYNYrA3tr2
bQks8xlW4Js0K9aiwalJmG5maBwimRYE31pRW7P8FHYT9jo+ShYoxO57xSjx9ZOPlw8nyj970Gn8
Htp9G0z3LptPiRN8FHKpbVX2Zqy5Yypgn5J6Zv3UZ2WA3dST43G48bmAMreaJObjMuxoIjOL7el/
YlTrAIhTPJqLBYoLWAaPcq72gE0wBrxOxgN8UM+vxY5c6wLp/NyRZ8DtJrgjrXj4/cy9evJBa8Cy
F2xVV6es1g1KcTZvrEUgIHOyI1By88loENRpKMmyfe/MvcmGY6TqKVnNJwWAt2JAeetGFXVyF8p+
anlBv0JIquCjpQx++WqvKb2SMDBx6zbzH1D+5sQibcri6WX9YrsidJFn33Slw3w5it8NqrGr5NZI
z4tW796zSckidK2JKDMzz2DIL4aA2+gSEenoZH1W+s4KU90cchwAUePzSouzXAwt9Wxig8xgIbBe
droRP3RwloTlgZp9WVYT3y3ZCHjXCAiyhYob+qqoBpo5cWLcOJYrGlm2YZQAT4V2Cfhqyy5UQh7H
oHtyCrLx1Iv8K+vPlyd3KmzWm4Qx79BX6ujtiZ8/LnIhun+6/EKkFG8PLER8KYwZCVfpYAkL/Qrx
Hknz47/YTFt5YoHAtQ/kMm01r5ctpjGpP+LRL0AMT0D1KaxoxlyUeI49512k9ayf+5REeptkdnQm
qxRw6yFTBN6QUhRI51qF+IAnvZo3S6Ajri6DTPDMLGZhQ5511yMLNDBBpym1Y5pghXdYuCtm+BXt
oMmzfDssEn/HN7dUJm30jXtw3+BoBGuB/4vGByLuOYqi+fTU72YJdMbuYCltA7K80n9fr+S909lm
piGuzuYpYBDvhQiT/Yox6JmL7TwCSfY8CBQAGNuUe0UZw5Rnh88rEosFdNBFd8HoK7Sj4qDtUEaS
AcOjaDUqzyV/iPZmSbAF2VDrHZFwtEhy4HOOkskXzfRdcs7+Q3HC7uBLKHGG7DPqcl3fOy4Qhw+2
PmYuI9R2xvQI0dzuivVLKzxfizagQK0TvtYZtLMsyCGIKyiTjRmbCfX8v8qAGiuh44HnS9p8acDI
3onH5CEtytnDrWoIK8vhZ5UHQ7Xk5qJvHaqMCMvxHC4jYPcRjojlnohHppYKlEav89i8sS0yU2/O
/Vg1CyymxRFgu13e/RV3JPLQXGfXCjtzBsCvYAEFAJKmpiKDfVunIWfmw89aoy7CON3be06xXHPs
VAv3G01wdYibH4CqbPUDJk73eluelVqolJabM3qh3RIgMVBcU6iI3OdxvDBaiLoOShR7bdwztdyo
xKApaM2abjVgEv4pnxotPWu4MjkTqUqYuq9Ult+v8FjYSbCXWkDQ485JQ5VvhreMiltnvd8LHJIK
5BcwVX9dz+Ng6PERtg+C+8SOOgQB373uuntllJvlHAwP0KQH/VyNwMufVlGisEEeGsYJKjNyWWe5
yc1l1YRA5NtO6VFaEw2oO+9p5IPtDEOvRR3C5m8s8RECi2vaya/qTmeumDc2lazSO2hmGCQJX82S
KX5li2++mVeezrj4VQTj9QXQ3v1RSsnj93ElsC5157OPLRDTP24GyFHXWliNFo04wrMv3JFf1RFX
je8dhzRCVV3nf5ClJxinsQsZybKzWF8gWqmKAIyv7wrLLfjpZJ6UqDfgzdPII2+1CJjO0qW5StYV
lJ9tgP3aQfRpMdGQfQYrbWpBE2MXw+uUPAeDi5PcegiQkGqhaofz+n3fbCBt3AcJihEy6AWvyWhx
VGi9F5sMbA6QhN9ukMl1Il6VGGYiki/ITAtWW9xrT12FrhtiAW3Ernm+qb9TICKF9AEVwwxldfOf
7UwcqvXcP+BpaoKCCE1vvylbI4lIIvqKmuLVLUNrLM0OJ0+VnLElD72wnPuLSglWgPOMqfjfM1S9
jAkIpVRGJ63+HzTkePKplqh9Tx7VdPo73XAEQjZE9D2spu0XlvTp7EEHCWJYAesPHwAP+1d2ToFg
fx7AUm1PSx31DR9K1ZSgzprLMDwCz0CToViGYhheEEEKWX3oWzBVfzzU8ZK/zbdyqjNGriwo6yV8
o/Ecyu7OzcI/jnG0CfzqEuVhg6DRGNQ3snRyuxxF6dtpCZt35OBoDaRgrq1dEwEcVVItojWXr4Yl
8L5LCkWGS6tj7tkwxZ10VIT6HAORXwO7nTsdQX9JOERQFomgbZRxUgaXDzM240OUkduNYaM54mI7
uS94iyyqYkP9UTZbYlvkngkCa42Dc5w3on0k4iKicwxhwgBPk+2tJNwGtMNIHm/d+/RDiW4Z8FjH
J+Q4lEMfWyldbHNIq5lfrd+tkVNIgRg/duAsmICSv0CKw+5zfYgxNuw/ppWDg5geHoykKU82oWjS
8/8isud1yrsy8CZHluadKv9WcWKD7vnbcSDNM0XKS9BLTUemwFzgV8FM27ds9T5v0pZ/QYvay6Z2
pFxm7IY5WPwBIbqqRJjqP5QjZBeEZ1HthO9R7LBMVdDuHnGXrJ8g7Vq0FL992AJg916GxU3H0XYQ
BX9PMY8B/07TaZiEVz5m57rEvSlZMgsnVhZWB6roxQb7L8gxYcebzFr/125T/pxoB/4V2haxo1RX
JX16bbh41r3fAxOF+xo+BoI/eaSGFSrznFZz6UomtxnDg2E9muAcvkNH4U+R+xVCcGul0S6ZQCre
WXfTc65pfwCsij7gs8zkgHlcVSh4/CB2qFZ6lX4ROjOaobOkVJ2taO1ANs2F6X6Ztijbsd5/sDJz
r+qxKHL1VgBVWn9xuTCpcUQ1MYuT0+MqeV4/ay26Tbmq+rah8inS39uAGbHEUG2slXuJY0RxYodT
x3a9TZ38WbP5XwG0OBf0+uBv+5hmx1rgr7Dp1kBEqnre9dOKxk4gOZY2CHd1OJ8go6dS9MBZMSIb
T8dmfx4NtKWMRRjkOj8PkDc14xC1dohJZ4SfvJQwrbsafw6QwWP8K8rqvoiS8mRaF0JSktWV+FKR
Nn2+CPeC9rC3w1HRhaZZgVGocZ7WFAy6sDNK8YO4Om8B0MKruqA0Qv7nUIjtgDvxwo+IAsc/ROt3
s4E9pSyJ4KpRHAU5Nwb9q7a7wdoXYodQYbK3UVFdyOJKSUNTKJrXhwVBC/N/0jBXkE670D4D3xuD
T4YxZpLdjLwUbK0jSn2NHYadTczQTY2+UCd5vB2/6zKza33pbjBuidzEnJIPB5O8ICAhKNxH3nWx
Ygme9ecLzrvKh5cCDgxEgI63UEkzP9o65gjxjc0I7sYTBl5TAdVsO9tkcR3UufgHniC1MJDfh1+R
VhyWhVKI3LQVHbkDsC8EUxQ2GjDvrfldTf8rpnykFUkC1bhuVoGA2lq5VAhnKL9f+wg9VT4B+6OB
x25pJkARBuGPDGNTCs4MtpPICnJ3Z4U8f+XNtJ/cWGwvpodUs5PgBzuIRxCPAbWmF+dRxqYN4nzy
ZhanaG0DLMBUz8COPa5gomjA66l/20r7S0DxwralUc1XjiC4RVe8sd6jHiVa4gddL7L2P4DJhNqs
wNYYMABFMpIKnRTsrg5aWvnzuCCs13KSW7gHUhqM5mrTgE7ldKjkQwBdfWvX7Zy3X89JA1STWAL6
1UZJPMRfXBcz7PkGD9q4NV9TH1CvOt0Bmn/BQTLJPMzmUfUH2dyJWqIoIBvEwTQWHvCIANqtu/hM
zamw8rdTs7yVQyVRHbHUA/odutuS3koqSHpJciO05USinGFzHVZojuuSDEmDStZ2JvTr6DYRGA4n
PIIdxVCGIuBmTDpKGpaTp1UyR0epAlmzo058ta6fT5KEIcL7JaUPmHncp8laLY8+6QKfQbRbvo4m
PEO36T0+ckNo3W7nh0LLMxL3/gmvz727eW4fFfJTJenB5oRtkk/HwNFHVlX++dloJ2VyLvZQ3TVx
TrX8XbUzRuP7hqYOunIGJHOl2drXU/o9EOK0/aPvBZlGEBTBXl3A83ic2Rjfk7lzmGxKjnnMoUK0
r1bi8OLnJ8EhmMKlTHC64JCHwApUwU9gI1dckmwc1O8YFXHWGakXqGopCr2gvQYSxjXGmpgoKAev
d1vrKGbL6MXZ8tqEqGFDGpjV7otKzMleMzPg4jP2rICU25Nq8lKXvtu/r6e8NSXM2WISoNNHqYXW
MUQkiFUvHsiBANZjvgn/Lrd8NrmMfUDZDgPppxGB2HKYpehkl8bcgMJnsPxj9rSk++Fxq5wjSwGj
lGNo3xOuJby7Yvi6D31/kmTDSSTH0rpyqKQnXcW2Mfod+l+qvUuFbhJ8IMjCk7R64yMsEeg0DNG8
JnOsuKOUdRFkL/xkMF9M3RVE/E8EZDBwJfnLDzePFvwRQtAnFLaXOSlU8eAEXaQFBCX1LelEa6GI
DltC7O458wjRqjyKngU6x43rGSq6iD6+nO9SpwdTmIRsETJUVKz6NmaKEhXM/Zx9HTix3FbG3FWu
RTCR/Pru7hhht8SOZS86GHW6CwZsUugpBD6E4fyaQpuboGEFOhFjy5ssHk8se8YhJTtILXP4b87t
TIvWOKPzTb9omz40AhhmuRjqZBTunr+bSe6rVlRSKV0hq5Wz/9BMrkfMDZv629KVHs+9LxFrRkw1
FvbavbrTfN3vK6ajaaW8v/nskF14iglq6eYC7LRzn2aGQQeJifSaEMmmxN/rRHksxug8+Ki6G1ma
94+/q5V8sSeGp5wh2qRmr19K5vNAhoCgBrW6HmHCUTND6Fr8asybY4Mu2XWyg1ZoQFl5vs7v4U8c
LH4/vSHVhSWlWWuFATopDggY14JeG6Q/cRuO0KaJSHcdtFAuBmL5/dRW12ljMyqVpqNjRWkrdI9b
yXGWQDMeXQMfcTZT5jl9j/GOq0fqtrFkvzG8+P4t2RftbXdvBUOtBI8aA14xswQ+AeOE6UPSkLVO
z409hQ7MZicfM8fscs6eLyy7jUvDx2Omn2VCooruStoFgIg/Kd7zZfXE2YsmGNPloO/GqoArGFFL
Cb9sB++h5ZHbS6oLbPu0qtukk79JQ70FVzfLDb3Oq9wxutClBJzcvyH6ki9TL7XPzLwDkeEkgv6j
EbUpDocC3+BH6bls/OpflwJjNar8bCBSC4bGtB1ETz5OwglCnLUZgI0GD9WDGAIvyj7pwKUiQz4k
xI06DQvBKNuAljuy4V4pXxNnunkC40YPXNVJnBA6YOufbKeB5Lo1Nlco1IExLnQsuU2/m6ajR298
Qh9UjEVNytEEB2Zr+aiIFN2cNmcclfwf2yBSzusB1nmXknvq9fBiUMj5xUKWb5EaVLSxK+mMki6c
WXDycK/0QSG74HKOn3XTzkK90+PXOtF1AF1QcW6BJ+CFsP1xZAFAmvJByroKbPFJQpZEpUMKX9Xm
0OtQaFi3zdDYhOvDuNPx8YkVIQdRiKLDqCsotJaO4adyFjKr/W4b6n6Cl2A1M+ugqGhC320N3lsK
wS9PQeDhoHyi2BbaYPDpO7O0N9rwdKNFVjorL8PAEC9DE94vQLNWX2A9OpfIg2MYY1gzW6xxj8du
iXQmTvOEhU/BnGjKIlH4yne+wg69R4wTPvQtjuFxMl58EAj9rk6m+JsorEwO9qw0SEwXUI6JyubB
GBNA1LihXDqSkWK2fMxLDl/lu1oZIgUbqCL1/zcj5mTnW7334pme4AlHjUkvUgbG4lDNBFTxE5va
Qo3b4VXYeXjFE5Jmac8d97OoWFI/evzruiloGkzgIT3yWhtoDPIet1e1bITntFFWLnpCFFpTuQem
/Fh7WkqdwMBO2LnFzPmQMTqeLefkENlMfcROacdZ3Q2i6WXepdBsFRgX2kcYp8iSsM19/12A+Cnr
g9MIu8h0C1UAKNPK9kvqrq7TAoaRvpHecrjNzqsXFnGzmYcW4b/kWGdPJHbVDzKdO9/c6OWrnBGg
Qp114gTD4FrPgtKCFora4Gw94b0zfJVOx0LJOZ98LAOXmhq/fXTYQGh0f1YTgx5U8d9kR6kolLQU
WDG4GVp9zISb0+oPzhOJdxjIrWGGsuebBTSYGPTd+3D3lT27o3LN6yCQFPgSCYnm9skxnU1cv5ZI
PD+v+MQkMfm3ZFHEyza+ONF7iKUsHrXkWOrWU7JGX8jcrBNyuo/OElal8xsvrE55uOvPbspM4G9G
OV32vEfjcjLg7ocFwgnc5+kgFCIGOmOtxK6wY4P2iOYqMjjCyw6bvk7xwKgMEOyloG2ivlTB6jSK
sUrDlST/FH8auKcLghc3Yhpf2pXGbcdO41YNmjCI7vd6I6H2ehESD892FUkigjRKiXdrGXg7xus7
UL77Bt++bKPj32tnaiLx0HotqHO3rp82G06t60jqkSL34aHRQVmQ+SeCco7+jZl0gGxC8zpyTHT3
oGqAkAypNgoVa9L+oITLSvJfE5PH8nTbygDPHcplYmcUxDqOb9yBhXEyqU5KPKN4LDqVtDvq1u/x
ujkc6iep5hBaILjUGW4SORP0whHzIcHQwx+yx9K/zbSrvurnsQd5Gdu8/F4ovtnXyQRSpS0tfJ+A
/bLgQeUR7HnkcXhafFDf1t+4+uzdAF8TcxnPXMHH2vsiEGgBEGsVVuzMgpsFTxVwBv3JO5mtT0zU
B/vr5BcZCgSNrQXpw3Q8qSD6O1LKJwdWscbgj25Rpeb0IMIwNB+7exnZAHm0PWrwtX9wyfuIq13U
+YDiRhu2xe2SFPDfsMUcGANTI/F+m+glcQzcU06ReqhM6vAJc+8EobFITKSNQ0IIT4uQYPZ1NYMS
U1TLnq15Mp/vAUU5ugnfeuWSDWJnTvjiJoLpzmC8gu1GRjgtDgCUKhsSTtPatosV3mAmmO8Wp1N9
6RSBTHwCWtUh6ee3mDZltJ9z7jC9BywP384FO94C1F4csZ8O3MjzkZikDbqNtk0/2mlQwCj4kDz3
vfLpEFG9SMhkwLECuykn+cv/NBU+tHWKoQPT9h9lvXhaQmsGKx6WOwbRtpzTfdjT5gahiN5+i32u
n4YPuQ283tLYyZW2/n8DOLjFueUuKJAt7s05UJ3nWowKB73SMg3N79OoIvqklWKNH7SI8ReHKWBI
RgN/ZqVUTHKXg9ZS4lHmcy3nWLDg4rFsne+vFm7km9PMgBMcxqFfWBv9q6UZIXwevNzeHyqasUzG
w8S3+C+piuEPozKwYEzgZT++GNkRVVWZw54PBgDr+RvpGor+4j8yVn7GcJKYIwCATgMBgLsFVL7I
/NRCy5l2HWJcnX2RRT+ZL6T3SsTsILmoWynh26txKvBJKYoG080pALb3IaoN4bV67TFRwjyniOkX
vBTiBcq+VBl0cW1fv77LAImhUPhLW6bG9RMiMxPLli2wPpynK2GLCyE7UZi+oQl4oxFQesMBwsY1
MiamZEfdG0v51uVKgluuE6Z2dAu15Ax32wDQ/YXlG8oD8tgFNE8a/vWb42ugWlVvU0kPnI2oAXoX
EsQREfBlCAy5WocL+TuljSNviNpxmTJL/ZNm1yxVakgyQEFRVHduH4RoEGZyprqwwMfWPSqqWWw+
vS1tTC2zKh915EKKmVoEeg3Sm88/TsCPchVeTzXxyFHu/hMnYp9Xkv29KVDDqnjpSRY6LoDDlP17
pa/eNgRwFMGGsWtcLmyahVWIO5OYJY/T0fxvq20IHrkoXosK5pZjX0zyZKrf2AIoYCKQztmdvVCY
tWpYSg2LoUPM02jH+Ad5l/vB6SS5Zd9uN2V2SxRqMQO5CP1nbkgn6pcej01y3Sho+yLX736imfoN
gV5DJsoG3+oh1+dzvJ0nvGoxqGvGEO66CsBsbAgaJWWRgPL5VUzboWLa2DIM726MoVzdDyQkuq+c
hyb9rn2XqjUY2lrS6Do4dFeyrXgPUbGzOyOWCetfZdB80kF+HIW1Vi+e2lN63dX/1kygOWqgRY21
mOS97x/N+nbPagZoWvJv5LxAojAGlaTmS13IcRmPMTCp7181nhLNpqJUdVdtf+URT3KtvjdYLyjE
5OiJElwTbfXIUy4XoP5YfNKb/kSIOuH8WTuhJJ4CM8G5xHS1TmcTEp6wCfXG1/U7JqEd8Gfg9F6v
XmkoM9M/pD77TfqjEoh/8hfpIROhIoyn/XFDC7aMzV818rKZ9EPD5yM+rQ3YS2QeyK+hDmLiZ2UJ
pN6d0IsElTLE+GULQMGm+/tm61f1rsi587MGtOkQEGPVlErLXW9rnn+qHwLnlxEd4T6UyUSQp3js
2wpzLntcUtREYF/LHmkbmImJ965v8tc5RpQV+xr0dCYTBaZqL92ttGi/5+HNXRxEE+3aWh0aAxSE
MTZGqejJQL+LENboNAR2SaTQsKG5mXiqGZ9KP7U/PGayrFmUQUKAf4MMoXtKBdybM1HPUOD+uROo
Whw/IjxvcW8YgkT6wk9ndWcdcBfAXPOek9kTH2Irur1YXXGZE2BlAGKDnRFXAFJE04x3b1xmOMIT
tfLN8srOoimx5Wa7i/WzoUEJgYMkr02RH6I/6iKXlyDBhlEpzMPDQpcplo/ZHZ85eVTv15rFkemm
Ld0ZxS7wJ0IXqM/7MaHx6RaRGRI7H3mXg07UgRwIPkOrMkMIoB265G9NSFm0d/ii1vzQ+zQheYdx
lUwKpii6nshVyXGog+8hOl0NK+uLTH1FW0MOXv/csm7fZK+5wpUAwYL5fYhsEtj3+AiVL8TsCfaA
Ad3QlpmsbsywBUR1LkgOquDjbH2b3oABwWFN7zn5WYvqzffg9JcnfJ1Q5Wv187rOyyMeP09zhNee
ds+6O1QS44iKwUm1khPIC74osg+J3BUNDt+uc0cJ7AY0sjT1ozCmSp1js7d3xC8o3YsuJJ2NAo51
8c5tsu3QnXYtJa+f9XXLMxlcqq65zBk37VST5m3fFLZoW+TTekKAgwO3JZolQJqWX4FatLwLSzG8
sXiFNGv6edlvu7sTbUFWyn3ajDUQVjb+ufm6LSDj+B1HVFlX/JIKJhrhIjvy+8XeM83SaelIc+EJ
7cUE529bYno1/Y5TXn68UKfAOw+lkDsZQPr2f3DYjf+SA7HsLNAuxdFQHqJoiXEpPknlfZGgw7ob
VTr3EI5fHkHy+kfC+4wtFrOzLot9X9qCOtEJz1bxUHs6RSA6WRCJreAFlyJeHSQWDIKJgqWkADIh
nHwiDt/O8asbvSaBdnyACZQpVsmgCla1CkunhHEwyH5wTItjZHY3AbmWneZ3BbZdgfvkexuHJUxq
Ya5RFSlmb0ZqruD4s5iti6Ctwv5oZxfQj9G6RVJhJpkiQzkqU1Nhk2n/7l4JncIQh2r2EIs4yUxW
zFxmgy1hmXLypuNyGqg/528O5N6mvREDNdYtvoLssDK/V2a241/zZlpjJgIDzrg9lvPqCH9xx2kc
e0VhDuYoLpdy6fssYxHv5iKs2xRyT/ztTAfgf/mdl7sEZcSG34iXJx57fpy5zOMUwtsveecfctXR
GekbAj3YrxLp4Buet43IAOTHriKvR6HRlen8UfE5RP0ElQ+4K1AH1eewsD/Dgz1tItVInJxFswbt
gDJ80OioSKIF+fBSb1YK1cReP02OZ/XoGXL2u3eFn3cBDi0RoYDt8tfin7lRyXPSVmjIOYk2OAo9
V0C4G4agxaih/4L4ULVg3ldSahIo9+yw+34vG0v6qMFwr7Q28iP8XZOOrN6Jg2LQyGQ9VhdM6M4j
UTvvmK3csTZXgtkg7XwpqwfUp7g5ppJHicKkuhth8BiZVRjj+5tNATCqbVg8jpo8vAHEo/CGU1jQ
lxvp+JK+jleqDcMjF/qR96rcySi4Yu27+VUhpHk1k6FdOmxcnoMalMJQvU6zEGyhNZ0CwFIKTNs7
tt2UXZpx1bq6Z5NlNMumZlf8eNbRxFw4K9wBUnMvcvZwDV8bVHxfc3C3wkM3EDDxKTTG61enwKaz
FEMxHo0u4VREl7Kwrd4C7YCP22rJAax4WGQQA70MuAUvnt8SWwaVH0S13yrw7+806vscx/hv7KhJ
kOwNgKMq/+5t5aFQ6n/7v/iA6Vq3540becby1LYco934wDohTcUEfkuBQE/DpPohd2CJFklaVtgi
3Xpv7Bm/sxoEChzz3UPi0cTFhyXrs0w/Y2ksI03HKTe301ZkSL7F9dt6Tj4d0F1z7fsy09rEhrm0
zKYiNGwTgkSvr1Dqf8c1UOeeOidV+0UdIXEMeFdD1nnpH7Bxm2vt10Im/GnCcQSaqhiWHJm+uNqe
gRNf3lJ3nAwr7G8aOOM5SFgaJrqaYuB+NKJwUXg3blq7yv6en7vBo1FkxzZa3M//GVOhJvTz14SP
GQ4IY1D2xFmpiKZQjJNRrSVEBWQMfacq6Ahibryw4FXryp5w/3CAmfPmiV96oY1xCRqRnIB7LBDN
8J27PA+IuwZoJXT4FaSZQGGn7JEa72SLVAK5zd+DnIUHSGvRn/br4US9JuRdk2ppIHZtjvJ4lxHw
JyUsgebDsKXSkShS2d1KAtEu3dSbkWqekdfXusKIXzML/b1MqujtPtjmLSpdx6KsEMI+cYybjYm2
v8aBfbQk8gqaLiZGlJPIUgh+KJ1JNkHo4RwQHPaI4T1xfyLMjJWt28V9tNWlHCRyh2joAV2E9E7W
XgfgdCDwU90PgfBuYzJXiJNCvDXOlYLk2ZQ/7dTlthxqFB7Q0WxRfE4bmSZBtFKZqGTnDcWK1V6k
S/5Ks5qH1n6Lw3U9dA+4o5VTCHZ+T9MNYHCkJp4niXzvp2X0sp9jIXeC2MkETmaVdP0JbCB43mHH
w+PpX7spJnOIAm8jl5z5mWzr5aGFGF6n4o9mii8GMzeR4ewmlyCEZsogG91RXTGJLVD1XiCXFDMk
u+nZhYffKizehS3MlQUdbUwUsSV6V9x+eOo8a4l6r1qugmHNMvjFf/VIdoKZHs+Mq+8hV/Aw73ip
6M+IzH3ZC5V0U7rH1Kpru/RET1xc4C5xQ1w8KUZrH6sQDZnhUjcDuN9lOU1I7sHUfJpjfga3pNVD
0I0uL7/iheBG+zonlnCzC8LU/CGLZVVRW70krCfGMo+Hen8CbJyP7G6UVnv77Xluugyy/TwPbzs7
4khhYyxA9UtNsHX5E1fG/HGxNhZu48LjeDa72JpCaKMycKnmKiq2cfG3ZSmsEJsN3Z5zGGyfrGXW
+31+zBdMdSsSgo5n0WyGImifeWcIKKir/y0qd6yiLMoqKVvhvoc4nLf/ZaNcW8+c4XJIM43dxnpa
jju0BpmPe40oSGFSPbFFTWjjRlqXOZtwBOfuaJLJW0FuHaEVhOXwFCizHpUFBG7thM8gUfjYL1db
9JW88OpMD3dh0LK6GPxp8X1sy1hKYyRaz1ekGK9jCFvd3OLEF78/bvjmUTHWMZIJs3esBFQ6vcGp
T4YO87QQbenbOof9n9akxwYasS8mTbIyS190rFI1Oyt24ILmYtHDcy0ACtnezVk/XI+GqSZnhTi2
ZRhZNh8N9IRswh4j7lOUfMVHjjvLZgLfeW3zNumlGdAm/dEP26MUlrwDly2nWO6L5hd8RRPtsooP
tPEm+/Np0BZ7CH37yMa3nBI30kWsguvmzI9hqIEOo+qEpf10lxATlDM7F8SBr+hzExzETaoRWA0T
DOcb01oJILfCgjePrbE0CGiA1IMBgGePIJojVBQ2zl3dmqsHg956tXyyOpfbaW5NuUO4v20PM8Zk
LZbF8nJc+YSTIXlpRvyow3kITKYot1W3D6k864VtN//9u9gjPpu93qjAxX0J82qpW7D20psBYnyC
uKwvxlmyrRrtIDClFYL3tEoAX1iKjUm3w+XlyC9dLMpUgebvg2VhNKLQvVHvIORJSuPISIE6b59G
pT5nEtNJ+LFsESJlMoga8vDCDOhq51vfzokeehAseG0bcvDW/uXGcg6Lf90XgHqcm/XqKU0tezja
M+KX1vGcQUdzXmrO3FNB5U56AdSMhwG78eyUR2VJ1yT1hGBdF5giAqwHDBljti0e4gBwtLD53APr
ZiMTas8FtK9pm3vgcFntEarhZHAqJJfqZiPC9/DHsny2Wxrlcc649cvWLI22MQ/ybQVxcgAPSEe1
WNQuAhzy6hQ79pJg0k02XoqvMCg0qEw03d3habuoWOnAYbeYhalu+IMfjMncgxhYOuxQPVVNffTT
gfzcZQSGCCH1KoWQIDW9IBa1HtGoMCnX9ST2vLSOeTCn+dYkkOWWfJ78z9SQE2gwzUzrR7kxVclQ
48bvnGTwIqT51TW6e1wB9jhIVzrbjHR5R/RIW/ku3LX7ofU3SyDsUSGbVGBlML7ajlUUu03VsxgF
4qyFaUSbmALxMZucmMBxpTDC3uTXNx4ElToipcB/y+eeFyRzMdgST2Z24p6Y3XeqpGAOcleZf6jV
cej6jMYyX8BHDoSdgxFWS5E15GMoO7wIX9iN9sol80C6HjllmjFIrKGQEVfXkwVlkP4cyD2Q0ASp
vAYSZQDI/sH/V7Yq1zTy6N+GOiO2ELbph2nkqSaajwWht2jM6MrzFu5ykJi0IPp7yA3FPklqVp9h
c2+0Fy6WOobP0oobxVLK9QIP1RZVEwZy/ReC8IcD2vHV/oadTX7abNvFqqzVRlqDI2kKJYdcNmek
jtYqAv7+z7+LWSOSrgvgBO7lEfT3mO8/oqKTJiJswZYszUgY3KCVTFMtdQQ8GHmfMTFVk8IlxcMU
IHcSfm8Q7FNo+7Ro+ESKGW0VNNO7iB4SaXr0tz2Lh3egoMx0b8vPx+Cj84BZ+X8Shdc5U6FPPDmJ
h44TVXCsz3Q2oVFn5ezPqDw1WgAifm57l1N83Xf7IclP5aUBWjGvepGBp97Ikte9ghDW9PCYaVvl
gKJb7/ZV7x5G/hAx1gqZrEEbwyadGlVejF4XHzTeoJ8BvUrbSXLln3dxxYiSLsTskLdDIO0zLqsl
stXbMGoI7GB+hTneWEh+2j7qjZU3VrbQOC64BrsNxbQrikjZuSKiLceO4fdfhYXDWDkiRCXfwyZW
Mg77yMnDREnj00Nxw62cqlDrBtH56c37ZuqC0W5xNNk8K7qJOYpLGJnliae6RC3NCdanwqXzxfy+
VA+/XEVAhLAjdVj2Qm8fk/V7qutPw696jSOTpN4rH8KE4Js9FCHJz0tH22YFC/TZV3e4P75SbH3W
hLyqF1zo01aXK3/nsZO7bCnuRsWcZCn/eSKsFk5bV8OpoXWqf41omW1Yz5ns6UC5kgWdW22jzuoj
tNxZLTH1Ay1iwGC1uI5oSMn/VmrH7/7xUQu6X3O1gQBJoNSicfLD/hJ+oszFZ8D7SvfAMGu76eJs
S24jOGpoc93RcUsuLKs2Ea7CBQaukpZpl3uwyCF6pl3Oe2I6QFuKw4P+N6GgdOTDtUnT7iCKMMim
5fYHuraOwfuSsE7N6JOAg8HYpiOKe9O+Z8yG0vyAeRqsF7i0U+vuIUWoRvedib0fSCp4/qNRZqw/
6HFhp0Ewv8/wJjQYXY8pXkCsUe0+MT4hxe7gXuk8f8avKShNvqSwvPdA/x7IaurQCR58eBNoQoRa
ptVlhGJHQAzpalxVYAyyQgjjvQtOUgHrr0DHCchc+gD7+FBk/WRYVfqwT/H0aTncIa7jmUfK4bkH
4a45ZxpKXf4heTL/pTxzRrumxFbn8BzWwM7/12bIXjyHw62pn6UvHjXwVJE/U9lFqL/G/jjsluYz
KrzBevLFyvdrAiyt7pxrQ7jQmbxdDMxmYSDN6ioPjrSPqSfNQmNY2Qkz0yBbhbiM3/JaFrJccYud
7GKgrpPVYT4Nfa6oFR/QA+lIXcuhbo6in3oJoe/DIarxNF5R8ZOuGrvSrgGmWkrXrsuHMpxs+n4k
OE6gkVo56lFX+snswtoa7xmacM0oKs2U65M7wsYcGWR6cqxy6ReWZiO+May4+pgn8TvU4rO9Wqg7
/lJWKBqmkuGSnGnoLvJfrA4jivRWnQjvcJdB0CdBt64i14+i4D56p4GFfCQT/2FtetkYvvhLJQ1Y
4O8KD9Y/5otwI4nmQhSHrKn/ZrFbWWyVc6Z/o5zp1PA0toGD5NUyhbmDDOQOhvfbvtowJ3WDqeeE
V9qGCqP8YnOVqq/GLk1jky21U3JO3Bb1sel2d/7q5kZ12Vy0NXbA4Z+W3ohOrnFZKCUrry0BYg4m
flh/1Oh7wvoDVJ/SpeKjYPFLmb3Of/k8NpXiAbddG4hNRYth2PQcjMlnH4d0SW0zhDBrqmBG4ubp
+mA2THgzq86T6Gp6suWSInFwOPgI9Z7rwpTSM09DAA6Z/YdlzeI7WguxEjMquzz2MdXbwMV0R7zM
w9eBhxfBXgE0oHmbmeq3jqgrelu/tcTdrFai7cFcwbn+RbEFdKUWr43aHwmb2KG9dr9Uu58etvdl
/pkpPt0obKvDSU4Jctd07468mX0Q0M6h+kmqihEXBqM3/2uTiO6uhl9tr9Kl+W7il/6hSgNA9rnI
lNEB0h22o+mgrNXY5hiXVNRTSIX+LAvedp3vXc9IDKpKQQHMmZ6ox+0x4oDXSNMCJuh2eYJfUQwD
cWhCQK5LzHEqkW4aGvClF2dqdknj/BL6CODCJxdEJpiCd25eOlIiCc6RnfDHihES2GvineqsMTmU
qapCGKwDnuxt1atklCZHdm5K9pCFAb8K3qIpgb7h6tkc+ZA1gHEqB/V5l0lI1C57U6yN9tB8hst1
Uzn3l5Dp3Ssc8AxyY1dScJHzzIwsvcDklcx6+hD2zJo0JcMzv7k4YIR1lHbnOGccouTjhcv4vOEZ
R5OV/aLhfaYd5F/wWITvuIfbEuowiayTKDYaCUGm2l2ADeQDPEcZHfXVEz5MBclXVtzw3LvPdrGk
u4WOuWWX+40EJ0JXQ4dX8PYxILjrNvoRBjHmXAuR8kEFiWaZNRT/BT1wRkiPkX22+zsma2lw8YGy
GAxUOVrd8tGATU2iQZ6h4rwEtee3yuOA8HmtPTbO/WhRt7iDJ8dLjkeOY7K+fN9PhoTCh77DzKRA
7ccYBrRimgfuotsyFEh88zF0QrHG1fqWVprbwf2XoucUsX2BhQH2wGUPaYhzQ7gRo3GaXFmyL7kr
mfSvNQ9OolJFWXpmExJZCZuCvX4qoj5yGjCx80v5B35efN4/2SY21QLTLTa8qsSFbml8uuFOx2wg
7dVETYrTBogECdBY5pA4O8pAE2hw4TweI/98AK7Oa6cR/YNoMpfIY/D8bbv05os10ek/KR/UjXDh
ugxI6AYhef5AzPuZB9YaFo1fSLHDSfzZkIJR9kbg36rec6bGL3YNPmixK6yUYFr1sGnSA7KxMGeD
vTLpjILunkbdW+pST5lePlAfjELX4dplOLTwxK/J8KSGEyx5Lv1pcG0kw6NylpAY5v0hJ9gFk9uG
mK47CaLkgWZCrqBt9H1sgjN41unP6pMJiKn0Pblv1z5DKFeGO55rbEPcB6PNzeFz4hd/JGRY6pDw
BhNM5523NvMbUSYUye7nRff0xQm5sxarBznAjxbkSd3wVCMdbf7ADvRcCeF+N8CwEnDFsrbHylI9
Cc/oYzljKhrHUInIE2PSMsaRnVbnZCmK/f4sezKek+rg89R1+SlkJxBPeDhD3O+fx/n042Q67aBr
opf9orrxZ5+gQHB+1kUpnhhhSRpUW2dQeK7H15+E4N5flk2GRrbjXJiAfmtcCHtv1xx9ZgJWpNmV
a9B18vx5n6fjE1CZiIhweB+H6et0AhOW6xgz/Uam0L0NCRew5YG5KIqmEu3EVxoSQUMj2YeWfT+u
GW6CBvNLErj4PyWOq6r6AlU2pVJiPAozRFkz6KMgRrVkeyI1vFEMavmZ0nW+TeiYvoF1b7R5TD91
LsaZvoacjFj78Tfgt3B5zMYjsyrBAF279C+s2DyCicWgeQdGVESd84LWRqWAUip+npkk6cz+nSN8
0IXDTp1lTmjrHqfoF7FMxqa1Hw/yIgDTy0c5lV8yF1YGbpUfRLcTNrtj7nRM56soqKbCUeDPGH7D
hrsy91VDWAQszj2hPMSLFFGxio+k6vzpV+nG2YpT0RlIo3HUi5mGWJSAuGWNN74i8V3UeCWM24+L
zyyvrxXIQvC1W9EtuGDKZ+0aMdvGS3yGd7wCAaSW34Pl+Sog4oWc7RHtesqegeU5SCwwAVGjC+zk
a/E1JOeia0FMB5R/eQWMLxskTzPviR1Lu9P3p6RUP/mUXARYlz4ArlEAn94BOssPNr8NKn2xIqPd
/SqVbiynkewtQHz6jDVuJ0OwcN1BjePG+BMcvS06WoMQ2BK6HO0ZYIQkcFoHkiE188DgRrWOWcHU
Xt15kNidN5SEVCPximPgpIyY/QRQrrx0OnWVT5iyZbME8E8Qfki4oB68dvb83u/ilavkepD4Zlp3
gZSGa65AyPtbQpFzavyiQmGwo//LcYovSlEGmOVk9rRnhP6p9FpjtOonV+3P1K+MTpCcroli783h
/fgP1enBPxtg+MHhoackMAA930W+Lk1neVm6M3NT1JvFQPStocFapZOUAqtkmT/ynVEUSi+Ivpgd
4jlFAOjWTpC5mNgZFdYcYyZ9GwaqUwizqxS75W8aP4yHpZY529Az8ko3SlhcNsMDGnBHEZQQnBqo
ymR3RA2pk03PI+ttU42pfHO7kKo2+cZKTCjse6c9j3bUIxO60y9b3DaYaT7PQ9Hdfg9wc2IjTv0g
BhkB2cxG+L/CfSvQR48BqtXoSdl6M0xMVwfB8XaAKIcRvFDRyk6qVYDahqRd/NYoWxRgl5V2pz/X
xuIDtZfrWuX5NaTSrrStP8IkUI+v+Dn8yawQlfudVyZsb/HNXOCyvgxDDTToOc0yGZQwZN8CwbhE
/8Bwzi1tkPJ3hNUUvm3ChG3DNuMOWaSAEysFegVZ/Qg2JnTq20uQFctE8xGiailb2EJnqkXq6/iD
J0GyMlrsB5oVAw2Xv1Q1r5SH4V0HoQpTykZjG3TbdFVYHpbNeNQJjZGk40juFoF/PzAA9f8vXZ10
Z7ke0StA3AdorFRQZzP00QO3zxJruSq4rXkY3eMzIMtL3LUXUz3UQAn8QDtNcerg1CTScr7E/58t
39aUPl+1rfWcEVdh5n+fg5HdMkwQ1dH1z9g3uWG9QPppU6hla+yAIuCCQer+82sA/3ZmIeUBWYhG
cCNALEPT5M6KMRZeikY4fHoj0FiujnWSc5/H7dIXi9q1Owucv7h4m/41L4WAGjP7HelAksmfFaNV
BliKaLbLDpputKXDXA3IQBpVyvGXu0WxRBFaC0U2LvWLIVBxOlB74grSYXjkilqemGbMDWm2q7CE
UKc2GCaYIiAztiBQnJP78cWaBC/5WiGKMW7GCQZVikkKqKmW5EjjTa4lsdQW2IrkI+S5cQ4RN4p2
NsP12wsgZZDZIrLevvgBcBHchxsa/7hMCIbepwwdzrc+stH1oCYyUGLJ3tEKar0WqMYWKPd3Ax0G
yetM+js6XNtA1LpRkMy1wjxvW99hEhb+3G7gqvgNEIStLKkHm+7NEmPvsNFmudv3Rg1aaV5H2+js
ekdjH/u2wx8gpoeScAuGru4+LduLLnxnQBk5SaZS+S5I9PREY8g3fxO3o7WxhXQPjbR6Q0oj7yY6
CNKawRC0Cff/mLOAnY1HGPjhqqqr6ZSHtytKBT5VxL46J8EdFD7BosLvAu2NJMxQYc+nmUgw+RY4
b2QQ3PJDCRsT+V5ZLZ/US1885tJB8CotEIOEx2Gnc9ZTaVqG8m8UyJ91h76YJQcuy3Dd2KKYjXSo
1+MyHT7drgx/41yhhc3bQFa8U2QJHgFhLQ9nKIYhP6bXVrPOluhscLkhOrvKQPcZng2wIl/ZSVLz
OZ5AY3IqIy7siNUV2O0/0ZwWGwarI9XWnuNdY0YdtuQlxBRvFot+fk/gmTIk/holvxyarJBzxSM7
fAwMbH+tEFTI24SiyaXWZKaoQ4mUA6kHyxBkz2rEup4XPrW/8P+ltLjGFRFmd8gwFEXORlCXWN0R
4qb+7y+OlmHmXgA4bFywfLBgvs4t2bWT9Xuy8u99PS8YgjXlA6FcrkW26GfVtxV7eGzgFZ6rF8My
NXkAxAq/+FiYHz6OcILLX2WBCFiTpsNdZolkWljSJpXUqqW1GBaxQiRvDE4AUbmwbc5ZhsxvGLQU
PVBoRkCQWEw4Q2EGktkW1cjJKqh8lDgJA58sMSVNcf1J+dhFRCOvBNfr7ZMvQmAyX0n9AgKl5RUQ
dRuk2o8KF8R3ZMOTbIHJvb3vVEeTO8sWldQrjz1O6pyI7EZ+YpHu+dTw9Tutt0s7x/SfKJ9ryd8v
VyDK1/Sj0lWXCWDLBuffLj2PdYzlruTPEFYi3NbzDrBPgafnh1U+eFMu0SfrNE25aJoHvT2Z0Loe
Yb8lnH+iIApRD1COVjHEhDvbLKYNABMPc9jFONBDu2OYIW1VEUvGc5DKltb7jZYv/UOTe/xUmvL8
33ZZj8Ly3lASUqpDljs/3bt59IT3IjX3TtNryJYGk8Yf6CntP9xnLV9wbbuiHqDIZpqWf06g/sD6
3//PIIdjxWmYNLricB7OKPJy0D9JFfyxVrJzlgZNxUTCuYhss/Mk46RgCFLrVSY+bNmPYrb9DyKs
BtPSQiCBvZ2WjFqbc+7o77U5N/9OZiDlpXY3tDAchhlzK+ZMyfpIEGKDrdT+W1a5dlg+7r2xhlIp
KvWAKrETxjuOhGZhSlHTnw91bgI/aGuh/qm4A9RkFZUrbd+NTAoKEelUGjjPmEbjvOz/m5D4Rg2w
zcOfIQc0Ed32OCSUX5JwajEk76AkOMDNRSqiSwFQQ4tqUFiBz+5bwS+iMiFOkqs6RC8jfuwdAFTf
UuwiMqNao01oFfWjOqI2jf2BGQX2z43wBAC8eZSmGvUe+YikF5C+/n4rtGacdx9biYJBRv8CqnVJ
9QEG0LB+8K+FFxkIKo3CL/w8O0Q3Ji/BD0Sp6MZffbMQxhouesdg+hGytNUBTiba8dfGvflYg0sD
RBa/ZFX6PnM6S+IWEe6mmWS1jJuJr8CNdk43w98wIEma3qF89WSWT6THSofHbdTEsxWAp+g7xVSr
qxfPKLds1cdpl1F3FphT3bn+l1qsUuIZTD/7B2TE0faUn3HajqYWRtUswQOPO1B/QfEMdlDsLcQF
5zwxtEn9OcC/wLxXA3l/sNoxYqea+wy2IvPmVoMUGdhKDV5ueoFCnaLXbLyBMHZ/68Ohrecz/wyc
mNDtlNVH6iB0ZgJ6l1XgUOsFaOiKRFo7bauhiZfcbBPwVxSx8Ro8FH48HYANSHymip2AQqdfdnw6
D4HfHrD4Kq9PcMLgVaghOA9QJuB1YyNYmYBDyzP0HHQiun1fZdYsFKaKFxBhYacM+n7uwIo7HkGD
FI+KAiUp8sdhm4gCXPK+5Lv61/sjtIuYwnAwdk1Sd1W9Oe0oyg3BD5PYRGEjuUMc35NhlST4cgd3
8WAwsqB8Dy7y9g1YLQJQLISa3SmmnjQbyjdwFLKytZtMpK3m9JUH/9Ev83ovqljY2f5aS45ALBOz
nSEQnicidGBQXQdZEtxyyJo99IcONK4AzZ1Pauq0QPUFItdZ0LCZg9tpBBZh5G9mxOazOjcT271V
Pu3ydI/ytyI64uRGtME3PR6YK9JxbXmhhApB5FIRL3Z5rB/oMUNaVuhewJNOUDDCqo7oNZiZJOjQ
CDKEdc14c6nCpdFDzo9NiHK6e2+ccM2pYoPXCG9HMzMvkvysZLBYAMVftqrTGvlZlCWZb3ulF8tU
lA/h7O4GuiKc+7ABNkestdzvZOsK7kyzykQelIZjrkpNuA270XysOzbiLmQ2MSeXTA9Oau3N8IqH
502mgZ7iJqp1peC6M6cYwCf8boIGhsNkxgTSL1halzH8g40AyodSYxKc+tWaVtlylzUF8ys4Cmmy
I7ulNMxKovhCUyJFjfaca+uoi89Azrh+Zu25rpcD7rBZbYAHOWrxIkMoSJXGCORXpbH8yQncLXz1
AjJCgo0gjLe0p61DeqX0UfmU9kqS47bESSM52G24GpvHZ9+kAAEjs+FdLSN9KyjweLD7Bg8R56Xs
H9RFjpZhK1m4mrDN4UGo9iWcHye/AMIEHHsrRM9wMkjzmTF+uv5qmLH4GaXFgJuO4zOuaufMse39
7Q5pFw6DeDLll+GxFmYRcgYQksnjeMl9jKSvwXtZhkXnRRSoV5DTdb5Ubu6m/ZDgKTK0WwVBmT3m
oSo+HWJ3Vpi1nNy1P0eRPqzFRUtgQBqscDm9DT00ryfybQmd/6jAI6QGF0/4b0Nlr6NMgIZZxyzB
SVSL+s64z1rx5Y7DvOI3voyUBhFmlASdOTiPDREfXGNnqgYautb7XaaS9H7CwknxBvr30haGQapS
Dkz4sUYbzOlNVZRF4mY6cPcrCZiu6yOqaFCIJiqfAQAEPzZwNzL6dcLIyTQfWy5gu86Bz4BluJGJ
Yu9dNMJO/8aJu9tybPlXgkzRsx4l+CWYuhFsqA5Sr0ynRb/ZuvYUHnrtkE/rxTt60RFmQY/eHgxa
EOUp/pttA3fekdgLr31KhLGNA/xjPo9uspBuvZtCw4mO1oOE+2LhQewVTBUI4434Pr7BckLFICEU
BWRkchqDWdKqQ+xyYY7wNUdQ3PvSBEsSMtbv43NgvGc3aVLJtS/gTwC6p4tiF/KToJ2NKPKe/BoA
KbsofesAxtH/g0f/1LPRGTkR9Fd7nkbJkZs0ObRdJ7oeCTMY0NapogBt0BVRddn7/LCbEQDuNZXE
x+rf+0nFPUNLG5tvmynAqiXWrL6bJndSxc/dGVIZCdsb23Ov13sMSScretvSBOarbBfIxHCAwRU4
JkfCfaIK+HJ7s7bb20Ijei2I4tCahcEhs4WED0Lkv49vCDXWbPmx9QapW4kqTbyqMi7pspuEhang
kYoevf8BowA7NhCt7tsn58VTWPETBoVVgkfrNwZompTpTVbgqqScIC67EZ+/mfAOlIkDoKUYnQQf
5irxyfJDb/gZalaVezLYv+182VAg7tdH44rr17hK6laGzXr5VU8nXw+oPlJWoo9/035dDWhhhr95
nfNOMv8WUIKrEnWQRr+bKSh87y905qdKeDzkpAhOW6Nud+64yIy2ZWBWiy4yrL+B/XEsOURfinSS
OuMtmxBhPmfTx+OKM0tbKbwEFlzz6bvgC0mMUHo8/+gVVEjLGGjYudsZaI/J1fwXHc6PoT+CFWW1
gFsCUkUe7iqncGFEVUZGBLDpHUHytrogUcvjv6SqtYoC5gcwFbx0nmcqNEnfyPZMhlYOXSr2zg9V
+V6Vdewg8zpBFYIxLuK2gnLVQD4o03VIYtbeAbOxP4XPjdNhHnq+HcWwXud/nsoYjqBTTZmFUM0i
8H8+dIviDe8ed49RXpH4MLbdQt+oAM+7VhKQVU4nKvwmNYxF853G9ArikmEy0O6+fu2ZwCtzkyGo
oRO3pBJ3Ci8EXwc9vQBRzqasPVeg8gB9afGZ2E9oudJJqak8gWT7xpYVOnIbYuOtdFLEnQ1qPxub
TgwUM3n/YyCyjkjOCHCfnnV/BjnHyRxhaleFALY8BclraJIie0cgBjV4HFQXvG4NxpYjcyWT/3KO
uGwHCkixt5U2KfjyFJsaqpMvXObOoLreSLcAYt+++Gbc7Qln9GHcsHtIT3IBJY33vsY/P089HK4r
C4a/3wkJE89KmFpUQ91MegDF6rEzaTt8DhkWc4PDsEqsR6tx6bCZ2e23sjELEKqYvOJRjkKzx7rX
rQexot9sCIRvKc9SMxwuAKgSknZVBB/UHJyzeegq0rGNP3Zj1Sf/ZBSAUvHC235kgGfZ9A4i6Otw
VV8mfAA+HwmbRUEqX2fpIaxSd7kg8rAdhytARv8UeEEodNyjWH1x9SXmUiMyAxYPls+5dSgFLmy8
4BxEqtCjvUFpVBhQshyanRqk/fNPchQ4LgCeOHQ89MDxMVu2Uc7d6KobxRx2cxjnMUdwR+iv/qO5
sDNvp2sHT7RK8SD0RFEkoX342nDm0kRR3jvTtGPyPMecqf3qEIjQ+8weMOwgm4/uoJZMCSZ0cm5Y
mvjDIhbDcAjbMMnu4dsvdkGuUGuclCh4i+hAaLvLIn7VVT2SvmVxzv2GexTT2xXR0f5vOP9Cxm+l
rVMr9NqsbE1X/oc6/P2bFO5ePZxgloiP/ma3JomJ6MYiKRx9AyvaPhPp3TxAHyoRKr8sHHxcX0u6
igKpfXIZr09xOySqdKN3lRKaBc020FQwKjfJpMCF+R4ZX+M2JFTkDZLyWckKJriaa/qteusC3+zs
PpzNqzkGYlWa+1ocSpLSEappOFmCx5lMy+YJy00xLiWEkOVj3nDJNu4flgglQ42pn8EADEBFr1Kl
i0h6+RQOBJ9g98aY39Rqw0NxCFd8hjKZxKBoVAEh4/E8m9Wob9Z5ZXArlgtvLIufgZHlRhMSGWR5
hjO0AoTwVQwNTbP3pPSr8MNMx9npLAEQ3Hx3dF6+XVyhB2O0bhZbNPar7k3J3pdNSjz+tWCEFz5Q
2jF6qCKvIikMgoc9Xh+QFJmuh2MJbSUtxOlwZVY8dMjFoFur2UEdjwY4ZF3wSjvH8FXaEB/KdoQk
RCA9nTgfEv+aNU8DgIfieLu2ojm8xGHTG/cZ3LqesoaYbGT8ZFMlAUyiUGpgHVikl+TsfEDuu1JQ
IG6MVTNGKa2TyGed6YOv9lqXGsyBLXvqsULfbkHPSuWEVVPa3LX76MWjqGpxfQmvpSX+4ixvB3ff
fL5sVJri0m4mkQUa4xdFkUT3gmi2Ur9sT9Sbn2k+t1iU3gL4VBdloAtouzwNtkjtPOaixQImONLw
IYBun+lxs3o3ZQzzDSGARUrmJbqb1eeTEAyXzjtfDmGEJtDvm2gBLe2Wb6Do1gLcLRKMa+ws1xaK
73xMUTYanZKhHrkT3nmBFfQnDIrCHy6hEMofnX1Xc9Y7csUeE2oV3JkEOGFQxdMRtd97nB5BQdCt
pJUaNiI+3sbgq66ZgjmWVNgYOYHDGxwxv7FmHPwI7l5vtWeqCbnoZSOeyNUAuIVscyLm6MLlcgTJ
G1ZyVlSpa30FxseEAweOPOzF7NnMPOY3e3oD0eD6MVf4urpzuNGsa4u9i0os0IDunvn84n7Go0Hp
k5xygfpumJcL+v6trTK4pz5rYQjabsSmWaKwX3hKszGt9uTAvXDrhia8Nn1+J68+2xXua4d8aES6
dqD2/hbr2KJNCXpYfW1Wu0LoxeHmuxt4b+it4pUDZymVEvQt6fUIeCZgDhOlvWV2BegeKemKmlop
0WHtKjMU7DUirpRGNgmhMWuCoGge/nZHFgLw/RugqstPIJaLGflC8ZvgcZRBUo34sP1tcGnvIKPZ
Uz4Ar82khrU+xrv9PDBOIEl045ISxKJlyhPI4mc0lcCPD+bu+xSVShYoM0yzvJqvsl77GiXhoDe0
tUPTFF3TXrka3NoU3dNuccsLhIHMJa+VcOohlTZJfdYbY59u4MPkapu62ujcHJ3Tcxi4zymCs8zZ
j1ZVPkxSI8eRBTCaf7DIZutpKdB/fOKIjOfAxUL1v8H7mrlU1LCu89EhD6EBz1/zQpCAHvn1+Bzp
sR+isu2xJeZLBmP1ljy7lak+fxpOOTUxLqkJ8F/Bvgl/Gp1P85QLPypSg2wIlco0mwSDgAPGTJSx
P9rfg4gA+PloEHmgnxPLfybO9hWXOBODhLwsGeH6+uM/clqAQoK1Ml0pc3arUY84hrNcBA6l494D
Y4/1mHkUw1e6PpIUzNRjmD7nBmhoMmCLeti3hUta93o1Qiq1uwhx6lefS6maIzIA2DccxuzFv1ZW
d+MWxc+XVO0pmRYPCy575d9xi8LphcPpWximYGVqgsySkBT/tX09F96vFRCQaOKy29F632AbbSS+
Fd9KCMcfdKT9MGKO56ksuHzdH88uNM1uWYCFQ9INNqwqxVtvNX3jDp4MwDtkpseIUlUjfgwnmrKf
qjSlGNQM3Ml0nfaCFeJv5CRBttOL3ecvjtOA1vN0KAI85EN2IoMpUF3K4iWeDl5/YFLR2GvV40hF
DiwtFVEYwxSrNwf2mLvNguI7L39dezmofW8AXQ1S/nUHjEcX3BkTlkzElwwGcjj7gKtv2ijCvTcl
/BhbwbJ3/8QqG72WcMeC2q27dj26DNX9ZjnnPed9iOklxWwjsrwI5Z13W2HCTO+bMxhnZeEFPZeu
Re92OmEboMQCNYhJrUX+mb9vR3yI+GM97/f8yzdaZCS6+DZyXh/472HTF+nqrVi2Uy6E2aZdHg2X
BYeBgG9zdm+j4nhx/99NLlv4/3V22S75CNGFftItuVoAyE1k/J3v78bgz49oIHBxXLcqNue+/q5q
K+Rtbx0hLdJc2eE94CU6aNMR5aSCp2LyrOag24bQ0xM0axmZkK3+ddynFvnivM0Tac3skmBayMNO
XcZchjkPZYYet3KPSVrOJ6/rtb35xDDzu9/PZKbmBGxu/BQu8IyoDJrL2+74EdApbc+vVC43kqoB
2g8xx3jNthWdUHw34EC9gNkhstbFyZRSQs0r12ooJMukrd0JFX9zSqUZTbsLiRzid39aN20J3IQl
txFsrks+yt9qYw0SDyqjHsIi+U/ehyzfNxX01MmX/uMAT2nBisB3T4AQkDNOjVYJYef0BU1wW5ib
OXsyinx193PKyOJen0HuKzHiaNcfc7CtBwIi8iJdNhVDqKcaosA1Km2iWZKYcy8mGr0Szo0BCnzq
ONFGIa678pbB0BsMKlSVA12n+jpjk8FVo6/48k53Sfzi58IPCV8Ylg1gaTBwaZ0dzQZPqXBOYrzQ
WVNUyiyr1acFVtpwPKLxD6CvlKcysp0dIaSeE95NFtpAnyCY6G5uCb/HCzw/mG/RplhisldjuIJD
c4JxbiAA1YoPKvlUvd6jK2SX0Br3ZvJEEM+NaX/WHi9vCFnzlx2TACF7qFd+Wo4SwVtpXfSh59Du
HaqbwrohtMHVYjnpyZpZ5hKzQRSzplmxCghgdRit9rZMPNyPSQYztDsYIo2oGqtQRY3g3pemI8te
v3eIXTU8YkRVstKhmdL/KaU5HUBINKRn+JUH/Yxs2BoIfsul3+57iRFeDm5HT7qaJaWVSJ4nElS5
rqtRD0pDzcejnjv2bPUJCGODL97+PjpcT9wvEbhPWxI3sad4r1/lgIgk4F7YTmz9SnyQ6qvVmgyu
sZi0xFI60Xm8PSCV20/EkX8BUFtbkFteNO5FJvw9HBuDq8w6YR/o6VMWGDRNbZKxuMIiSqfLmS5k
bfuKJPSlAKaWKnAK9UOSZW0HWmeFfBswM3hN1Bpi8ANUiOHZMUqyX7+iAEE70VwZGsop81IoQAgG
QsA5uJRz4amaK7bC7RW9rV8ku94gBrykGX9qKWk3lRJ9LQg9xvxCrakg5tVeupySZj5qRDoIFYVu
jfisZLJq88GWBAmqi6ThpbHHMjjouWG8mb11WR1K5+J+WnsefjVE/lzCc1ZtPaUtKB5oKt0wTuD9
uo8ROQ7Dc5zDPX2X7ZcJ95nK/vm3H5yELDitJlBVBh9oxB4OSFVdybBXXPqMiY9+egPiFrvgCDon
S2o5oZdm8jNdkmpCgNwJRtr2YpuuPEICNMgztPOoll4cFD+WtRCqecJQYmEpDnolRpqlnjarwHZL
tFPzdCixKp9KH9ERBO0SDb284d/+FNh5rPPGS2QhZyyskmy17todB9OI/0s//TAojfNkv31pZpUP
dGKFpg24voowKRjnTezxF0r76t0P0/5rDRRSXT+ebtm0LU9lLyqu8k9dJ8Q58Xou/qztxUoZUD0K
iJfuRHYScRpBDDP84/fjbDWsfn/XDVY3NgWyGpEphxiC+jtxr1VZkgF8dpJXTupJf8AMJWPGRSHM
kM9pSenKt6c/PoRtaz5Zb3akmNsNykk7opj8/6GrHb2SACfjGNFHCskm+ISmUE9VnqKDcunHHAqY
rpZ90ZeHZm/ETT7/5Gnfw5vrT1yTJOEOvgPWpDhEKZlMGFi3X8UxQFrwtls8C4U3BnHERy/CTXhe
s3ukvlYt8RPE7FRv96mqCQNogbKicEiUTL139+aLPK8uB+SBUQqOlROQIdnnE8lQeTMxtyseJy53
Z/1OUCciVhxc37K4rbvdqbfk2fuVNWcDeAifOTnl3gf6KEReZ18Ybg4boEQpZUPBvyDbKPEhmqNU
vpHcOEnNaB3TuLPTbxgkTHZzXfhrtnAcJa2qZeejrs4g9fMHjyG0zi63J8rRibOEycrwoLEK9JlE
AIe32vWA8AWWVGi+Kesut+45U5qWEduvoYVsRz6ngafA/OZGXGZgkPfzFzoQrlbhtSk1fCYe8PVD
LnCml7h8yWMvE9z9uyZJGgbmRja7WhsfuCrUSJ/KsRwd5rUSRvzrF5K8qWd404+zSf2sPUGjTUMI
vuMkXoAE51myHhT+xVoPWZq+SSYtZAX6GVavPFH5Mhmv0LySI0e+ct3a/bNd0MeJaAX124XiPfVR
uvpgvwDYU9NMESbe8e59ZsKSFwc2sVvzYmKc6qJGkMjEZmFoxfSd6RbV+39R1OoXeLxCfWjjqGC4
0FAbw3O8vjUqh5D5vpsWWiejJhMe0gFQ5L43vXFwij88b2IJ/iviDlktlnmqQMjgYkcTq5sHRCyK
PgOFjL5wsxO4Srj4ToZwNuiJN55EZcDTenO+jFcias2fLotDUNKL1m0mUyaFQvOC7u2ZnIwk+KnJ
d7SFRrFX/9I3mluv/MQBKVjqYzButbnn3LZDjHXaHk7l/8OSd0bz4UdYcrAxRppFBZp1T02o0RZ/
72CX46WfaMOCtYxW0ccNJIVP4xmUOzr42o93i+AslfDhhJ11qRnvo8UAnVqPVRz/TgFGb81cyMqt
nJ8jXKrIS61OcmrY6INOFcQxPmoU5FXrD9HEJlvhBsTEUqcWbDqTvwdVmXQU+5L7bfZ28hlKXNxo
5dZ0RgPtK9mb1qCy+fkCwWwQFphM5iUQgpSexcJCyFijOmp5ZK70EUjVWKMkYgtFYp4NgftFlrOg
Qo3+EvU+l/vCUzLDux3c9w6G/7FDCR4GobblZD69Guqi5QNYuKEtwMvOvx5VM8RgOZ/9UFI6SLcB
XiZ6gSd0rg5TvLAcKOnbpL9KgzypN7NvH4suz6CB1d/Rwi1dnA2aCZEU4bZmZUjJ5kbtnvU1zaS/
zw+BGpIq+P8Au8J93gjiBR6D2IMMiwJ6B87RxZTZFXlix1mdZ3pvmel/CjOh34ZAOUUsi8FgXOzs
iKOTRhkhFTIhpD6hMN954gE+TiDkERvFaYzLw4nK9Ns7usTXIoVZtNiMIex7nuOvQfZwy3kodAZH
QADxxuik62LGQKcHlDSlf6vFSOtWhwvOZZ3kAC0gkvFbtMfSuzdSZFC/620QREJ31bTbcFQtBnLp
iCO5OkYC8/DL1+IpfyNjhVHCYOgR2+lSVPz4/XnKJHLaoYWAJvIfnLBb89qYP4iUVK1a+9/sjyOY
EOjA7Phq2+0RN+3906UYKdkxBmg8Ybm1BXc6Fex+j/DLazAGQDwC1a9+RkQ1mp+DIrukCqj+DMPM
u7zWKTelTNrT42McAvZ9pBurAypHMkoyynkwn/j9WTIoz/keDK//uhwtI5eEH6x+dPocJMxx+e1I
JNcmMiDUV8KYWumRJdPdOVwtsovERPDED6qg00tgu77CNmqHNp8YE0PZHRUgCfVVOvUggzuIkcrL
PO6uQqYDvWmcyMDuIjNjAA6HqAsVvUmT5CHWa4RnjbCmejbQIv+0V6WGrEDPMOhMYsuPx3M/U6QO
o+vV9BckehD3IGIuGlAc3N+GeMhEsA02ER+v/M+wIuzZ0+jtcpz3i/tORBgBsMbSTeY++aSsweYE
QVxkYq8bk6IOZyvUdwvHyzgakGwodJ7ikdEcvrmx2WdmQ98H6I7KzDn/IJm+2MOeGB9/hXETBfSA
u0c4wrdrXgT6u5pb/pUzwD93KNVi2+S+2Q4eLy26ej8dQ3Ww7xaH2TjpUxydJ4ZBzyOboWrmHm+4
dQKqwIcCOUOC+2zC9LXA1ig1uQTH5ArBwGHfWXtXhV+P65WZlj7FvEyBNN3iFRN66g2oXwOLtCu0
QLgUrC/dFFJq/wgNktn2C2per4egcaq7VvJo9gjhpNgTs9yGF2GO6gO8Ib8OyCGkUgVlWYb+SChs
CqGwzVNXlSe49ZYl9z4HsfHHEAN2LbOWMGodK47DcH/PDcUQs9PACHTRMH32NWn0eVIjQZlpn1ri
iv2b9YTGpkaSRajrtQvULpOGUSYJRT8DpVhANz726yKQ1RhCqBa5PHc/4FojzBTEbAsIx8KFmNL8
0iF+XJ9XCHXiU7AkGork4TajFzI8NJdXhJRWgSwbpCqiJ/5pq+Z+rQ+yqjkSP8J4VDpOtRGNzYcx
mpa2dUhnkMtm8vkYEXXaqLGDcGr0TxtE3wLmVh/MKKvhAxlAga7Bap9wfxYahqZQ4nljrnep+KRp
FtmpHTOIn4BPNUAAHNPh4LwQEgzdnCcCUk0Sl4E5q6f06laYW9ioOTss7ZiEtJA6ideoE/1BCszP
bgtDyWLmYQsZjtgZfuWPVnqv9vVgD3gP8B6PuYgdWjiMs/ciNey8UYYqbYV3Js6mrUVnARsmDN6g
1U7nv7nPZYE4zg/lRG9OFDoVE0oVo5+3NhLU2oBqQGbJkzQTYySU7ebZhIAlcwTjY+gMczGWeN8T
a16hN7QwSjA+Tynkua3xBg85c7kM4aIeB51gUk5p3dUKpB+lFHgkpJ6rIm5SW9+S1LbIbvReeTu+
loZX8uQ1QfioSBYgiaG1sLkiJPtSXo1l2yRxqg1ZVsbqj1laFnJLG/DnAUHRGupDhW0XU6uLEOSF
/xY+xHKe/V7wa+3IElBygMaOOeEO7/FmCc6hqif515rdisyfSkVkuBtca1JeNggR4cPdxjDCPnLT
5YBmZqXZ6zWfbYXwsDJoKgGhfnzfjykQIJTjBrBpoEDmwZY9lyB7DT9Exyv8nTzHpO1I4gzwylk/
XW5kdA38l8PoSxZxvBdHG4dtZJr1D4pk7wCnBJS9kEw4xW/nfKG7xR7xUhWb/fgV06W7XKYI39Cz
QP2SpnpNGP1Ecox3sNzsi8fohycbDiS6M+CFNm7p6YHdOVyShPkaEnGTV9HtyK0s1t1GGXCYGww7
Mzn/NRi3s3wmEJOosS5qhRkiafNC0/qM0eZtgDtZMLG21p1exjRctMvnpNKsi5ZgbEy7e4xQYCSG
VuETNsmi6NLGUk11AHtn4xd0YidQC6Tv8p0+Llu7pTRrqE2WBg9ccPSnTwEV3mIP6CXvup4Y1BMq
yOqJUNnGT6bKQ9+l/PUkHoyQbmVixFdyxU3Jvyhxs8xWNmsNXZtxX8TrLIvJdfle6vYjq9jP+DbC
m4rMYJ8Dixg8bpAk2lXcTDbhb9mlyYQGUEgE/oh/9JfPmDoN1+Vy6raXPJAzVLeTg0DEaG4JVwxL
7vNSQ1IiEgJ3ylZ9TvYmyxciJ2VVPC2p8rNBztjyKdOKXMPtQ8KnS9NeaB3FlNryrz3yCTCIA1c4
6x9AeT1CF0ytEcv7AVFZ66fhHYDCr1R3+poiGoaHQ13EAGJl3IJPQ4OYsAtBDeMZcZYvu5Jex/Jn
sOQZldN2spK517eASVZRss1clDHIPq3RkFANdc8ArK2nrHoccm4xZhAV1IoResZ3+h6O05ZVHUut
rxcQIFcs0kFJQrMH8EDW3LQkVH540msgavSddvKY7kWhTU8tB9C+RXis0fVnxceQw2glnoYHmI+r
pAhXBME3QuZZVEGlV3TbJCee1J4TCAF77vMQZEsi95vDC24cewfnwn1+bnYNxk6AdDHbTOXTqg6s
asBJ1b2s75SVdChRd7Uv3t6eg8RbWwvsNm4mnbpG354hhDEHXbJpSMISIeoD9QwmkdjvUJeOA5vd
5GeLmoh9Fz+lbIiOX6h++foLRAJX6hICTgQyhEhgt1P809haxnBd7U5jY9G+z8mUMXd7gX90uUP+
6yuEy4gBo1k2XIevYtpCFgTM3ZyshCq/g4xwwJApDBFuGVGmVuaphSN6aOx5D189ZYQImOw/KbI1
HHBPEeQOBIFKd7kPL8HX3Kv8QSv1oQn6tidnFizZbfoFT2buGZyOqq6hlsBOc4DNu8VOsKn4oP08
+mfW3xczVVrVAD+8Qh4mME0p3a0rw9p4yjTu7yzNpPPSXXS4Qs+ev0QXhlXq9FwAoEqY+6UsbIn1
COdrd073TzYoj8i8+Ec4Kk6Agdeeg20YxTSgK2dkqiDcsLdjwQ1MphGIX/xCdJl8Sg+1BIkJWnvb
R/R1tCzQFyshmWTIrKanDf6z0b/x1jewGLsiKRQ0N27SAV56/7Pzg4jBHJuoBSbmPmMhqs1nh7qK
WDaV8/LlIvdRkTc+Uf89eqT5W5DcbooO8WH6nHp8D9Wim9r5n8q3EguDyqFlpvxOiRaxWrvIwQgI
8+AMXwd6/A1W4OAa4EG2SEXmg24fQ/HNaxaebji08nkxHO0AdGe4EJtcKQw56hj8hAQt//WAQcTf
fDP6YfMRRAfff3ADTab+ICKZw0DM0Y1sbyFCE2/CLkVbkM+CcAQXVI6kaDG2jOBJMYtRKdaxnpd8
k9FL3WBmLQ9v1NI7QDGwHFcHOGc3tCqyW+3h87TVGTVwQaqX6+ZbDJm47B8ib87dAZlYMr4Umni5
w7/g5HlGGjGIhQ+VD/fknIFyUKbkWfcirOCKR74ABS8LelfNrTgqjQNnpWRmF7rK13cdI05fkBaw
U4vBCz+Hb0tDhShLglNtxhrjaruMG0jUVFXKkedlW+owgJqvIuoCPaMPHMLpuSqBpJQCixzYHvsG
XL7XKtUFcTNlN9+nRftcFoIKBs5CCtIT7wET4mg4SbaD6Dm2E1kBmxOqU8Dr/Z0hvyZgvK02Aime
tEiWOmOYv0XoOQ47znD0ZlaSVr4D+68hklgzp3X8amB3tU915y0kx5zTOTXqV6tRWS8NYeUwIE2J
8D+4fnltF+Gi4Q1Ph6+jerlnq10inZESznxR3rhgORhhTE2ZptsF0aNT+HsKH7LykoamMMfe1qMG
1hWHb9Wmv2aH5YS2Pae1p+jks3yVzP7J1UD1Ou/3/eKpeI9FGkukr5ZNf54PeQ8kCgz0Td8+IH8j
d7qGfDHsReGuqfaNow50P5pZGNrmWZwwTDmei6YgY22jfSHKCELPHeImFzCWFSmXEv9mX6y31hY1
vYOyN2G/XYkYut5HSRBUOfYMewM4s+QhsE5uW/2Lf697+jkHKCYEBNSbEYHpBZVvNh5m9apLwruH
Jk0M0o5EfJPmm643HJgEu4mhM6fZEvBc4wszLgd2ZtylhIXZsDEqxWFEJehml3ETJ6rgFo+K9f/Q
btRQai5TeMlojrV7WoZqrK1I3dyrPZtPthAcz/lSkZxmFUNVIiZTgat1AM29UAFLpVwmZzG8LhyS
H2xlyAd7WmaQf8ZWOzd9dXZvzlfoCbugtFAxp0uErQTqwls0oI6SXJvsSjoRO/XW+lYJBtBLsE3N
+oic0HNMc2ctfjHYi57pBBxAmpGvOLTGT+XFJd1y0uw/yMnG5nu4KxquZWyHDKEFFGg2fuNF3JKW
0IOjN5Odj8GJwGde2ghT/2fXn/Djr2t3s3wooYVpMt27GppYbyTqDVKvCGd3eBuvtNB+DCDmiFGN
FK+VuBNP/mTi3wBxOlIoZkVWyBVt7GSL3I9WkH6mcY0fdvuGSTPWWLSeez5TWItlFMUyyqtfs4Ow
0JXK96OrRB9XGnYG1jxwJ3whYqEIMvoWd1ke+OSksC9UoQKxXUT4zuXCn0Vpw2ylIuV8ZXRyU8Qw
dcGjPDSvzwCGfu/GeEhNY86/hyiPWeIj/26WJ1Emvg0JSs7JjuhLe5PqbUzen+HqB6okWLz9nUja
kytBiyqseJYOZkXj1nDf0bJs76S0Bn6g6BW+5xVlwLPgyA+/hcNBy64m4BBq6Q7TbwIn922Y4K4V
TbDCR/WpxJH106UQ5x0G4x1f8KvLumRkbUiNbCA2RSsZEw6EFTZ8ACfmDzYzqr8hrnVBTJ1Qc6N5
pKLrwo6L5eeabQabX4bznHZgT31G/Kvy6mRDxI+JQ8xhphyKt7r9daqnULENmAheGeNkUD8TBMuC
r2LDVoM9xeu3CCJOzt+la1H1gODZnlSp0Sc/gnbsoEauIUjxkPSQDhUDRpIvDoBD5GOUXboEXRze
f4xKOkndBFR3L5WEYV/SoNIF8hHNMsU5lI9fs6v1+VOyxQ9KWlL2GdZfUOp2vKTq0VpSq6t/XJmX
e1gI6I7QinZ5ulvmmdw4k0YbXfnI8uDkhYxPpssMulwWdZgsE50Zg01yLSCLL0lHwIPxLrPCpIg0
U9Hy8XbJY806xN+v2ntgCxlArtT+Gdhjxycvdhsyts1Gnw2Jm9hMn+OC3O/Z+INfDl9qL7B5LPkg
PIV6TVVucUNjUVoSC2nYmXV8vP9nDO/W5FOEpTqTE6uxo1+/ljP4wKsk7J59Vs1LEB5C6u9j+3AC
umrsVI1rYob8CwStTy/bhvF+Ascb3abchR/AIcJaqLFSHBarfErjSq1nh+k+7Sbp6D5j3E5tI9jh
ddyBsunemCwfbI3kXLu0YmOR7GI2ROvPaxuvaJlJiJduD3M7tdclP/d14B20p1c99QzG0lQCnWqO
ihSm9Hf9/Qaxl7C1rMdZgxMbUffOIMf/Iot0kAxENwi+btI+vqUCQgQ6t37NCchb3I9l072zaO2P
r72Vts3e+luI+Xtq9B8jzp9xi2kUkrUaEmgxCS7Qd5DbaEhqyY6GkTb1e1f2c4EilvC3+6fM7frd
fMTWPNaTpMTZcoV/nH0asqdXIpnX9oMmQxyJBUQtAvK2z+WgfHf/JAV6tmrl2mM+/9G/sj3JbcCO
8y7zkb7FjzxElLmCsnomqyJL4D8oFmxab92AArI08pjj535jqy8ErfSvLiW4CuvvXKtjIhlHhIhT
tVYFtUPQXywUMa9TV61ZYWz6X9RqmEOhm2ywWYRNuEMcq4t4Dvtv19QFLQ2eRIKKnNtUr1Vep0jD
6rRJgZkwEXZDZwwb+v0EEWNaIVyI7sWgUmh88gLFVnw/avFya8GvnfnnRDBRLOyQ1+v6tpXgt/hV
5uYW4ddsgvLbe4pDfiFJG0lwsdeezMx9O3f7x053JyB0leWf8zQqySoGNQ9OQyqCxuWLlDnXw5m3
Lo+Uo3cx2BinS8kfGgDYwbAtJXEjOa9f+wGcA6Lf07AIbAXUL0aMOa+44Af5CcmxM8yfToNRTDwF
SJQs9m94SB7jiU2tkjZIbdi0NZCUcf9N6FdXKlm+vrtoew63btPa34ARqmge6qpv02+DUgmHBEps
gN4bC0GB9ocZa/2YgcnmZdb0tR2rHg+A5XPzCmv8w1lrQarkT/E5blZDwKQ/VYwva8Vgs3D8Cn4b
rKcQSDiilDbcCA4rzHpWFA8XWiNZMMpNAHJWevgX4OMmwLTny3CHlQ5KOmd70hFrWukaxgRau/a1
5aUdtv9qh6L6Z453qs+xKx4x2EmPpWX3EA1Pt8iZfb58M+Ay5McYuqJ+MowcEo7L9xqW1w70pT2j
LZcUyEH8eDvYa2kYnPfB0bn4DG0JjTUICuKJ7xwFaDy6yymlVgaYEV9ebVkxMncvWuhTG+oIaB5P
bzyCfny+I6ABYD+OnVTEjajXlKl303osId/YYetnuPOHuo2Dk7afDQfhm9bIFrKCHhl/34iyvYQ8
sQIzF0bk3A9JeXNPzD+Vq8v4Iwrtbf1CqKa/x6Z/bzQzXggE8NyT9C0JQwul0kmgYBpR2AGkbJma
l6yJCcZ8huoNvng7Fu2znt9TsaGISBiRC34Bsfw6EAfufo+j8qpfi3uL43yw3rt2gjiIzkfkBKKC
7zlLB1Da0rVuaWOaOGb1NWWdrDmEAxe5UKz5BsaQAD5ZfJ42c2QpbxKgDLfJ/37sxo4OBmxh/t24
GV6LBAtjvdBg9Qnr1M6YX4yvUpR1ige1g/p/4aOKheDEQolqFWuDfW8wpewKLOQ14uGPDrqN83DL
r8eSXIaqqjvV5gICkSGyeyiYuD78SoBGo+BE5ILAfxc6DILEAQm/HTx32mcD8uyBNaxOlJCF1yEt
bcdd1TFIz+ckR7avrf0+waf+Yfoik7TdBEYgmKMWcWBFs4flpioJn0NIKDTavMOPLiRnaEr7YqZt
6I1hB4BGbLd0sjkJoj6KCNW24mlWApWpxUiZU+xZIFKvEZ6ZpGSu2kUHgezrH0VVSRNrRJWTJ//L
a6EXOobmjTEa2quW+HxZs9P0uNMWoplUOqQpMq5ScFiO8So2yIEMYwdkxsknxKew4aeVCj7qI1F7
L9MHj3VaVi554hMTc/+XKsbjTFFroaSLVeuMSHfc0EEcTBnVwkj0ipEDxbx8WHrK/VrxRHWmJpAh
WL681rrwbnSR2vBwobBgKax6Bb9wObmSrWmpkbRRrrV/TPSUjjcAWBYHrb3rITmFzw3F5FuP13WG
TMa5/9rLCwwmp3Gp8pTdwGyFzH9N4VduXeKSfsIr+gC4m0dJhYf/iB1q5zm44u71CuqAKbhHFelD
YTLxdg6zeqG5d5fgaulqWgefuh9S6eshFyo3M533jXurC2wabaGOBBhVCij+3VDyTbHNePDXgwPI
go0CfL7IOFRLAd2XKZEKarj/I3lW+RqLmHwjBV4YVE8yUFn3wtBW+mVeIrhbMPRbXBugKiuVO8Ve
97DVMMP1cbC3iryc78RnENWsLtqRwqsAphkfhB5QcordgQ3nckWsMV/P+gdbRxOo4w6sbSZXzP0p
sjeGEKQn1YJ87hLKlLsOcoO6egphI4m4EkbQew2h4rP/PheZx31MlQZwZTriD001bIuAAJnXFPY3
Et/w/TbD7B5JZHY0iPNmTOTZFsUisURDmV8d8OsEUvm/yEBo3iZPib4MF81Pij+kywY9CopA6nfJ
o66KPr09ISJ+HTLD/C5WFO7i27DqTb86gmIT6Pi93B5We+NN3F2NSGUv6AToXelzbSCFVH92+/X9
WRYW0+qlYQELaCGe5+mJPLaNF0hXJHBSq6nZn6+GGRvppAWXptvDs+g2ePi/MrZ6sMiIzrfwG1lO
wXJOybPwgT90XjTWSC6purovyu5uz8zmShzXsQSqq9aP10Cltd8VklJv6N6PGBUwol1zA4RT1g9H
480WCTRA3jry70JIZ8AsY689DmRpJLfJaE7ufRV5yVoZJiCkhhi6owkf8+kSqJP+Z/xxMi+FVXRV
Pm5xypqb5pzUtA9cxUk54Uhu7CyLrtyx6sfI7dbfE1MXhmKRAiLpy1NowRo025OcaLj2Dsb4eOGH
B9FYil/4090P767Ihk9rOcD3PvUMK7mMCIpgDrYeuV0G1rFIhpERvxlv0wUnRJXXarflU4QYTLQb
sIUKbErF8m7iOQLM2p3BCfWvyuouAI3zo/9RZihbfH9qe9AwJkwUHZ1MNI5p92hEFpw1Byr6dalf
mcsccL1DE263Y6u8z9UAJMtpv4cOdRtx7pZWEnssYkD7J3W6s01HoD/AAteLERZFIlYOZ8L9It7r
vLHWqh3pmM9IcCbonBaWHTa8HoEveXQBvJKgPLLeT5Ew2A6NqZ1WboJWoPiwNsD4KNsyMSaudkDO
maE6io96H930ZH2ux1+QYmkY0TzGA4pwuf7sw9wTM0B/Ou0j6Ya/x4COR7b5PSffzmmD+YzYd7ke
QLhHOrbrZ+t+D9fKosbBLKZQhqqJpFAaICpOvTi1BN7caQhPbaeXqoBoWfCGwHfFaj9sigPz4pAE
TUiFZVt0rliDL9kVaUDUngScDW+LdxzM3/phCCzSoFPn+Ja35W1SZgIvSh6xNisyrSA/6a5goSBI
Cw6l1mTnkutuPwQMmVIaxPuIwOjsdHltpzLGw21TquXC8Bsih9vjWEoe5LhYrH0i4crI96FlgDwM
Y8Bam1uSlrihCM/gimghaRp3SPNSBr504TFd44M0+TPCrVfL+HVo5m44Tz24yyAErjyALfw+qSnD
y/4VS75nuYR72Gv74g7oZGuQBlr5Ce0xVAEwWeFOeN4Z9YqG9C8uUy0Vh1HyqZnb1CjB8e53XRzM
Q0vkHPJFT7tWwnRTS7KrLIZY0dicYrC76mqN1ROm6F4LHtyrGmfBNhvnWf8Oa4HKDqKMwsJ+zPu4
BkiNcToZXrug7zAV9J3EeMARLm8tG0Qp7CDNx8EVlktjUtRIviWjJ8YQsz+ZLM2kFQ0Z4mwxvBnj
s62VskTW33humKsSW6I/oIPVoiBkQA3pz2ofIvPT/eqwzGUPNPeGyPYNil1iPTiOpSq3IXHCQGby
BJmW0kjFCaGTHpYPwoy8yLevMDcNorhyf9jpp4Y7khsSqThl8a/xEgfXcSlUIpZIr5kC75W/fgzn
28v7vZPZyJmDNVB2bb1fTFAkP0mXhG0Ko7YbE2FhSSc/8UvrtniDyhsEwd+IkWZmfy00BYTWDNz0
4HDCahjVLJmLr0pHKVO3RVUTAkMfDDAnkANMssopRBBfDq7xBxBDewo8GllPZYJAAqxeSxHK8Odt
pIeNWkVkXR3R5HEM9CrFaczelC6jmhcVq75gS+6oWWg8NQ2EDnL2If4ttjLdUkPIzTBd9f/U4B6i
g8GXyrjpQNsd6OBBxMllrbAgVhtNiG4xh8zl0mlZPnADLvRb6NQY5OMyFSqp6ix/aeAtAFOUiI79
WCEyyJACeMP9Pm31RaB3dqrODV/wcuQAU7UXv6JqLnkDiiuTZfpNuG80sUxd21Xep08Q+sw46B7f
8ythlnw46QkpCHwgw5dyvxw4MwwqDnegE811dMYO0BIOboFH+rMIIRF73tCGG/FJaPctkEU7GCLo
6UXOuHRYuvFAGDE8hgZcF66I32njOwc6Ecg6DKkXozwSKll+flxodpnkoEOIB0nDWz+gnk55iCIw
/HJCQWKcC8elzxdv+zj6xHO+SGN0pcz7SqtffhSwsaeX3o8noBjK4XgcZ7hAjN0Qwal/LhAV0Yi/
/kJbAKJPm5OccASe/4Fqi0HOTg4HQsbJU6ELu3txh1I+KPYOe9TAjGQBgQIg5htLMwUGfS5kX20S
LTKpvMpl15Dgkx5gF1bf8pGAum+bIoaxYFtm7TfnnJfvey2ujqEZeKgKGSvLIkBPxrhbshl8ithP
eBEG+CHBobC3F08NNOauIMuWUvay2vYtrka9NOUKV9DhOfs/sV8OivxQeaLjnnEGNAEWfH+sev0C
yWA7F0d6iWvsRK8egvgoH8X0O7XgpYaav3g4KVCSDnb5ScXYdGXH3O4cyp7ok1ws1J+xTHJ4r7uA
FKAlbozMK0WvOSmnR9Xru101f/ldMlTSn7eom278Of9YGSs5I6oixVbLyoVSFG6XkipC47g9YsPM
rlc2OVIAos3xdAJCv0l7LMinlHLNCoHwrZ2tXN/l7fwPSB+VPMI7K8PTKklXfqyInXD78l3n2Apg
Z2Gcot0q0jUqx4DYwd4fsAbV/fTSd6AauLVNcYD1ORu+WPzmvUaxUBIHJxIGk1n48j5IaWiADBeB
BlXrnQN5X2nf7b/LVYtUTBLkSEk/+hZkVw2AHysdAzwkjfK29gz0JXlmohOm85fy/sJBPhHwjfcX
cLG/AwaESbR8MUv7PbaGp0djGDRffPVCFFUDyOZF4mnKeuox/DS4F8UyU6CA+9n1mJbOSyPFOjkC
0R87yURWKa8NQKt1HrKX7xDkBVhC3E1FMP23An9wnmEw0DVNMgMV3JvgnJpSUxWUYulYiadqI9eg
zJwGTxdDPyAZ2GXv90VMLPJSz75kdZa6PC1oLxgWoGqcyZv+NikZBmrB0LMXeP9sMRdFoBpdXhTO
9BYjl5JRDtNlv/uOjdiEon0iatEyVvXQP78XstGtDOgzf9MT1vMhiQYSQnATAEPVSz7s2J+Lmw/1
xIJ2ugceh99/iLxiiSRRAN7y1tLnhmAQqKOvsgZ4XF+Nv09tuh0SquShIOLJihUrFGpMPCr/PlFm
jrj+L/JK100vIPiGDf3JzJIZTcEFnE8Y2uiaO8IdbPis+6BjgbOEUNR2Dgr8kaDFzGVFO9qx/7rW
5Ts+bu6XcZHWl46UMwG7dGRCQrzzHpKiiyOFQJte852WNMgU49d5uCn5WV2QXdMfYRvbdpbsNuUu
HG+CEQyPfD3Q628bfsmKXYHJSRfizn7zgTMzHIX1A6AsYyuRIsAV7cKzy63aonCvhBylcCoAdTVF
6t+MwlpBS6rDhQizEzSXg5tBh35D6maTZ8gaH2Gm9gS8ZT7ZidJp7lg8JESvw3KTh2oBXJJwnryr
VavaQJhTL4LXvkK3MsRyEas8BFr3K2hcTL6C+bSDv/h2inHhOmg/8iofrtXdbxy4cK6pG9UZVDQa
gbQJdWvWKFyo9dzmLvxgrRT1/pnYsu9ZOok71PPrwIlVN7RvfRlu8SM6twLVZkEEzVD4osedXFkR
K+2QpG9TyKr9EQ6ZLt6QW/QPLyZRD9EOO8fS+XpnKD+usFg2Z3Wb6dJQXDQdRZpR6AK56Lx7hOTW
ZJD5T+Q54iaVB2pARXdzxHeR7KD9/C6uzSenxY5QMrMx+7jfqU9NHq2nQ+d3/G4p0Kvhw6PMb0Md
fmm1saZK0w+vdS0u7KBH2nNAF1ltFVUX6y0EwvrylOwhJn2Mqs0Xed/WlqP1A/4D78bdYuyrZIOo
Yh6FG9phAJ5qYKblxtMzrb0WVttEo425LlWYOVY20oNIvGDocy6z+rlWtIJgDwRvvZOOi/k1vR35
4hp6hY0QSaRkaRxms6hfHiVAixmIEOip579piFKTYiHFp7YBzLNKcM3XbCqTdTdeAQXK4ZrHpxnY
6FgqLXODWuXMm74IMn0aZd4iogYkC20DBi/7H6aeGLLibvqBEXVMO8lGWQ7AZTt3gCTq0xrTsDSh
dtWYz7r9ESxcaNfAFgSAyl02T/CPn2yhuNABqKCnkXxQsNphPlWKrOCOrsEgfJu5dU3vQl/B0mtW
pCO9U6q2oKZI4g4m+JWr4+wXsqIIQa2LkLqL9O9iXLYtmXF965TRgcJUtiRDu573C73N7NGTTJrr
PGKrX+X9AYvP8M8gpqxalQGqlJgUPreucWr8O3Dfn708EjU3PzHpuf3LnTMes/XPwZ9NCYZ1uYio
DbTOoHPjId3ptUTg6OhvXSBTWsn0Jq/s34aHqMrZeG0qb3O+eqd0DXR4ZhdeiKO5A6OEXpvVa/J8
u+mdDnD0cS51/dK85mkkWdlIFDoL49CSfc4if2kiEq4ChSXAH1Mh9QLhej1IjwGTrH0bG5Dgqz9I
g9Ongq6bDNm1TH5lzVOYFx2zbxtBGOfkhBg5ldzvdUfrdzdvmgItqOaXVzoAL9GQxZxed4Oxxrbv
flNL777cm3hoPKJ5Wt3ebagXu2eKRWcBPoE/uLDfhPQVkxuh7gWl/u+pB67BwTVADR+idJvYx31p
sLqK7rpQULQ2JFH67sb8vC/NFvzCn4v6vyaeoZDEv9wgrNZ2EJ3ibbacKFV5/R0qTJhkpOMQ8Kka
m3VrxwjTO22v5IkzC69SVg1A9+ipuKor0OWFEYcz0HtcMc8NbpCu1njCRpQjwdn+rd5D6L0b+aCk
gpmKhp4R1WHVAaTVM9QOAIFmWOtvDL+PmS0gFEn/CteNO391h4U/wtLXCGT052BfwpDnKtFC/iWO
l7d1r5q9IQtHenyvAVkSvdBqPODYm6NETzjLirgqXkA6kPFkvcZ77gXvzvaGU9C3gTRY8e8FDhU5
0UOG0CuJLBd0CWtnxio+uad8ZQlj/f9gs6bOowSliyoY4ZSUOZUn028DSUxhi2USCUheClgrQTnL
d8UqR+x/sjsGj0maR5efjBP8lhxr4Xqd6720mMebHXEsfvHiV/0w8g99bok/1Q0NGCpbsJe1mKJV
5TlsBmE+jleCbzE/3XnhcY3veyyAJNIub/KwtTqu3JiJkvCvm6nzS9CyutzNFGxSrxmpQuCkYUun
DBrGd9mm7gL8K3d0B13SopIEdmGZwvdpdZ76mJbpQiYbBGByqzHNEbxUy2PJZAnaLD5JoI/gEXQ1
F+vhttnZrUwKHlyDot06glYz9wzmi1JBzHlS2Q3QyX3amZ0T01/RBnl8qtmMRmmjtwV+4Ae9H5s7
LhzblFazaxxQPQagdhW5qUbzomz3snb2PDwtSI5QlRbYcWsDtDL/98gsIKDwa4M93aOfm7AkiRCv
27Icy14d2Cl0H3Hg3P7TwNebuoIUfy++ttbRflFlummwr4i+yihVCe0bLVbp66kkEeNAkGsAck4y
S1XZKjLwI9VIegHEzOi6QZV/gWgen/da5e0VVR93LPRK/1NoBjKUrQILVgZfWjHh8lpFrsnFwtEY
V/B+iBmT4PaOViX+mhvL3pOyD4wcHsrSZQ9k9v112aS9caj3G0x0W5qID8VL5wV4aqfHA79yI2H1
WGFiG9Q747pTu93+ELhG5bGqwSYkqR5frJTkXOJAwkJd/5zYqMPHr2jMUEF1enKky8h+nFmDjOyf
g/oC+d8jcOY5tFYbKn+UPbUexPUlGDmE5BdMsdELuAK2ij7GC0gk6bQRTcEpuXrqgR4k1nWbASRr
vWV4AzaTrDVOc2UvvRVOM1tiIb1VDDMUuw7Xn+pldJAIl2SwBmhozdaw5JuAqEEvwk1tRPK54vcW
pNoUlPYbn67YWxYHjeMgZjddxrhH5575VqzwxlpjjKC92q4kOGHBZCEUoHiplNrLuV5aBJspw+HQ
bQqUndLNPLLREoHA0UL/5fCcq51Yzmuomv5k/9BwsCGEp/vWIIEANfCDhzfQFv38Dh1fRJMer335
BjTyJC6tPRUs1+r1b+WH2ULw19zYjNrbYpzKCFz9GGv1ECOaCs0rOI3gudVVev06c0C4puoQ4Hqu
N07fXcXFouMkIMyjDsxCwsG+jic8nXa3PiLAh3JmBXLm5FTOo7NycVK12R1XxVag+wMv3u8dfDzZ
c0zrs0O/iKg5HOPA0uUkDJDbj13PgB2vLY6C3otbEfwfS6AjuhP7cc6SrXn65q9913Eh/9SYW+ke
Rlm8F+BGBSxbjyVVZangO/ZNMWHR8rglebPk5QA5ziG4C+9SGymZhrNHRPIhgMsORg7iJb5KEemp
P665wr0SPW2XDznWjpVObPSwkpYd8TLI0mubnt6GUSa7TiOKv9XBiky9WWlZVqAZCwAXYr5zueOg
ngFqK7g0J53ESq2l08g0RH63NnLSxfq9pYgb0/eqPcH8GvFDWKz6bzm/IsOnGEMMXT5IvkGj0Lhg
YsLTTIuUb1WHHsrCboRf/PRFnwcu65+Zf/cj9Glbob0v1kg7Ff9EItfmQOygaJRWVNREoMaZrTK8
Xtrl18SgnfdKDzDGYcamlHpm5hstmrHKhdO3PPmyrwed0W2dos4W4O5Mw8CPFRVSI2fRpRCeEO1B
0CNKpvGvjMOiogoQncD/p/qizMUfj5wu/hIpccSJLmf//nFFpHH8T31T+rMCVraMJCGVGeXzAbp8
nXdKpHHbcCmGbsQvm3PKevGLyZ7ZJAt4B9q8LYWhYDdDvWTuO7ix098VJ8zhKpGJmzfkIYZza0Dd
W8WFLwGjNN5lQprzD3pzOU6j5fFR9U5J0FAEW5OTWI++QTKf5B0U+q5qDc0Q83IZfytDJndKrpe+
DwQkmG37FP/7C/diLOqgqeyD3ajvzUDttEp+rIjm7qUbSc2XHRIcqo+Fs9e9P1TYTqqCdCme8ZxD
3f6hr6r3QZSk2n5fSdd9Bim/w+gLKwfKxQHx2WLCeKV/UMsOb173E4UKhS0WXmyNN5ef5m12GIUl
8gg9rHzosxBWuyjTrlVW8lP46M+tF7FkgN9k6KwnLpirsj3939crxaGHbft1SrxT5LW/lyTPDJ7B
/NVsof/a+d+FJmVtB6Jz/BBaM1AxLbSAjLGj/wZfDgYeJ6DAABOwzZzeO9jDjLXD23AJ4EGxotx4
hfwJLkKFR+EERrBJzwYnCta1gubRTWd1lmy4Ke4n2saBT9D7hq9yF3Fd6a+hrzWQxL6FTyA3zgRP
1IeEnH1AHP4v15Goq0tqQZfiZRxg8wMTNa0PNNDZXR+9epKSeboA4fy+7WrVklXZqNYhJe3BUFui
LELoXNs+iIZ5pqD7zzgyVdvrNjY8UHZWzoPqXrehbtlmbqxwWbLsO6YnO58+1AyP7ImsXJ98H72q
OJIHCRaPrMw8QzKCWoRctP+TU+fPixikvTOm5BzZ4qWyAMeeR9CFu5IcqstnX7ekXw7846/GWePt
8uWDH0/6wUsDOpG4L70tfQ2ojp5jxaPSk5z24SYW9G6yMkxYLqn28CMu2fmZOsXvfWGIWIYXp2DB
H2n/lXgwD1zDXL/ycjybAa1pLa6xV7s06CoAzPyAXQoedFAgiyAivDRfpKM3zwJ5pOD/Q2Zl3nNC
k6tO/RTUTAanj9J7CUuDTck9ulfAMVCO0Zl2uae6sFvFWZRIvCSxtmuCQC1dsNQq0kAJXXRhT/aU
W3rmY3f5xnpktykAkLIhblrwMrent1X0UfeJdOCyN2LvgQ8QO1C94R2XOActSxFTN7kJyD5MP1Xi
cDPSNaAIQ1R0rUkQ+a0/9YrxoL/Y8keFa9TJ7YShmRKJr8VQH6nFCzDp5jM+1OIEK+wys9gYvv6N
VNtkEwu7iKfJWq1hZh2/ztQZTWVtDr4n5oty0TtSIeFHLhpkp4UWo4NqbUBviyrl8N8QtXnLIWI5
rhz/JyDjLbXNWbbXSwzHwqj/PxgiDzoCnBxwWUEcoow147pZY9Per925jpPoBtostfio1hq0b47x
ZyXKi6lQVXd5Ch/xeaTV6eTAaHPAD5vcGKUp3QxsRvj/SsZyN182ti53lGYBdrYaVRl4wRmjQiVu
8Ap/tU6j5RxU+/ezg+w5mZZqDqiOcs3XoozVVMJJM1ivxfuylwvETC/M4UpfY51pyyvzt6ZX0YtV
ZYhwja+28+6ZYwpSWb8fXgLVhWPE043R2XDV6/dApwroas8bmiytG1coXrmf/ZaNiniAga7en/dV
YoqNrwH1M3Fnk3AwahzuSLG6N1HliaWYaMKTqScYXYLJHiQkigMuWNoCgl3+c+OyPizb//D/Spvp
O9I8f8hRinA5JufNzp9gi3tqPL3ys8VRCZpySFNWq3a9/p2rnqPZ70Ug9fRR/rRnbw91s1KSC97g
BPJa6U+osj203aXZU6oUsbhou2m/Qm9t7M+aGRd5OcKxYOEWZ26yEGwMjV0+VqKhbym4xoYtcETB
alrpbK1EagEpsiMc6xUe/ZrTCIp1gkpjN5Oj1Q40gZ47iNAM+fh6C9YRtngii6f6tjNVYm/K537z
Ppy74zROJvWgeK3vugr5quBjn23Eo+bk8Qs3eawtxxj3X5W4LRXlS0z7avaOW5Qsn+Q7iZZy6NUD
9fwTfeqdkrvpnrDK8WPpjlq5GiUq/+v1xY/yJZmp/zsgNKzCKVPFkZMbF2lPjBu62WkkhfZE0ltL
TJZPxE5X8SeZf+hUCKxOo2vX3Fl6Qy5aSrEM+v0WXUAs3uvwhjQDTKvce+thDU0cuDKsuIqptZ/L
y/ef4KKnwg2a7IuzJPYs3UOg8z1nsSC7E43yPeRWgXOxUSErDghU/6ziHCGTPbG4k1pH+cODN3lq
ahl1ONVZwNs0hg5DKlw8/0RV6avQzTi7jlKReM4uSM1+RxJ9GIIBsPQtUgaMhbh0Vt1XR4ezGR8/
AltcP/UkBuAaQ3qzOyaF7bC3yJ7C7bN71G61/xxjxRdIcffcHT6ZfvDgYU0MlKbBJKgkO/vLEE0k
QN0Y3wM821Z8QEN9q/AkyI7WFbh5xxM2bpnO3WbHVJoa+KeOXKaBvhvX/RkPSj2uLFscGJJfzaRq
TWUjXfTlKPT81JQGWwje+j7JVW6tjLTHrr2KWSODdkwbPXKAYclJQUyCx8lcWm5eXs0MUqrWtCsI
Da169OFxRcF1Pj2ZwthCvw7eT53dWLd2XSNZcqGrR+WxjkxxeSA+FibHiYUO+FtOzjvD2bIl6dx/
5yg0habJRPXCvvtk2gge/x44pu8DrVXt90aibchO6GHVdMKyCGKZoGIeaan+QxAtrWozr++MK/Rp
ysNpwKLCXWlQb+si64iLbJB3287HU2lPhiTydRRXARPrZVLf6tBf2dGIMgkDYSW9Q451zmRS4rDy
doadn/iem8nXjAUkmUYXHfabRqyhMxnqY5aUUQkVxf3xOa7M3NKtAFzcXH+MrBKp6pu36TNPoU1q
10GYoYjinsgEB1kuE4f/upsuKfIN6GBOLwzlvBlx0pvOMdeT+FaK4KNBl84WCne2jrSxiwuqESNp
sN7565HwPG85uy6y9jjnLUdP6sXtD4Ce77+TQYJCmYZOBXK+lrFYD3n26NThpk8qNbEXCebh4MwC
mxt3R9db+bFgts5d0u86uM6gvDsy+y0Qkhfz/QhPnbuWTFyfxldxHsbpIqvso6JaT3pE8NLb/9lM
1z11x7H8dTkuRQv8d35ypr1bdueUcK/jsZhLGehpdD+gr9ij2kDAJvwDyfhOjM6pEFbXK/KANUGD
ODFGVf/1lGRN41PVi21M1kawl31A4lP4YM1eL8y1lNxYUfHOb4HFgd2ukAW9dFfSLRP9U0+/pjkI
8cFG9LsD1kt+0VpgZzTgfq9IRPqXXAwMiy1egdxYI2fC6es4T+qP+YVBKJe5ZNbYfUlP58lHv9TE
JwBMI03YEVE+2U+AE95MBA/VHsJ/iucFkf7vguqYosiW+nrrwoGoDVQPR4nDHo9Vu1j0k4k8iHGA
tXCgWPtZh8qE1wmaiMgzmdZcDFn1No6FWznf4ZEJ5uYNEUu8MEZco9EfgMPdvKRm/p3ojEDDMH8N
jxVVaWBNnAxSbUK+sYwgSPNHTkhjaAOx27Hi3FRQ4JTgG1XQSzE86C+sdinJbnBQ8+5tSTu5pIQT
HrJZI/zFOOHPithxvYCcbUA346YJPQk010jiuyEvcAYMTHN5rN7J+1v03wy9sd6uEtF2lhA7FElf
dxYIUBVx7UWwsdcaHM0SbnBVTTMPm0WPyRI67aG9/5ZJJ6cPKAWLQlGvWXzUeWzZ/y70Y2H50F6t
8NR//Hkg7b3eWi/pfWsQSXOymUK5qP29CN+rTEbRYS/ZLVNZq54uzrtJBfejUFHCaGTHC0PpSDVH
GplQgtbV8gx6H0Wsvd/Zyp5JK6c6/GYM+slYbNyGDzVswlLjJMeJRhT/1YsvdpmKFvXAFwaeLSFU
g0R2yQ5AmPAd3mQVXUxhZldm7g9puBxkKn2l2/eXCSUBeYEflHIBcVRbn4yvCNL2idRxfyyYKLGc
/9jBUVGMaYz/0TSfBTg1PyhgW2lK6IWm0W3Q3fSTb3oMLq8Bv5TyKYx9NBtHH2jEcYtj/6HG/ej0
ndq8VVzC8oUGC2E1yCHe/QbiXZ9x7knmOjuK762pIBlxgcTHkBGVYUvfHns5twVcSPYWGSaFCSko
eR9Gj4qQ4BSlSlTL2Mg+V1b0zadeytdv61tRMPMJyP9UTRjBN5nAf54bDXSB+yZd2B5BTe2FMztc
dVaWz7qZUP4LS3YckzW1CufvOBWsZWEd83jJkfqVvHC1a2Bx13NmFzXiPx7gui8ETcZ0qGHZRWEI
q2lfAxxPhy79Sholsc+vYl9ljBHqEr+I3tes19EXVW35fdEAx4zr1pccuzdGf8ycnBxlC5aC8tU9
3mxXTuZMLDu5Ky0miWdoy6lkHQn4yZUlJDrICoor7mniLPjzqnpVfNvUS+SGfAlYID+TPqFa/L0i
kGUKiFOnXy6N7FGJC6gL7IugtcAdBjYcK95+Dmf00mHyJB8hW5kgYoZ5QPq+OXNG/UaCfU42H3xa
3yDHEIsTaMPegl8noLFjOcJ5xYWt4vNHUWYX0TxO+hvSFr6nTRfT/0AxUpxyRE1XNpJkXoyk/xIX
FdjAnNN8FVH2T2M6bEIHlSafjBd2SmKbThK68g5VmgL1YB9wzbW4mUm2WYCbQkyqqHZLxgrIB6wi
rgCALHNa23hWdifWfGZJfE9dLSpiabzumbhJ3hil3aD1wdMyDrlr7A1RYgT02csIdNXVKkIHzidu
XoSohgewU8ZWcqoZt86CvrPnG6m4HS6woMFuPpXEbCNTA2ZURYsluUFVpGiOoVGXKUX898nRuZLY
oBrRBGtn2FbDDGz3FzMLv6xl4h6BdkW+8Q8cbfbbNiTQmQYcuZ67Fx/JhJ7dWZnEtdFWs++36sHT
CkNp/cgZrDDdb+IVuQzlx9QDeimfvQdTqgwnnKY64N0Dhkc3jFI6+PCCtZD5foe1TEKUdqS+UEBZ
eWOyoC9UdXd44WbbndYuDQi2fMb8q4SGNmPTq4eiZOU/nCI99vvKiQln/0qmDq2uToUHBedtoANa
Sc6aSvc4tUt6U7bgpMeTWmt6A7RJukokIgm2jmWp85LdvvSte7NBrPAYrpq2VP07JD/w89kPR0AQ
eh2Tp15AaABjiIoEUWV2sCH+Oqm0pvJBI2hvs8y3g5mrGVPYTGnT7K2y501APqsGD+/H9SQuZa2G
BPvsIg4AEnv7KxA7z0JtQUwNRNyKl8OQpUUx5AZtQNqOwihJIHxn+Fu7HaOsquDqpuLmldR54kFP
zQGXlHVRUzMLlCSLs8Dw4+jspHpxK4leBbqW43x5WLMHh7RROBHp23lxHFY6k8ttm7aM+Os4BxG+
CNyHpH6A6mDRDr24NRaff98VzGbe/JQWZRCUpUVqJECAB2a6lU2hIqyNLQC4sAoQbq3zPpxicnsE
Yi+dGQ5QBYLFl3gU6+37UVaunCqh+wcDADpl+7HCFlC2y2nWarCBomhmwNjWpX/IHhdFanAJDvKF
9b5LJu7VQ0HE1rxAvLkSSTDJCK6I2iz3g6TyQJnUbnj5kXShuz060Jo7zAwm//IB/bNE2L0NUhaC
sdtyRBJ6/SM38dBt2CBoQOrYm71Ql0voc9sMnY/sRZnKS8TUQJCCgShfQmlHq3EcNkmCSfoCitnu
yI9DXV9sg196/jNm4tlrHab+6v6vZlHa5+AOCSgDVLkoAC0y5d+Mhvm46rquJYAS6C5iCvAy5Qn+
JUiSFRQyAohyFZGjTnk8FescoRoDxIbjvoWyecpXZ/UZyd4vJDATPrvUU0N5uOf7qn74fEH54iV9
JxdmSURGMCjL4z9vzVG4mVt6Z68mNeaUBdImS0MviniPL880WZTi6NmkucWyhPwToFxj9ZwPhg6k
cZKgI7ldZ5XEtkegseNwLcnIwyAPw47aYWnqPW5Hou2VK3JnsfcqRoBePD22UjTrtKKyv38Bhzt9
BX8G2gGcEiXAE8F2SK57CVYo25V1aMzCOgU2MosQ9i4bsl6t3g32Ec87eptJ16hi634FejTi+WpE
YMqSFtxVo6mXOkXNExThpQJoF8oBwhC6VckN8rLU2LbTRjjYGbjqnPh4AuSt5uK/WIDHSO30ER+l
WGvbT5ZQP+iRthcoWe2yUc7Yxr0etPcqN94H25WsoNpZROc2PM8KpvTIHgM2hpKQxfGdwhG2yw1O
AA7Po0kt+TLdiC8XWYcjPcEXAW6EZTsX2e51LNofvuC2TZgUhf1y2JpPj+0sa1QkMu9xyUTv1tcY
IFGQcWsP9oRL7J6xp6EkJcZWHte1+2Yjs05ot9GPZNLr4E3bBizuQbrqEK9xTeM/Lh1sR2EdJk8c
ZdDOCM1LiNoYIsR1vj4jkR67PWUp/B81ISnc3jAlGtc5jmPjTJyIFlm9kKG/oTJ0jdT3DDOWOGA/
LoSkEfuWmqoEtN5vloFdVIsDBEeinp67kkuxm/vwG/lFWNYRTwnPW2n1wH9U8j/dHrb7K0X0eT+U
8UZDQdpzNji99GRHbPs1DowSFCWdHi5ur6r6Ep3E0xmdAOdweYyiaGwA2Z/VyLDAjGJ/9g+hTLL2
IaqiHqw2ERqauL5bIecGqcvHZb82jpkW0f9JgZ62K1numF2eXSZuUjUWCVr39d9WrZWPhqySm5V5
ng4LRoOlmDSGP7uIwa3/W9DBS2jPOKKrwRTLJj8RzwO8qOlAmSkc+SBgeaPKkQtvG/NMDQetQ8WT
7U7KrjH0GjhpLEx76KqYU/2DxbHMracykq6+OSlfCU9UBRl3dipMmZFgFBMN4eT6w8oW1jorcAIP
KcGkxPMF2dtlzKNTccvvZ48G/gd5UceLBXksCHEWt2jYW5n0EN8nJcDkCxxV9TtYQHKkRRDEqLJa
DKfMsdgxebrl+jYkxh9/rRyOQqN7nPmeIf/Uf7cvHjLe8brNRkp6P/VLxtq9xjgktncnbHQ40nVJ
eG+Hh93oRhsPqzNQWbBnMKwi3evYFvpyPqsgHkGwIHLKDmrQL51eAhCfZApfHtXyOmhTM8yVcI2s
f1W6+fY1Y5XLiDOScUBUbtjdfFJjlgTUWs9o405YskwxTe2kIwMplrIYOZ4+/szXfS+nMIMMynIa
qbPA8/klHpTuoGgBTJ16KVkdN3QXSkkfTIdQeWS0s62bZ6TCHEakyZ8XY1YBqAIcdHxGJYmq+Mm7
trXmi1nGzXxM9K0FuOqCBnVLHJSKGj41XX/9o77ih+fCFxUjKS+PGnIaRkfRrG5WjZx5VERyh4k9
V/V9HjoAbTvu/Uw1DoXgRebzLi+keaLqkAsf9MKHGeiSJkjAfJSTeS/FImOcxe+O5WJhmVrZqEcQ
eACDrjzybKhhlnfJ/JY+m3PPeTauU1NksykzOt3zLRKKh3t1PZ35AeOk2zUchvMUnDmNQeTgSXEX
ieX1E3p1/31ByAey6DI9xEQknYiiOJH5nDOvmNxE9zScOD7dFOmg0gVrEx2GRBi1BK2AFkbzRArm
g1+UfPL691Ik7fJPYiz3pmx6fB6wIW96MXFItrbo/o03tgWUrkhQZn6J0iOBCNRO11U08Q6f6G0L
ExLryEfYNsJ8AgHie9T8o9nToKIh5Ro31LpHg1x0dsYUM3aM9rGddEkNZmlv+jmAMpTkv/2jjFgK
L6zli/ZDwvHkj6Y30NiBt9roWQC+HgJlgm3B0Q6mGqUuRgoGKLOI/PahAYtRKXFimAoXhsg+Bc4j
I3aNeWJU8RCH7EgmeU8zUOF/Uv41xnrTFjFMIXAJYwm1jRM9PfIQ+EbDuN8FLodw8SLkV0lr6Rk0
Qwd02iRfsZSfbXlEpH9Afv0VovJATPhPXXX0yshUVik3PuaM+rZivfiBOXcheIcHYpsj762Vx58l
dqMM7yMoPxN77l3UgMNM5uMblKRq4epfjnX2jqt5HUsRMeCRYme/3dsfWwcMVfPw70I02p8f2eoN
G8Cbvz1X6NP5IoFewwNLtyOnU1y73/xK0ZuSKL0vZdwD138jEZyGemnv9CxCXF9d4sMidcBQY4UG
glhvVznLb/BG/RNa0j8gmCbaZwSPBjekn4TmuBf1YTv67HzNNzFx747pudvQFY1/+niq4uSFSzZl
kgO/TpWOX5E9z0aRszC//yZGhl2yBY3Q9MVQWvAJhoHqJzBYoBnpoqhuA/baO9jTb850NuKF5Uzr
wLM8UBJKr5cIFIYVbT+3Fh8rWA6fTV0WaOfv6UAqiWKsa/G7hBNcLrkYhxBMQ+qEPzPzOzf5ICsX
iU+9It/3rICwqwKY0thaLQVo+epNKVPzB2qrHn4wVXSHFfZZ+pQ3eDkbtuEiTXCTeReh6wUriNpV
FlmeDaGs5pHTZ60yTdbl9/EoVWhVJIzM+TTIArGg+2kTGWC5GNuaSD9szKuTpgli8X2Bd/tJL3Wy
dBZXWsK8Y6YDeG4sgWwtDzFQd8YYRJo8d6m0U9NdzicgBqcednGvThyxqIEQeN27SBtSL+dZNfPr
5H0qWtOLmauFIPlSxrkqwfUzOSvyU0dv6BZD82Y5KcO7p7twAaEWRsIFpFdjKqAQEDhppz3z52tl
zDCqdyU5VilZkpMmn+DXB8HJ3tFa/JkdhaUQlLkoNh+zrPNiouYJuEPb3XSYiUxbPn9kA27EFu9Z
jhkEVy7lVKcHp2tA9SvKbO3EO+Xa0ylDq6BWA+XnP1S5hKDlODcpACyBjga+fR0/fv1XPD9OHaeq
5CIs8/ToM2vhXfKE15LWlPv4c26tM5TMZrpuIvOuKmlU/93SHbcwxs9uZP1tFzRHGE3ySS/tnAbN
53wrL5AyxBT1u+NVuUGOR1dQOWUfgHhk0LwFejQlulPDvb9RsoQ+lptUZKOiLLScITAGEAZ+a+WD
/MLhDwGVaMY878+z6UoqnsHDhQy9jA9zYY5yO1r4aAXjPZgpQvSa3nnC3aSaAClaRjfQm6w+32mK
JKzAtRSVk4YgqEBQwtt6fNPaOqoHciAlkMyNGksYdT63B9Xq244G/CeaedZbp5K88te1MgkCW6FI
LPikaBiIpq/1ng1w8QGFCnVyDdudHb7TmJxi9NtGe+Yp+IMS/XdzYw+gkSgi6mnczYvETSPlTnid
2gylqBnIjAAkQ1JM36JgCsZuVbFw1s0cbP/AWEyjJhG4z+CfSEGx0gMAwixyYveaZqNi5buZFa8Y
F7RUlgF++Mr4WKor7Cst0Hs5lf2jEYt9lUtI5ew3B009ai/19sc2qGEL+FhYZRNv2VIO+ELxdJbv
x3vytgQppzUkesvtTBPAi6BzTk98osp6+xmvP6xI9oBFy2S2gptgBbFGSLF6qSAF4FZmO8/JjjXm
EDDXTT3+lmlBjZDziT5gDX7VDtyTSqk0IF5WN7sHutD1RYeXpU3XG1gLHPZGFmp0n+E7qJDVZOLs
eDm98D0kRcDV5dYdep2trHnnfO5jcMYt+GRsPn2TkX2GVe++vh6jzaMuw6RELvyt/7zyKXAwkyP/
erS/USxBNxpF0H7+O7jT8u8Sl6Jx9j5Qzc23HXWQfubtfsucVITIb3naK9XDzd7rNrAHXxPvnNyt
DbbDZl3WaLupK+vfGhj0Itu8jHhdA7vSlh1wqNBMluHhZJmqDV/1WNRs3XWicgMnofE3OKiTUA03
0WugexfTQ8dA/KtL4KsTNn9gO2NtpKIt2cUN1az+K4IOpc7/8c/QPaE4QE2IeuD2+v3XlgI7w0rk
cnt0h8WYaSG6+utVukDrgmtFvLj/1l4MfKNVUXFcsHW0U6AXova8sBFIM9L0CZdxE717n1yzwGKf
Vgmip1cywx8K1NDl65T1SpNvkjKBDoIP/enKViBhVlccjwAP8zUqfMAVYbXOkDC1Ol5guQNSA8yF
U9DQYA/TCWpZOB/a5F/deIjpH8S/kSB/jQv3pd8IW8yADmpbF+4mWghYSOdlr1294Z7U18HB2VLi
WUfMaICS3rMxmUeCqyJN/tqXppAKX3mmeYJxjAxhhCxiFYDlQUbXajuRtdwax4vu7zBAMIxvCJe8
SLB093WBlJGLXTPbm6TokX65lw+odjvgo72FoGIcV52AlUqjbiU1CTuG3UUNZQ6LozZDpgrBcj18
yvnSCZ0x7D+/SOpuP0MwMlMZeZUcgc6hoW4CBJS7p1GH3HhSh8TX0ntDvle574zfst9KpWS5oLLY
lZnZKKuWwLUGvPLPMt0ftyV8NMoUKrhXaG/w0YJ5Stn8GQFHRr2I56TNTdBc0R5ANgSRsuY7BfWI
IDT9rbIuN56mdJTtwwci8wecR2FfIOYstM0cyq+vE9usCSsfto7QpSALxAKTsmqOmDXg0FlH4fcG
SzDQBABBQxtIEavxkVsA5e8voVdGBZWHdi+TDzjxsDpVhCKEQ1MuwolWO64NeveOQDP2TniHIKjx
E4GVkIcX4GqZSewZMqvLShRISGMJ3fa0MsxzLboCXQFc+ilZ2RfLSt3mYdyPJKeaoansEY4AtPV9
iFV0gzm1JKhxve6WLLcipUfgGVN8hvOv2LoX6DaWHLKItmVBwJqVmYvUHBpNPYUvpJG27onh4BBB
UQbrNZV0QwUCoXRrrcJPIVwEtrk2j/0uJ5vUgIig2x79EdXM6lEbOsBSHPtYR3l0x1RvDZBVjSmr
5iAm2veib/c9rHuG8CrKhMg6C19KMlykxHmowXFRTstNDip7m/vDxpUCzXxzT9JND5fdzdW9KsI0
XK0OG+r0UgmLDtpLlHRrFRruLN335PA/RCXxJd//xETrb1Iybf3xuQTY/HUjFTTUK0p8Fe7iiO3V
0AwzAli8QNCfrpk7kVWN2XjSODPhpDhfMAiAEPhNZikCD6kw8we7B5f1+wzeCdQ+/ABWemrrhEwl
6OwkMfdGD2tGmyemE4+lUSX3B6CwkNuHR9vuGyfJeB0mrM8ZAC3oyQFIp/2pi8cP/ioeMx4/clDY
le7+zALV5UE1WvfToZWZLg/ZB0ZzGdIJrkbPUuY7Z8I72cIj0130KRO+gZE9MWJqccxe06lqv5V1
67R4H/BTpNFSf9hc2jusD0B/bLuTHWHXI7VFL6WNvgsya4nP5vP7Yz2TjWPao0dbT4Cnm5ZbXUBc
cQ+oDxk8QMfYDkpe6L8tyx/INnJt4ZNJqgTaDwkgZxudrnX/sdS6vYPdFBPbnAl7T/pUwvqpsJim
ry050GGa2JEusUIST42ZJZ5O6J9aoACP2TAmXaynFs10bkSV/UrTx4FSeWNHlulHF9LJFal2Ks5u
ZEga63YI3NpB9D618ryRolxuuPRSPeefkQJXw45ZCdkCCdbCYZnwyfpHy7bsDWlFRxKCb0lb0fjS
2sIRGVwuGrTztIgiV8F3hlY5iPYuQXQZHoa+0+moRpRzN/FIZG3opSSJcpwH/ff6fo85RioKMQ6B
T6wgPBeapCsI+G4TKDIjowBbJwohg6RfBQAsXnIA+H1hPRVvXSK+i38ypvYdODyAKZTY7CyQOTZ1
BoiG48q7KkFEdF9wF5AHKiQ+qAE/mvFdTidOo8O/0ac55KsC4HVNLifsRzOhGDickGMvHhzq39Y7
MbM4LiUJpV+mb75sqxpeqP1t7epK4BaJnlt/AzwBBLQWmKtkOs/fFhGkOBNFXEb2e8YZdwkqTSbA
uaDcYHZSggPHf+ooqCG2NJusTNMCkJyeraXPOF/UqkTIINokz3j8zwKfAwmbiZ6pM9xQhbTrR+DI
f8aIHZKgIo0ledwmmFiTKDPtYzegGAjYkX/oviIEZ85OS09Vll5S3gDSlJvLj7uxmHDNTt411b5S
k9Hv2X/vy2+Y1fX/yHpiuhcg3s3icKl6fm/FNAlq49vPL9lvhPjyiimqLgVhLrmBJQ4B+353FIfe
GCgqfg9/+eFYqHReR0ig7n4qleeAVdJw6DnFIDCsTW9PkUIuNTVh/TuK+/rfzcM2A9SJl+7k1Ob/
e0SzPwAW2sSsGIzfukOpd4/pomKRNzcHrAkaurUOUD2Kfbdkcwun+pmQmC81GQ/1AmNXRw/jGEGv
27Z4wd7KLaXgYAbvi/RBgx+U7nArUCjupIrcR+OIWFmlSizNFE3RlNAjW60hu0ynyvrjKcyoTRDj
Wm5U/cyUv0qKGIYZmE/W6bk/d2Ya87+vfB3MbXzfbEXESTgcwNJjHJ4No0p0pf8WsLy09raQL5Dl
yG19gkE7Ym0cahzU58eFmrcuL8lXQf8S1b+ROvJ4vq8sSSf4PKbVoUGmdw0cGdHNWKyqdqGBa3gu
R2RkDZs9qHq6HlkmeuuHjQaHsWhSmph5mgnsxLTghuM/UFE1hP/cX0SHogWcwti9jyvu4G/cWMp3
WpHXd5k3wClV7IDwpLfCG6EoKQJcreMgxSc6EtUYxe3iEng5w5j5v2hdmLv6kFgX9GukGBYoa6yF
0oWlRi8Sauq2SHNDRWdSCzXS0Yu4UMXrE8CMfugY62Fxm04sy8MJ+p+S69b7Hoyz3rNo1OqK7VSz
e3XWbJMl4udfJF7pMF2V9TmUh42pDN2anDgV7F2m/mXdCDXI2IpW7YyPkdb99fCAdI6M+vqFJ/35
sXbaD/sxBtBRg4/nB1yHWtxKzqMNOesy+QP6U7PpccA6DySWY1dL24YzzV8z6WI8ZDqcQIPITl3b
e0H8eHJB6fTQw/OhbVHQ2zuwoa7PAzOgh7PuJzjPwAjy0vRKmKkAbMlx4iBnh0Z7DWgsmCTRbYWQ
9lVKWSCwGr/YG4PiXsAOaV47/xzLJPoQdJok7Exfd7aQi6KzpBlX8/0Du5lvkcU6LXYAkGrIdYnX
KwiScEF53+9mekDE7jMsLMK0MNGN8FX2Vtbp2NI0wr6nCovXc0mjn0783MMaCGDnavXBF23RdNhz
YBoaGC0h6C67lUDWnTZngCw06/UD+CTjpnXQMqY/uuNplJjoEsGG/08LF95eUvScsmjYavvQe6LD
6kyut4hNe4TOIpC7rxxEtj5I6gfqbKgpJZzGohWaLJOb0orq6EyXssFTBmC3gnMfOWqzKmeYdvvO
8OQxHsMWumtqED5ySU3ENZR39GRNDxC4kZ5D9btEKww/rkuf3AkFtbVrVtwHp6nOOjulacQ0GV21
Oee4EhAGAHPTKgrc5QsFjXE5Tim/XBlUmFOWvcB0Jzf02arH0LpEHSUy4uJY8yHrL7Ep4+UQRzFB
Fd/2F8nAVSITczNAN5HOSSnYC++Ylfj/EhF/XTiZsvzh3YlniWHXSYLKHOUUoRQOGU/nxs7BUkc2
xYPGEzUEZ0xHZMcHXbYPfw/dkRCfLHlx3/3v9wLgu6vUSyX5CNCy6mQiG6+r3U5XkUj+OZFWZGuN
GDw5H44GCZIo5H+2rK9jwD5L2kCZ4u/1RY8XeztPjLEvEoHt7sBksm1oSEdY2kZmsFP9/C0BWdBG
RxLPsr8wadYkcY2MSKTQn9TdU58809onGAxRK52x8xMzvgUeOVLbcA4bpFMjEvyZUdQJIwued1Wg
OS+kOGEf3pu9EnAVwF1QbuQTIOltHDkGqax99L/R3YGXJmFjru/aTV1sSS3GX3uilbHFqfxF9Tck
SJHhwicHjucrLhAkFEXRoDAln0Pr3XU23827OkhNjrXO7BGG3qg/BnTT8uLmHydseKDtW33BIuwZ
tDEDJ0V4IzZOqkfcUR529a5E4DwSuPdgOrbmPI3xPDcaUAjEsXOGk5nrIypRZIGavVWrXRZgeDYE
DJH2s/CTUiklBhXrimTMYMGXmM1F1PPhO5vwF7mxFeP1l4n1k8+FBaPN5CjAufVvIUAeh7sjjBgH
5JgZJpVuziCT1XJ2V8FMWaO9C4rR0g4KWEWYKctW+CApoZQElQslTfYxkzSNCdsqyZDDJUC5VkNH
fwaCElIubL8Pyo6uW8ytT6wvI4em//a3r3vhJWpB5R13ikN4Bi0KOuQtA+EPgvGzw3gCmuqAxdSW
mQNIMoNirqj4aEyOgjn+beGyx+Gno+prO72lgb8RU1H0d5NmDfVqMmo1mCPNUVAVN9FJEMzrgSkj
UhxhKf7itfzzoE90nuyUX/kKvMinJVF0I+5xyCZcbBSibcaghz9myzBehjpeuwOjA6PqI/CTvJN1
BBL3aviyBsuuGQEvQefsxE2yMYgIqKLb1dn8OCGZ5ougzBbT0afJ3xOEWxfJYweeHSuZUUEIa3lz
g9RUFZJxpGDJmfQIx2NQmCsYMd+UC+W8bEEwFdVe/r3IXECXscRE44neiy4xEQGg/r8wcSPxFfQi
H0ZXhF7ROh5GU7LVmza7nXE+81ESiXsdjIsN+Q/lLdrZbn/v2g2U2fWot+CwdeTv0JDRKmWdopx4
vKrZrgtDTMSaM12twPQMNgDMhmqZYWZYYsFzGjPXTHmPsSbboXyK9qZ2QCIgEPgCb1z7PaLA1urG
dPg9WE4BLY07CR0HdBvvVP1VrlKLKa01qTYl9SzwNOg9u6h3hbMPeGKoymuJV7pwu9ugV6tHXZK3
bW5En3OpwMtn3c4Uf/XK/Tl0P70xZbQZzjq97atlGjOT96Abp5wpq4IrvdA0CjeueIWWVEC2PIg+
SbIIOJydeVU6KNr3tRQVKYG6+3tk+HE3ORdoFLQzc5SHYUZGe2FKgQap+ZjtKE68n2+7E1EWS6kD
OBF7mepgVnL3/g8vVdDsmkiqmq8Qeeh7apMsZt9OgODOV3C9cjw+rM0t+xwKHoDJXaTe//jHm+yw
60pqojR29J6Ya50jJ+FfOKx79THWWRLL7W/zPfP845QqZV1lj/AmJRseSRgGdPXCGuz+noW8QxcS
qelovM6ALq8zAafwgJt2xHLYCOy8w4BORt+BkaGBdWPc87duedlNh3vF3bBfeZh/5jLB0nG9V3Fv
1sPdgicwrJUeIHlnBoFWJNpY1MxGFmBTwmQ97FUfgCgHC6JLwldCjXNyD2RGcNhNl3miCZbzxMEa
7mKoIqoFX95EKrZrKM79sGATJ7AVcqQqGWlYo9UgqLRJRZU2iZyvFQsuBCh+wEP8qSyp0Id1oiae
vtInIG1XVfFQf5Z4eevdpD4ABTothQNLkUpHxF8d3JIagMZcmGSBrG7tlBPCW3DCjo6O9ym2kOvY
C9cswu/S9LUdRtJYGIUqgdFzKFwwmY8ynMfdMaDRNd8Bh1+JkHvdR4J4gsOglQL+Fw+0bYe+W4pT
zMr/sZP8FubiOuG5Og8cFk7C1s3aQm7TK2jZYDnDrrIFgXH0IAADTIbigDP3DJtqRx7+BGFXaB1h
1623CaTnkWno8s0Kzb1+lbHmPRbbc4t0Sio1Jm6wcpBMNrZ0l2QN8s3Kcpor2YRybyEwqwityz7X
kmeeqxBhZFA7wMnWFUmiOswjTfCwUmLTLmpA2uVGtGz3SDmTSCueUS5gpQ9IkZHKb5W37wE30M0j
UpApoboIxSxFYJYltZjJ+/auOvMsEBtL2OQSLGQPw+AJgE4CbdGmU47M9VmU/RzfMtAf8Hekvzmg
giWLquCy4t+/REX7F83SLvgLIA9d51+N+Y2OoxZ8dpMFLhKsk4W02GBRQNIzbgRVR9LONHPlWoe/
zEAabocy+cn1zZnrBE940svBUUjUOL+RoT05sY/BJLsiCfTvV+L+Bi6hvjGft4P+X/jTxOyWINSS
ObiqJdo89vU76jxIdnkg9ouEVOgrVy4vtd3POYJZOhpSTOl6BSLrfAYTzBDeg8ddnrUS//z41lKC
I7maDMqFaUxCZz26Gl1RxHbSgdsO5Js/+vc+pjSPfCZd05AjH7GNSkp5d3TmP6fXnNv1rEkjSHOa
C3FQiZtioQby1GOWXZGWPHHVNxd0IYGm9F4TftwEKQMHj36vibI303icFltHi1X6khalvs5xi7Zi
Ysnr04TXynqDUZCMTTwxahgAqX9dVEG3dLNQO3rzdsDjuMRsFeSpFMGt0C70j6NZr3TmALH1eKUy
dEdqY2SD53Yr5qLJF5bvH269NSuttrytH66s9KnWh+GHEDnJAlVZ6zmeoCok7oBsG9JdQpp/MdqH
uM7FfK3x4BVZ9BgBMQMbAw4CbMPGlgQHjjutVDNl1b6EWZK3diWNiQs/DjqeTiqCuRZjT0saiqCm
dWoJpeeMWm/ymp3NNdRnm1eqj2hAnhr6ZC7+vRnTtfcvhdICUPlhNwWsJd1bZrr6V2mZkLQPqhmD
uCxWqdxwZ7yh7vTXUYphsAuBFcV1jZD/komLPrzf+eZWQ1pbSFxiuf3fa0FIcwZe4Smo5Muj7uFO
ApkJUGYSgihFraghISeSOOmyxN37Y378zzd7dej16vlc4iSSxNqfKED+RnZa7uRormh56HpKygEc
xBQsLO/mFRhxXS/6NkkFBh7oDFw4K0kb8lxFxbxou0bYhaHygPxgFgkeMxXBr+UCIbaHkfeZYzW6
oGHOSKHCjAqOZWmXWZYIHt7A+gno2Buvwx1SBv5MAy7xSXWt2YFI/R1HRigjc+guSpac/PEcOChV
lcCA954G8or6cAfZEWHlHXrXnFnNS6MPWmVmW8xRsBfU0Qe4GmUB+cqa7QC9jxsdiyzIjf75+e/U
+mYF1JDspup6DGukamsSYT3de6MW8I4yiF9osNkGI/sqebnB/yptSHsBKsVkxWF7/prHGeWNyXO1
KEq83j9o6mzrAW9xtdVxaL8+jhpJpyYBjHoL3wZ8nxwqnB3qo0+n7A2Ed8faPQpZb3C/ifazyJ2v
n/7Nk+F0h8accDtNhAUslgzj3CeLLrakotfoh6y+e3u/9X2rTbGlFtLndaYCrbMH08spyfZBiqC9
N/5z4vD5xpZAZpRjE5P/TZ9uXUqTr6/ETPnQWoPN06lv74Q3J6MTYEd2Kt/Zm2eZf8BER5ooQYbB
giPiEYfWaAYwfnxzTO+EPAdct39RwiH3BhgWUwySTWSXwpqvxhng1FZcn/dyQC48bI7wEuVvH/Pd
QSLuwc1JhUR+vwO5FYWkBEibRMIxpg7V9JfKNgJT0zdxBEJxeocsyb7SqkIwe+4VgKfvaHG/R2OT
NraldG5McDuK3f8muv3UOs0eoEbJvjdLCv3uWm7hoZzFl8c1YKfddmziWuC/owYEBSZsRiFkVmBq
ZBSonIi2VXhDhfDaPWkATT82GeSWODYErHj4k70OimHlxj4aKIw3uaOhtcoRn2f6+0seu+9yR5PJ
xv4930CSK/zOaqYua0up+UhfibDzYEeDV5tdu/D4dMMnuiO/jXT8zRt0HyVC94RcnjrAlD5qef5B
JdiIXcsAce4QdWelzLfSXuSFggazAtdGxFF/riZn7EMCIojUPytk7OxjU20Up+fI3iIrt1VUGyTU
CNRPUgyXmmWxVLIP2gh8gxwUVbQ9rcDkpjh8WaL6y+5SYcNT5ZA1u4uvYhVBgRbgyjbvCTG1wbRx
ToaSqFBqsvIN0ELcXZTqXABR+kxOY7BGKm9mnfjwwYeulVtCGMvuNUXyfnmx6XmsI8X0OwFQKUFm
EJFCPhvaw3syighuPX7jZMV65p53IWPTFTcaalmhcckSCXAQ1pv9qTxE7B7Ks0Xk5td0G3LiwJt2
LobwPWmJ6kmabnFgLwmYdhO1CupBEksyft17vzkGBJ6KeuGzdBCrc7i4ZHYE/KPBpO9aBPcmfnhA
0qKny7zfEkOT5DlR54YCHV+hJT5WvuUan+tCt8azi+HBzx0jQU7cfK5HaA6JPnqhtl5eHBCn8VDQ
/PFODf9tgrXUYP8xkfc8UHUD3hRqOikjQrD2xW6zgku4icobPPOGP/8VnYH9RnUZeTTKgKlG6VG1
GTRyB1JQwcqkCdznSHEdBYckLLE1clPnKtf4S+psp5iwrpexo+BUrTV4AbUm4jT3grPkvDGp21Xh
3rgrYYsQ8crb9NJc3yyMkQdwh42NLyvvLL769HTnHpETopvhg1rLHtYymelDAkfdbTtKBMR9GFR+
CshVYw3hJYRI/ua85+8yEojnUDo3fbF59HKW7o3n6tHwa2RQ1QYMFQK6gwD0GGBoMkKbeZrAg//q
vKxsxDDskbfq9izsC5gdfccpx1ibPYhbaO8SRDXg28vraoIXQDNI8+EEziAAFy2YYNAyWHCBWeW7
p/3N5eUT0HoT3QeFAzw4QZ46Yrqh/n4dxD4bGyvGvxRXoFe8limUCC8Mu88Zt6ERVbfdQBQhNIxh
HwXeQljh8gwvH0VBUO+544LYDXFH/+/b9Cu0eZLw4fvkjyH0PylQcVTX1ZIujnIwudcfrLxYJbU6
JbMCjkm+f1j2WCqNxJRFdlD36f60gZqafijFi5BddU/Vh3V1miVdJ6VcUdB2qgHxyJ7u4FUomhqN
OmAhXYZuhHIT0MwMdA4XGf7kmK5zYTg+JWdj1VC6seSt5+Tp3WH4SnUVvrJti+I5hKcQY8TgBLJG
Ff1c18e5rojVw6x0rXrQDIQ8A9rDBbvltenA83ByY/ptN4oRHK1jHflTOjG45RrvZCwnOF05UGct
HBSVWHgtJB7KkfkfCu13JpcTZZqmqnpLDE9Gw/Nq+cEmCJZVpNcUTg+lp2Rf0vSlLWUxAySzamI2
oppCZoG9pGRTwndV6D3BI1jDSIP0yMljFiZrt6WEbozlte9SbJXZdXwVwcaxqz5XTdG6XCf71Oy6
AEz0QQD4toeoEx+gQH32xtD3OKCC4HlsuzN7x4/nSkSar6gBVj+1YA9LKoIo4FAVwmWS58Ueb0ph
9+wxBzbx4B7mSkXVq9JQ+Wjbr+J8zAxqcy+yEbFpiUiej5cR+Ye+1moTMSNj0UccPLWnnuvd2qCC
RTj79UmXcyoBzIhiaEtGde035M4hcbvXqhDN9N73Vq3IAwtuxUumnDEqu8fMXMIyAw7fqj7jDMDi
ULUigQ9G+tdiVJn6muuFRpeHhr1+zanlvZjVxx7gCZJiuX6SwNmUVl5hplM4yVzClJg4Z1s/jRTJ
LWCuyFDh3KztxSTpJ2/5kZh1al+MJ6haLGiGwN4YYPMIsK09uLigNlyzgQbrObGawfyQX3iG5Ucg
/kt30nZy7mfV+V2Jmkit8CYVXjsH2pyjxybpDl9TAOMDA4BMSXfyjQS8cFctQH+m27XjMK+xvcYs
YczJQ7O2W/k9Icu2WC9wJr/5AcudOS2j2qjZUyhgdc0b824iTtel+BbyF6/yeWQrWmoCVTWw2TKk
ThM3NUUbhm4Xx6za+HEyqcDDNe5BG8DbQW35bVgR6UwDMZJ5qUsX94Gi4MlDCiiBAK9PAE8vGiqs
1qykGmQsLrlpIcyWI+UbXGFjXdoH9ZfIU5Cfe/ab4vpPsQ26rIqqIMGcteDS3XXFBpUfpa8thXiJ
949iFqOdAbaARQYe9/r096oBDzSDhfQCucxmDYy036NllsCN2kGUej1GSual0THMQGzzn33ZUf0B
FyPZfr9vX1+G8GyOnYn4+7fdenMJIYmaUvVLib6/BVUEDBU+D494dU+45RuXFctCLOMWlXdAbPFG
ygpu/dkxtpclWchHVofrNZZDie7xkc9Oz6vlOh4Kc5UcXtzXyrDvfhvXyrst9vRcEUx/qbhcVrY3
+k0anfufasguYkNICVQGNPncaD3liaOHicoutyVQb1Bjg1C4U0JZBMGep5ZbTip5/mMrjmRxJz+y
401uENAHwjSrzwe12mkI/QbwoXHJfjJBY6XK3jNN+hBQQ3x7et2PYYfLG/BRtsQohoU/jTPAbR5j
KwfTvwZGKSyXLhcAMPMHTVY7ipEIBoPZlYbihA5V+a2UYD6LU4kHhdk+jmiXXCvlIKV+0TbEoLDP
Xjm5WBc1WFzLi6ynPTojySRnUYG7HtvWcsuiTOKesimOSFOZL3SUYzkCE3gQuYa1YvxRr0pL1wdA
lDNWxgJ4+QXsqmH6Foyc5mfdUstKAhtv+KU5nNwc6VYYiDPJMGtJS+vF449OTuaASIN6l7iVCoag
Emh3UN92S6vTT+3I7BSRGyMUZ/iwiov42PRIWoKQP8vfSOQeg4i7Y4pDykQIDp4GEiVrCuxMWHdy
mf2w9s7VCS5YrIUlxD0WtpUSDBlKPATl3G/26SlbUBYah+O9LfEABRpVZySIHLM9pq5aSePvJw3s
g4Y2TCYjW5rH3GQGybZoREsxk785w6/uCsbOdsHVq/Qosnn8kA64f6Z5N9xz85KpI2JjxVSpBmFa
evVCV2MneI2rsd0wsqoxpmpUcwL29yh6doGfXt7yAhehSuBCaxlFUKYLszlLDoxUJv3nJmoXbsAF
3C6thtOb5VZJ/ck8oOOdrY+tc9BVF63tJKjRuXpcgmkrgUBOCCT+CiuF/5nesUlF7JBCCOj76g9Y
tdrKQX0UjVHmHeVdBIlaH0IgKGnFWMLKWBpmibc/JT+gmKvIW5FNG6kgDI5ssTV++7q/UiZd9t5u
hFYna4+A9ETITPTped93UwBtetrynVX5q19ccL/EXj86VVxzMxJHZY2qM6YAwKFvSrNvlFaU43GY
lCQpLbj2P4NFKuKTJ63jjZ5uudGIzK0tomD7crnzKtVh5FiFlHZetArthU8ite1rcdCq8KQ5H818
w0fPhJECebtM+8KWK6WFS0yEQcIpMHzimkyc//q+r6/sCybmZNEaqthcd2qUHFUC2DvRvEgvLBx0
7MmUR1raKMAZSdmOmruF67H5sR+3HeRiIwlTSJOv0oZsfPzczzV+jdz2S5j1CP6Rc8y/1HQdkfmW
7AYdsn6wXVk68l2BT33p4YoHg4xWQOHW3SPx2r8PdgoR3YRuY1hEnZ5rKw7QujcKaL5Dtr5R/7MU
7zji1HGilN0UQRKgdyjK+cbIONtdYftP2ZPM9kn9lGfTUQaTLPqCh/xcj1xJx8SsYeNcC2W/v6Df
n+SZcFG+XaTCrCuzMtGf6sP7lefhVyRXIACfpzEe6zNh/knLuB7ipmPzF7FiiEryAqAzD5zzzCRX
lP8n6rBObSh2oHlfqHUO7K52GgIzxavAQZRTcRgDAxpq8y38SgW4vi41CvXxS9+SILY78phElIEv
y5RVx9KKSbOXntZK7AApC00b3ZUuwDsZV+Rkoa2VWLBhOH58jGu5GXvXCWH8XlODl2FtlzKgEfPF
7kzI9oWjRyd+ZEWzNYfh+e2KNouM2bgLiK5kJp6mxaI1LL0B2fLwWGPXfpICnRdF/dDI3BOmrN/z
9oP2bBZwqkub6EhgUnbiQVruGULEXQcp98DE3fJVyfcg6VtXsiCRlVweDvG4bappvCbR2ZZV0qeS
v3XHJvHvSQA40t3P3VCdlaCIntuXopNcXIB3Alwhh6T0KJ/xUIYgfAcOp0YZgJu4lGSqv231hJms
qLWsI912CUu5Wx4XR5TeR8M+awEfyOPV0+/qxFe7xroosxvArXEye3pqesPdvU1vd8hFbmL0I/Zg
m+BTWs15XPl6lylfv4PZe0lNDx9EDmGpljkuGau+maYkTrvH7iuLVqLkcXrVQH8lq5D7sxKwKVJ/
Iu7WIo9kz+963kYiUvcG9v19TyuR4Xysd+Q39q5jbTYqhpnqyws+cYcE77bZDpfB/KABPnlxnUas
cuGc168I1E2RfZ63dM5FwOBTVomrcFTY9kWJkvavxA3nROoijNtfvUsqwS3bSC1BDpWR5AY+S01C
2HU8F9GTgecDPZLqMDFcLIu/0ZvupfvBvRn5xtAVb2W/wxEKlB8VISC3cq/h4nxUshbECbXyyw09
qATiMwjAD3btbwuJc+uOG1qWkZMr5qi65PUBvqEQohnAFIJ3YcjLPgv1KypnkLLDebjKGovbs7Sf
FW4S+n0TCkyHhLZCfL4EhwLa+Skxa/2STacVckYnHNrRKSKlEQbvVVKCWf79jmo8pFpEp+MT8iax
bMovqL8mIDLy3H9MPI+kHZ7nLn6xthvjI/o7MyWmkK8t1Mh67JzIqTGHeVZeBc+zb/YxdbosqHTy
2rWUr3iOER73n0OSIj1x4wvMK8QHhj0lbyOtKtA7wC34+VSCyikQ2a3s9pS2MEhGML8elSADFraW
JvpMpFaXQzOJtMjbFiuFE990TU+gYAKrcNoOsdFoN25O25D93GzkRB7/t70c/zAeEJjTsphmo6ah
z9T8wgxPbg3CmWcUmRXz7E45BCTvt0IaB8i4pZSi+2PGLORnvf4Al70mRgkbUPb3gB/rTNsBT7Gf
I7112siM4H5Mostg2Eas7rH1POrDwB7kjCY9trw3RUrsylfbDtE34XHNFahYMzu2YI8dMNsrlgZd
GZtrU5QO9zAHq9qxBSntMZlYGXoMStmawOWaaymJ+jh3uvkw34Fmi0FQ+9P8k2dfgmSHy0EJnFA7
89o4mIjUJ2priM6wzd626oLydNZBHSog7faQCTpywutARu/3Koi/taLiRCB1H8rl7bzqzTkuGDzM
y3R/7hhjDHEunJN/GQR3VFbyeRYIBeeP6oJCheRmYXu5L9kKIvtM4dTUemsPsH169mvBzuZWRp1H
F3IRBZ/FCiY4g/ltme9eHsPinhL6BRSI+iRmdW/z82SA3NdoE76Zp+5iu9g6HRRIXQV3ZgAdf8NQ
x7vM5V8Fe7gfQPh5pJW9iC8y0nGingGh9q0/9XU+famvTKlXTEKz96ZNWM0IaYADri7zpwwrVYIR
sNTkxFsHYHfGFDDAzTPBoLv7a66yVel9RM9iX3TBzh7qQAWVGoLYb0wmH15mWozkIomZ/smsu06S
8PoUlZmMe+4Kc9WiO9Jzw6OUri2BTEm9jgoPMXJ6vyiZjV0tLndt3T9K62JUxYhZGc+JhdP8Tr0w
PwrMucc0kQl41ayo0h+VC5Q5NvRrbraeX86dmP1iHSEcZgM2QpT8eTUxP98gp2ja6fZaysG7p12O
Ne/BdJHm1EZPQ6LJeC4+Jf+puaYHwiEzi8cW1DjfsiroULmxV8jVcbEg0Rocijq71wg9SzJ9aSl7
8sQbpfhrHckcvSKUocfzz7oCcR1mBWHCusaOqwpoQztMMhfYqJXvuJ9Ai/kgF2pIwg5aQ+iRNNAU
kvLR/vm4FTAXEMt7555ByBjVw+nmXllrtJcBuKOirDs00TnrIv8LkS9SF/SURWATyHr0X2T4Ryvr
RK0cZEo+L5uQmrKK7iP2t6rgHsUPvPzZkRHzCJMQ48b3Rwso9R/dhXPeRuGzfcK6MHaKEE/DJc2R
MF2z2wpQv3Nz+8TQmmyXBT1IdTPx6p3wdtrSf1nsswRulGiZ/IPFOoW0NmCXMs/Tvh2SbK1ruzRe
GwxHtO9lMFRPkJdzInQbph7Mip/mjHsPv8jD37EsALIP/1D4pKKJxPnIselvFvA3slVIqxt8//QT
wvedwF0od4lopUQAXzSx22uc9wADpsOcURILxKvOTa3bf92mobCFdUPG/TJYQWfgkNlquEYx8fSW
QRwE3FGL71KZD90y4pdSe77VKmsD1x03VYkTi1hUBHRmPctX8/RFidqUp4Z1TAZaeEKVvpqVMl5X
ZNiUaRvNUErZDOLKoNsJbJQDuwH1fFX5jj0qRYKmmAi6tB4aGg6NuP+xrpvq76j7BAenrFJisHPQ
HJgrKHA9Lx6TzMgggkaNAQl7xPhR2oqt94bU3MLxu4K38AJYdUeviKqTkqMJZ0cBfgNPgNUv/MtG
ZMOlLiYFGZXA9gXY7QduE+hIwhbdsMgX4y6VWeFyW4ysIbMt1qCeks3PgtCNUsopv/JFQRFvrI8H
+6jYadRzilLbLaiPeIjSax1ZpWcWTsf08Lgr/QGKnqJnQUXQDyCsueRZwIvng/y1JQBhbeuqLQ4I
iPhDq+0XkR18/eJnqPhWMyD5IaRcwRzQNTLqzPXwESX+W7xiD9ib3aP828tDnOqhvz2kQHqzLndQ
yk/pJ89dd3RK+Ox017KS/yu+NZL+3I6v7E+8vklAeyXYBhotMiZ9DSu1BrOUWe97uyClrzeYVvHv
g8SFTh9yTGadm/q5WtKbs/5E0ClwRbXjoEJS2v0TckHvn0S3plv8GNvQ4ssvv01LonDjrsEZFS4c
Ccy0MYSvhQw7nhxZC7a/pg8xdAmr2VdRwqHpaADqezf4b1qjdB6/DeVBVJ5Zj3Yl99MLSUddW2iX
2APyWOhrW4uiWCAWsv9GnwZnjHsiTvvLmu/W3UHUU1L+crDpB3hoG6gqsbsMGVF0wGwqPHhdmRMo
+QJSI38Jg4X8e1+JrbDFShlObNZhunLARuXQLZsUfVIbuqnJ9bJUwVtwc3m+wOI9vU5YNrvzOka3
p6evqqTTk+mUulXjlCQ3s6bPgovDDA4lJoQyqDRJa4yotJ44YJuV5Hx/B9dP5U0LrAWfAOJoszZ4
B3wMZKN/GsuvhIJFa0G+hYfDAsqQTVesx5Tsim4dU1lYpt+DZE89gDzr9JCVORO5qiflus8MLZxm
/i2AXz7w6OKQHKXhcyjCqWUKPAqA17MLhJYmfuz1ypkNJrvvoBdhpPpf6O1Wke5O+aDBIdj7XW3G
Ng+B8X0b/Ic5lDioXHb3Ya2EM0Wk5XlvGgzxXVNZfXj6aklC5EGuPlajsvtnUmPwimpLe5ukp+nR
4TDe3zGRNRTwpdJdSQUm0ZRqB7MqzazY4SdJi/QosA2BkpCbsMHpUVhhRxIumAo/kM7v3ig/Q4QG
GUki2WFPYicyOxrfP+K8Zl4XdxXFtN/ID5RCuy0effGHgFx4yUIn3uC+EyRFl6dfs67g1jNvcDyh
acg6GkVANKnjTHHW8+U42c1SlJVw623h1GNevb3/sKwDUB03N/oW1V0StC4WAVW1OQ+8gqOugrQ1
VU652Q7CE52ThEJP/8Go3f1DG1a2bV+KwjAZYVaK50RdjLG9CHvOheHE4euvPcX0fXNuENbIDxIE
vrsr8hn/KZlhx3iHAN/bnmu2zcmaMQqXId+CK6T3NecZEm1gsue4iuwhtLmanhSErZnAM5fsOBbD
cQzKLntQv6BpGfGQGZGkL9SicLPYaYTfMKWQXImuSYav/M8+dO4dcJDOMGRn8wsXYMucPrgC+3tt
qg2dWapTsnIm1Y/J99m6mtrElxHTOQ7cpQ1/klsZz5+w3Vymv1x11FKhXwAav+hw6P+0lR5zEFPs
250zsmEjuEmulwLLvBh3C2+V/hVUOzkCOZowydHcqc3FFs6KryGHzsF6cUesEcPWmqkX2uVpkOHr
9QqUbkyC8rAslC9+m8GDNiIIRsQZSxG5wDcUvVwr4bcjWPdJxDdIgAiWPvnRWSN9HRHj1CFyYeRQ
g2zjtcuxz7+vNMbdbcfrcjlZGViSlbcSeIOYtlhOSWf2GqmP6UBSCqsCphoTWUeBddLRoh4c3ap5
Sl8j9rNuo/TJY1009emAKb5YDURm1iyaQSb62JveBkGK+JlU3ppaYSAom0h2pVEGnPLAvH5tmXMQ
Ga1YDGgSxrWHnweB7mZvvtStRkbMrte8x9zDRRc7fSmlbotzIMnQ07yMLoYHBIxtDz05qZHx1fGi
vM/PyCwF/GnboOx2Wn4ACkuqKqlZT47BFkN8dCVdepu09NBJlwfwlW95RICutOfFw8k+BvEkrHjk
/9c1qferQPMOpTEHKsRiF5XAPW4Awq5g6HCqqN8cTwsa/ePdfkkhSQISGKmQTFH+E/+6mo4yFFpv
A7XbzlOeG3hgg00e8SZSCXHaOmvm7mzkM5IqUgRrdnk+94LaVhSzxTnT+4V3B8hZobFjFq84TS/t
E0BFPtFBE7eKLHG8hdw8d0MljJg2y+qLfP0SqQ7ltyTRPVKHtDSn6Ik2QHa9F0xZXwDyR38IgzJX
jti1W+A0P8OQwujpz7dgNXlhrurSvGDtEIy6jQk7nr06m8aOSBPC24s4vZ+3gNP6HYvRHWc60z2B
PoIo+ZHe6RLyFcW1sF7CkBGcWmFdEhiC5/OjHt5WkzLR5uD8R+ui0XxFLyUMsPz+122HqRpnl+9d
PB4o4WqQ28RhoTukzQWfFU6oa+EIgrqrVH0/nV4+YUlot+hxS+oQ9FMR4SVk9ekYGqVjZxqUbumw
VwhsZ5FTEUvUzHncczfDupHui1x5iAYBLZUy/tKsqUolpzgx7LepB5bVIm3d7cIl8FciG2QkLISU
s6cvayWo4o2+RW9vbz6yLeOuHVVmpBjZwRFi8w9SidbQ5PfWuuwq45qg+67pfDV71DE2c5OWPWp+
aYwogBabwpSGPKZ/vv2yF/0V0M4RiiaSXLYq+PsvMeGZD+5ZpzcBTlnpTA3Eqrha7TvRfvj+dTWz
1nZVgupOOMwQ4wLr5lQfE8kxdEXc/bYdTS3AXjd+Lyek4z2NJ/xXhrFRBG3LOwJNpWDAx4v2TOss
jksoYxN+gpderV5YP9QWoUIWYx4OcKlojYg25n7aBhVANJ8xzum1zanw6ux33dn01vD91WeJIh23
4KnWKMaBcNEJqq9YNP2Dft25fp3MnLwf7NRG3FMamnsKSgdna6WcriLvkBIeNcYxII57nolxlrV7
OISFQ0k7HlHv1QoKH/machN7BG/FuqhdpRKNWzINBEQRGE0H6tzTWnQk9eHJWSURRomJfVY2TuU2
97CMFPPaJ5E2h4AAtwVKNP85PpZl3wKbkr5s6kidBPpv9XLYVEH2x7iljto/7hOjlXGloQzTo45p
5Rk6fA3zJEfTLZzzgyUtrXEZhMmZ7j+MWgh/QdpteqIvNulq3IvkwvMZHGnbmQaqfORLnbKBMkwl
rLKuYMXPlUOer+ySh3iwhBtwMNKG6W2qidlpz/nezSeIV3LgBdMbCpIP2HgkFhdsSFNlDHhf2M0D
DKNRChKnsb7Incz+ZkYWT3wHMdDi9kFSO5PzK89RZDL/PXNPbemMoSygSIrhspALu0OY9p6zywOc
y/9WqQRdsY1lhf2Zth6CzAAAy5tLkZqQ6FRQre4DHcYqFXE7DbmWTwC8YChqAAl1AR+dV3WE87O2
PAYhZQiJbCKvcVUnY0W5XfOkry6y82sYYa8Cf0z8AKS3y7RvKoYKcMfoKG8Ej0tDKvCwx1GqDFG7
OdgV+t8yCLm5nocRYj4vLy2fH4r8ffGLoYJ0wVGpFqEg5Z/enO+ioMkl3O0zf+CgjMQQDP1TR/U1
iq/16VNadrm0GAWGMneZNtUgkmL2FujMFmO/2wEUI03NU/4V8hsvvmdftpHDzFs32+8jfrz1X4TL
Fh7xVQZrEQ9fXmQn2Rts946yPQ/9FvMBatrEeVVTWVpjaNC2HlHJllTCOpwdHtlovpE9TOk02eup
dyNgPkpvXRynw2kVfhoLpJAPoJOICHxCsQL5pBEkNxZ4JxdAS0MsD4wo8YK8b+tvYiVZOg5ad1cA
mWDdBKN5Cu0iysAXgNT80ILPVj2zF4sOO3sMRZp7PvxUpwwn+nbm9YSbtyzfBqBYMCqvPTQUYneJ
1/EUiHY025qU20p/Bft+JA/yjE+Wvqht52/D7pIV93F5PPpcq0eQ9Wip7xNlkZRb7LPN7NZTgUO3
qePmVFi/8nUvEWmky0vtz1LtaQ5ptClXIoYFrSpYxNceiL9itZtvPbjofC+p+nhtvE3mkX2vST4h
6T9/fNyX1P296AxaALAkz9ItFhcsQQB/lzbDuoIQzQ8hR24fG9JZmbX339iso6ClHJrbvevj17lf
S60jK2dDU6LBrMtPqlhHR6NJxuf7I5kZXk+1YPm7bCIOft2fXww/eKR60Zuv+jVHtGykAV3W0VZl
r2K+j2wwuKopIPS8aK6lTQy+jqrN9MMPi7Q/KgNajlX5z0sOlzY+mscd8m02Ym9DnXpnmW7P5+aV
p/CO+S8l9sZZ2KiET/5Fi7/daeAqFEcIUnLbecl/17pUYSvAlvCrusaCg9H2f5PJAFgN566WGQ24
HvvGBeXNd/jVYSaqzexTsdTvm/k3uA8z2jLju+Z9olBo5b5L3XsTyeHj9vt73VpEQ6j0G5Scj1SW
pZTJNqi3MG695S3h9BSsj9aDmEHi/jra1KHEwtgLAXqFB00hoh8tEyRuYNQpJs+LxDUQRBpzFupR
dXArja1vqCDkvJ7hdhjCYjA6vkT0MqTqAMdPihe+PldbNlPEXV6qQzFK1iljrOrOXpFyKvtgRDqD
8y1VWjDeezKYC+rUhwHnZj0kQiJJ9OSSovEWqGwmcrMz/r/dcy7SpSWa6rJrtDeVyOJ0cBtmKe8p
9khp/sc1/7etRMBqKAwhnw/NOaemRsH0yoyXmEHal1ClH+O4QeTd62nTvnd51HH10b+11LKWLxa5
S+v2bddKnw04x9c/kXr8kHHvmMjTOy3rf5q3dD7H+DJIidQN2pIqGk50d2+u+gTW78aM+QHPlqYn
s4dHUI+PC2Pm8U1+TPjzNpqqYdtKHhmGxNSu58rHik/R3/36xYjJ9yZBKRmMFwN+xOjWUXY3ObrK
rD2cCxmF5qIEpm3tXmcEIwinD8ojq9+Qrp2S9A3BNLVTio3huA2fOQtJF9rB3p7hA9vf9jW0Wfbk
Ge6vT7hrNY9KGjUITVecuSSJpEpaaOrSZUKMrVnICHJXJyUPoZWykr19trxtfnC+6G1ZNdWoQhef
ETk0DROe/n60ZScb2MUQKB76NhXihE9ONAvb0kzIpYGJfci3hN4pz7LXZoTtVwEOoGfQlpeoYlIP
Ae+1ZLoUDgXKmYgzFWXt68x3coMr2XR1ac8M1eFzwyn9KQC/ZxMoT9XjXia6WLkECkSc7F5mfVE6
NdAHrfRQMD7h+ExWfVXRH2O7TOVgeiHQQxz2Za6vJ5OZE15GQ6x0V8gO8m4Z2c1K5raK3A05MSiQ
jc3oj+N8LMPFzTg3ZDfu7NAejcRrc/sBLac1/QPcPtAyc5PbPP6DaJBesy7UEHfbsOI2VQgNnH4z
SHKR0ENwUoOY7W9otnV+JPa9ydVyjeCNRj64CJ/m0ve4/pRJiX7otTS8GF5K+jHWIrEnfID1bV17
0WAf5BFVHHosXC237VfDUWm0WoGdqegmbCU3ETn5eolIrtps0vcCAfpZj3WLQmUk5czxoKs/LU86
Sv8qcStjpfk8GbE/vW4lbAAGwqlUMNshlY6d/elTPVwyjVDKY4uD2bSoUY/jBX5oYo53L7zYpgv8
YNuQ8v+TxuJhhVxixkcha0j6rhvGwn601tEP+pKkELdHrktQZoLDY1pIBh4d0FzP6KcaRgD/v8nt
Nm+6GH7dQniFiaRi2bfROML9k3fGN+0XVGLYjuvyVg9y3Pj6hmzJPpbM4We3syXW4PoeXOiGJRtx
aQ9wcFi4WeG958GKgFrDXmBo7poeSfLiD1pi2fQQTNHZE8J3HYQPtpRVxbtSGLbeJy6IE5cLlzOi
V6QqRPELMQo8UOaLwO/Y9VzN2cJRS2zwbk26iCwv/tNZa//FZtPe8Agi2mGYScUIL5OZUK0ZhBHd
9TIBAXK9g5N8Gw6f5CrTEkM79W0LAYsSZn15fudItlH3BkfTPR4ObxztYNBQmyrIrXreCuwbN2oU
TNbuleDD3ftzc/sT/Wj+BDKck+anjXqsCgom3YMbuWiaYSEZecq9Bd10mcGc1WsJ5GssBovP0WYi
rOljFpabu9KC576I1zUWWaj/QJrMiZLE3AiA3GVcoqOfIL8V+xZamLD0eTXX1sJGC7RhKJD5QqNI
C1MY8q+KYwUztKItw6FZgtQ6iWAVOpZqsxBNtIUVyF0QcYq08i1KpgJ5y++/QpSfVrVKMgF9efgl
qE2ELDLki7Ieka37KG3+jwSAdZNsUzkDuFY8xx0X2yWxlm9o1gpiFlxMoIE4cK77y9YItHjR28+C
f0U/p+YfIrTkN0qLcyvkquqi29mEeL91SOmwRVTXyH99BbfjqJubESR9oii0KMV4QJurwrEz9Z6F
knzYd0eOYKS2aCuOvmcheoGPALBsLTAs7UTyca+MrUhkH5Gt85rNG0PIrtfNmCv2WIEuAIsCHNUR
VtCYZuaePcmINRoJSnR1Jea9bmdvEvT8EQxuC2lC093jPcx2kb7qFgBPxPJDRiVA7SvCkDTjghgH
J82u3XtaULE6BvniEfI3WQ6EDAh/pq/WddWxoJg80UA4gg1PiUA1E9NpH218VqyJgMoPm2QlxD4o
5/BlhNLAAPO1vZeXXieYVec3JKkH25wazFRhQAtfhoeftoYTp0wAEk7wIp55qO4M0ZyeowSYZunO
SLQz25brPpHc/NLits9zu/vLRqLpG+ktcnbFQz0eTIfCPRBczBncm8SpD8NsqzKbY1G6k5pO8oIg
IfqVFOdYpKjkJ57Ujw1uEq0KuxT3bMLXosYHhy/Ne7X6gAGbp5XCzrzrfb6/Rbth9uI1JWNZn2Ml
P6upyY0Z9YW74W7/ToyEnGhihJQhngIBwJX70E+gm5G9GKjv/w0dd8xkdH7Y/h7L+RHIIs/ip28w
SC0FDLm1uA/PXN6Xc9w+5gigv97M8LYLtMHzd3FAqW01DVPQHm7GCQ+yBFaqRQzXTYg7MiH7Euur
WmaJNjEiu9wOn3Hg2NEOOWZagGT5ujtdT1GW05Bv3K5wSwgLhNm3JGsLRjd7j41tuJibZBPNhh1z
DjwfqJ4UiFx621OCA/w+m4CjlgOCw8FWNi2PaBhgtUJG+onng4lV+0rRS6a65VY5wcr+shW66uaG
3w15aAPhiCxfh9ZMhBnWcwWdAbRFh4EGXPrhGWuceUA3VXtBfeuV5JKl1q9G3k0SvnlOtvLNwoYe
X6DEPf6iiSjWH/MHQsUP8dRiK+RTHTkZemJlysaKYoPoPDER9Ft+gpcTNt4oPImKGH7apliEAOqG
2PgjYi+y2+8Pp617prvbEHe3mlQ7wd3osCw6WPu6Aa6L2x+Nhtx9eMCRxjOeoaeFPRGSuX6pQW8Y
PoQwubHR85OqIuVB67bMNZrs8UDKClJosKHz4w+RZ6tprUPijQuZgK6I0mOxHzm+YUSoNmPR30QU
TCxqPmbLUT5DNKkzZQUxiQjDYFZUB/fPaFYCg/W/qTMAsUUjc61cv3EfM8+uGZR20sh8zy5i9DO8
mrfE6dm0OQDCFXb77t14ntmH8LCyL/fKLSD4MAJ8ITO5/d14xb5VpVFHN/sgLfyAhXT6veWHLKxo
AS1CCLPjbcHKC17xF1RTTCNQwt1TJ3/KSwIX6eURntOszA85hIiziNcnHP47HKBjTZbU4mSNc2fB
xIXULnj85Qa2QvkYqhUu/fEr0ONNYUFGcRKRNTZ/ExbfZdx2WDvaftSHSGHt/CfbSHSduZ0+v0NS
F1ZOsaCt+X0YCPgo0QMqjUtiJLUd73fiw+gK6amtm285MDHVxAWIA6Du3DFtGJPTORmMEACqt9rQ
1+4cr+FQD3RweU7TKH/VPJFsXuO1MMMGWNMnxHIErU5PNOCY7TdffzKWV9T/lSPlykcUGfz1Grqf
3c7Erc5YjsOU/mlemeqwiU3J+7exw+cHXBaS8GcSRQ4oZa4M84lOVhw7wQTGrY2v0mg2WxPd50q1
MbuLfEV9FeBxkZwh7WWOEZ2Ag/JZH+rWQOwmMb+yClYgc/7kAL60NrW4TOdyUYK5ZyfN4oQczXZG
bW11pikdeW29k54w7EE/Yy3UokBjqMFNWBZh3v58K3dQsfilDSkSEoZIYZdXW2OpoGgJGcZJaEZ8
rESKLmLUIhA3ZH9pLTu6BlTlcmqUUHJRLxI1ehnRQQREj1U1bVFFsYV2y9GV3uAGHFjFV8qIipxU
MKmwmEetfu3gjulys1laMzbt5Ug7gUSJXwtMF6rKj3sx/lVJqbiw38q67mRQGI/V/fVupTd4DoJo
cqObKRf736QiGfF3EeRxZt/KSRIhX9R/pq8dwL8FdllYGC1graf7pXVROh9tSFbNZUVbTsRAmsKe
JZdWS8PBmtkmB4CYwcICgiBCGsE9D5+eRx6RoK6TE3HemEaSud14dZpvXdTTo0ivq0iwLB4tTev7
mwuLHBBcE3kWsNxhWhlBSPCjKTZD+1C+uFrU+bk0BDAIW1mLIfIr9rYONbNN9hfrh6LsgJmjR1uR
nCoph/VxtoBBmTv0MtkSMpXVRKTBSqqhFVAITofBoOdZwvVF4G/zjCucc5vZE+npsKYEoRyLe4kc
UY51FWp52p9IBlAGeKUjumOmi8rOaSN8RmfGf7dCVVi3pNXhLOG3riORrYPNw5iSincAWQpCHYXu
y+3e4DWyAXY8+wtNQr19aNm8jr2AurAySHicQeeGQ37mCo8KCxD2iUgvWGHgtsjkfbeZPeshNZmy
ATL6828Xlqb71Wt98F3a8LkWMhn4La6A6d7t5VLTCNGdpXKiQgO1VLwZjysndKs2cjRG94zy2mIk
4E6rd2WQzJHwpi63pUMZR4F+PR0qxfxmIwJNgOtWlhxIBMCLAGluhexzOIo89GJrRpcUZJnMLuGr
+RJJDQVKJ+3bpStucqnTfPyV/7JqXAB7rD09HALhrZbwmE9vVXcS8N2DwzeNY0mz8N6up6PpZ8oR
jVaJjq3ZIREYXUYolHMTIK+5qG6TsHA7gRjD6KpVWn9U4GZYEbOSETVwQASVelysg1LdpSxiT+x5
1W8ZdLQITPFxKqnk98cTtgAf5aPbGj3Ay+uyWrNpZLUQROQ3ksE8FkIblpuieOQ+aF+0F7sWaTCY
U1tBQRcM9N/6bDnyzCkZG8Of67fBDuuOIcrb3N4sCBvmZX+6I1mLpG7GAMXM0h7zrUn+FQU+aG27
HwjRvie8Aht8MT8MPIkqHSrTqdboaUrjVUkZYkpfMGOSRoq7vAtovqvK9GuYfI2JqpWC4+DFELy+
+Eeykhj0haktN/2+gyqP6W5DdJ2tWc07bkveE4raHDSKbWinzpwkjcYRMKjZ8f4zjnHVvEiMUoh4
Fy3UlTvVbZpuaHe4O1RsBcFKSbu2ndQJx6cvVMi+vZWm4INfzbBr5OdEDI/weGI8nQEdIgZLq4WI
816SduVokdiTCXrHrmw2epzLWJYWbcuyfi7EnWNcaTN58k/GyLx+R2FmRtpzOl/OHlxnePIQQp1m
SoGylOzWn7VQUg9zkici5DY9O+flipAudi7HkS0XM1dP0HlLNq9Al70nhFER0qxXkfOH33AyOtMx
Lprzzz72zr6GmzK2Lcy8oA+0pUbZ5E2u4+MBvi48tz/IfD7NtaSUPGPW4oUgBTCIH+JMKE3s4zpN
iJ3X6BhYkTY4B2hcWWQMpXCtzIyTRYYEYDqngNzHpn1ZpgMc2EELiRwANOJHWjAJvivwCUytkuqZ
dpHRytsfYkgqi/92JC0LQ9idQQX9fQlupVzvkYhoXietGcQPUQjuJR+6vHFr4ta4bI6N1a48xUMZ
GcEcKCpJuX1gjuZpV+WepM6CYkrhzfthlBBh9DO/wFttMu/6DnoeE6jlanShOJxu/cgL8nWOQQFL
0+cuCUBkjvvvhO+LdIB/um1MscSJeIpWfrJHsWbs3/3nocsaJlXBZiTSyKefDKd+AYP6recZ9NFU
nnvoIT7yayQoOwVD2PXCz/atATsBuUkCl/T+baGAwnSSrH0AtAz29Mb/iOcvNeTJ9v9EmIbskxHP
MiVWZrJCGZvKKiIzhS5UMRsjndZHAgdeQj+4pfQkPK5Bjy1wER+1Dd6wr65Yf/fsoRwCDqwa8QNk
PVwF8dunhqLt+VgbnrgjygLf3YQFOsbZHpQFyWT9u+cF0XrTn4PNkNt57tWDR8JZmxS4dtaqBuQr
IngMal8IbBzNmt9REyhaZU8fw9Y2Ggn9nCLbPCTz9D3rSdKt0VuO3fNlCcU9zqOQTCRaRvQRMrSm
qt9IZMFaM+zu/vOwSEw9DvqfoTrowzz2kDaTYt1skXKAKWvqHf076M0pVHcuvq0i3DJZepDeHhos
/0FSA9Q9BHj7kq63BsJsNeh4mzXAgAa+RpSagM3ss6BaeSqHI6Ph9FcT/BRmGb29qAtpBT87uFVK
N6OnUe5d20qCskTL5JvVgOl07VB+2STMDR3EGBcBpe5WnKhaRPSrlmg9AJIE5/lX4AL/JU3cFA48
uEls4ZOrSgBy+JsTl7x2t7KS96t5hzK9xhAAqx1INW3OzE6Ks8gj3hNhlBG2u7xDkUGDlZLeqOjW
MxP3MTOrkWFfjfPMEEcYiAdy7LUBb6LrW0O6VMuu/xugJCSNsH/gmXstDz/RvVpmGCIKHCmnuqU2
7s7X7xBPilyyxKuysp/2kjnCkBDV+dNBsvQZb01TwB4AheptTxRzvQpbo8JyQA2gI/9VFWfXNxxs
ZPnzp1gfwog9k1CAusy3oTFbpb/clScceTGzO22chGkAY/JBK1+JLyEQP1Tzyto7L0luHH32YrX0
xigAWjkgLyKIqAnMMsdTiTqOtKx41tfWDeBZMbCKVc0vyuIABxkANeTxyxdc2ZGb4432YMc2yp8p
2opktHeBHSiR+wLq3hwCB2dEL/ZWLfSGwzaaYKi1Uw4miSzrFQ0QS7dC+ejzkOUyHsqctV4j2JhY
suxcIyjU6Zq5xYaNFpNqAmSRpX+Tsf26n4uoZTcK4SSE0uQkcxPA78QJggR1hoH6rJYH4lD/yz0h
fpY6F5J/LjuGB2yxTvqHyL1XI1FaINCAyKqtOIT7yjWeP3fkm6ylrmfOovuNVH22kkYzxgSkjRGs
z1szpEHrAJOUh0pCg8gBl+dwoAIWcQeRZkg762rZYtBv0qifMRdmfbe4t/4KM9m8FmFQaEWx/ai2
OWKzKvzS/Hwlbd/LcVNUA0fCKdmLSbg6J24cffBdVsA4mBVfthv31ETWtco8YX+YfMrcXAWQgcvg
TLyDn/UkrFe6O69o00VxaMA6N8cdKPgPojhQKIv15A434aHw5S9AFUClgRLrTnsOFSITUrmyitmC
mP/EzXn42xm9fh3DKvQdGoGMZFea4q1Zl2lX2j99hoLYnevxv1VMfdo/aRBgc6RJMjh21gqS/sfY
kLcGMf7PF8tMd71yyzqJKJaN+zokCWRwVQwKwvcohD65WoKqFsXZ9qANyvLuS4Vw6TNN+/4YpUV5
rANvtJVWCaeGhlRbjaaPstx5FZ66o5KFYWM+89StbNYzVCGPB957YM1eGVVF4pi+H4iykxL920OY
ThXorMQww9vUfeJLO66Hh1pWAnfad3I8KcVO8yT61kRfJD1wYQupqAR8PZPaNHUKun7gWWb41EI9
jpl9dm8HRiryAlHeS7/FCUFFQ1brAIPCOL/xvsjqbCM18lhhkjvWmIrFsRwHGP7GPNrLXg3zg62D
ZBaEZ0rZOCstXm7Se/id3eK74urGBQrmK3qoDJ3QyzPrbDlbBkzWHaObiA3BzFkADdBhQAYhq2VY
/yMWtnhEaknK5MeXJ49gck2TbKWbIZC7iimBx27eJ+nlCDg28HMtTNwnbuxVfAI2Tr627B6+cFI6
1HOXXxlGOe1zd61YIusigoKqBpjzVMHofx5G2krTY3kyy6oCNwjmfV7JECSMrsJV4QB8dSUwIory
6bMKsU7ZYfrkGjRKGZvBnQOmFmuB4ubjD6iFpdY11BBy3lP1xCSzRXkpuRBDT923evIbbXb1IfUq
m3CDhSEK6tcqwu26iH3pwlV7tX+O53+0rcMXsCOyAQu9MI2Cb66tZGo2m2loFeyIutBrbqPGOAoe
31i6TISTECQe6JUoLQZzWBB1tIjP/XTELePlN2ebZUqMruXRdaeZoR3+bxz74OTsLuvwsnTSQRhj
5slkK/Zd128QH24p0UgGqibb/hkvD96SSaRkJnUycwnucSQAAC9okcKhpnmqbCozoeRw+sJh58j7
e+Jfcp/K6JDS/U38b6dXaAyV9d2RgADDQKa0QekPx5/lVJbZQBx/9S5pb2YBO8ClD+g3Q9/S11EL
m2PwCZAVQzZJketXl+KSZwoeVtVh53SdqWeG4u6zTMNDpas+thvyWmv3F1kbPUkUm4emp/3ZSt8h
dfMnhtnKFnu1poL4vDU6VwuJXX3MIn8adzOgCzTTvv3cKMWsz3QkAd7xCIqL7i/eYNunK81qPIUE
0e6vph4Rj5rOyYn70v393FrbzSQFdUevwVWES609py66jmuGZXq32Nz6hzulJzX3BVpRyX8APmOC
RkkDGIbpkf3Fuzv5fAMVnpQB8l3cOggjNbLRh0Z6HYhYa7aiuGa0+7MQLYsmxQTSV2iSz3tazVxz
ehV6rvwjGKWVSgs9VUePxnPYO+VxifSYHNWHy8Rc8b1W7eluisNG+DJJ6hpZHRnF7D4XphTYoOSY
0ccN0NmVLU6reL+YdTIY4Km8B3tCZpPIVhr+UXn/S96R8CNM29KZAZrM9L6BPLAa7Qg/h2Nkgd2w
VGbPZXS0ko7VSdGLUFR1MJXrNxdzkHKYDhYNH3PyxmA26YXnzahRu42MvfBiKuU0IvIBb9KSDliH
PN2BlUzs1oZnT0tlHmVpjCco4KBTaV7HpHj82Rhdu2MO5qOavWxivDFVjoPPcvuYYM8vCXI03rOA
pLAEXk1lmoYtFtnR+d7laWEgFHn9JabwzEWlocZBsZWnqLRdnSQyQ3ieKK2OTCH2B7ZlOj0Or6Tm
/g/ehG562t/lvc3AB/OnPHJiT++Cc2/z9UVNXZDbHbdLVj494De1w5KE3enRTY1wIUXhdvwHIJJj
BPiMM/8L1n+BQ7SfSzdjfNMtSIfDRGkkgWTWlmma4OhNEnFXiMgGfY2NhnB4380YWVahtNB364RZ
sTqOYHmvXMx2D5b4Xvnss5TTNRcgzNAnCJRv26ia5ZVmYlyiJWVbQA2Ja9ZtP6rbQXx3UdQZ3/t/
KGNRAm3GoweQAOBPbKun1QFtB2QWxpvqZOZYXItekFxJU14PFO7J/2mP6UEMPp9OyjO6LTnx+ip4
R3qu3yxNXi0JqlRmmGfMFo/Ib31ooRVf/8AnCEo6sGnuWZdqGS+SegAXhmviUNm8cD9FcD22amR2
FyJNET3MaSWXGN2vO4GepF45QKq0xEiPXoJdT0oyTCJQ3d4sJGBFD/pjlXxYPk4YnOb91zsNkcq7
8RXfyfq3IXjzQk7qkpDPOV/TUoZx5otcAhf9Flg7Q4ek9B0eiw73AefAPtWGvBBETmqAmMmGAdQj
d7/Y2kNnlyYjhe290GbndaNGQ6PF2xga/mG3+1ZpMhVpAEYW7rMbFYXr/zWfbmGmLFV2ZF+9tGdp
sceiYuZhFlLj1pAHm1s0Hs/x7ieZdy+M6Ns3Y3cIfk8ZFsQrjHs3muYsI8hdbp7V9x0yjaA7I2/z
hJN41tsTssyPdE9QW4ipZ9j5AMQ12SLX3zJMQNh/aoiexbe5w8787Q3HFGDbJ6SN61RD1tlMiE6V
2c5R8pTP1Hx4myYy5Q4NR3NlMBMN1U2pTZfJ4NJKyx7j/lI9XiYyeLh2mYW7YJMOjMgoH0ImutLv
dOdKvi8Cha3fRSlcGtlCZhxy/Eq8QPplElsAx4nl+FXKrvscH4i++CH6B3xicIHXWudGfvW2nenx
80HhIjiyeYzOfNnHxoxx4YzPi+cfJmDWVAlUsRYYTOxCzbKgsCit0lEzTDHEhEALeXlgIsvOxm0T
mRVNLF36jcVj0N4whSz9gXbrrnruMaOwR1rb/uss8xdcmNsx4Oc7whRzaE0/pvERJX3HNI3thi7e
pBcoCEi+b6xQyhkfnEJ8H654IUkzGwtBx9Q7F9OIaAN+lUeEL8+1XTpqbH9DmQWzd3pdlg5v+byP
TTRW3nHK0idCug+NtJinT1q1srS+61iC89DODvfvIwf0Y+DPcjodz58dX/POPlRDJI/oSzu9SqXo
XXSXXbTk77hSCPu8Jhw7eJg0FHUla+xKCLmxq42bEO4aAp6Zxx5u44e4nVZ9Vai1On3oQzVNOCCg
m3hci/3eiiHneLEQe4lzWyVq80dibpyVXLdm5lrSePKdIIapA8FS8Ngh1LIM4vdb83AqLJ36Hf1P
k0Ap+WvjO3V+uL1gEUQRed1ybOkN+ck5uiWqLXuh8glVV/cWyooUm/tu7UVfucE+8blS2gO6Q0h6
mt+GT4QJ7HNNFdvedSReuxHVDUZoRTeSM48Ig0tcB4bEG//NqKIHb0vPVq9J47Iiy5yTxdtJ/P1q
Itl2Q/EpfP5CLuSIiHlYcofkc4wcO+gWRnrIQUs6BOdsTJBVd1sxYbZ7iKSo/cjEy1cRHtnpmjxe
qv4kgdxs0x8SzUjfusXoRc5NXk/4sBhxMXG305ecuyAzKUh37AJ3CaxszM9UPvEmrW5XhOcMIv99
LBpLV1hlg0I95tESHIsPY2mHBjjNbcL/eoXZxvInAPUp0Wbg2oY//FlhOkV8olejOzR4EhDd+Jst
v2NM3Z3zZ7WPDQMRWCSfc2MLZ6EFvjjOU4qnIxRj0PzMHLwOyi5FePgHaqlWbtRYW0atv0DDhwr9
DwtVYgFd9zkBqhprDRGIhqV7eV19pKLFjf9b7+kwmCu75MOPL5qfW9YzxBen56MmvWaRTmxKuHUy
6W5KaWj3XSQfMv33Kf39pfhqThF+h2lpVdM1Nl+C0jBQmmkg0E4bShkhhndJKCzJ2xh/IjswnXRA
Fe8T0Fp+I+HyC1egvLA99CXKV3GBcRoczMDhxiZjWoX94UpjIvFlKPF2YU3EvVCH+vC8u8+71JAU
1xO3/Gma4h1vv8CplhdUQ7dmp3EyzhAmmSm7aCGueSxYas9lNeyix3Cb2ATlP2LO+P5eFTFYl5wz
QLetgXPnImR7dcPCfcOdu8dzME+d6Qj8X4Z+N7LGgjjidWpt9TFwfgQyomEMCDqk9sev1ueJOeeV
T2xM6MhHtdoL3FzHrD1YseBxWzMpoBjgs/dBEuYHmqyv7n3enNMXsUBNLqCanSpJezls89r6irF7
W5pCDY9UF04F/kKXDfUGXrea6SUTHzGeO0f3PfOxSos9UcBL+xVoesmfuBHFsqjYdJ6KnOu3k/7j
YHV06Y4Cw/yTLgfQ6V1KidVQqLGqVwYPDcw9D0q/akdu+w2WJUfcWS7hkLZjacWtodx9vAz2kYbe
Sk7hLwU1PvgPITbTpH7iTLMLP+/Dt5DJLrp01NLs7kdSulg1WF/qmGcTGQ0KBFNkCLxXn3xNhhpZ
3mYYrOL2pGjFG+UrHMyEcx+zfyckO7pqBuFUdqwUTVNKuMGY9sn97c8iq1v2firxEd34+jZXHNLQ
CVVt0YUJgantjxowj4UlUNoXl+ChsI7hv/hLc4ucQxrLlthwkQuyeioBpskIHcgpZjwSoNd4wky3
ZeYiCkfE31DisP18mmmJBBb9tPB8xldxi4Smo76ehg8Y0REea19AF8RIx3b6inSOFAWQFRiOkXAZ
OxR/hsO9D7F+s2MF5aym1iymdH/uoNoKP2VxsieAb1rQPpM1wLfFwuio8KER75BjdyBgCTWTMa9I
j5/VaAqhNKk4JBR2j3PV3TgLCAlKQytoT8Wtso87qjhNN9ErhbHQNTGTQihNUEAdKNKrXaVah3WU
Qyw3c7kc4CoGoeZUtM/W9D8taepgsONsUtIT28LcOmvlvNx4O/lK4mk0ER25wALrxp6b9WCdYyQk
bX6SFZZcismDxWRmboRBvvAUJjhBanPylVrzvaePRI59o7m9EgYA4jCFTRM1a/VrAwd+EGSGjlvv
IaCj4VAIVoM2DGTVICkFFX9JcXEnv1C9FVEp3hNHMjOHsq7Axn3B6FSOBSEVQdalBnmdx/vlr1BA
O318k3VEWlrUYuIkvEd5UXUBP1d1EWbupkdCndvKKi4kzKcqzztEqEhY1qgfsjfxCaMcCaiUnMZd
hjfARkKxmShG68VSlPBWPmIoOjsdZz7jcCiE1s350jgNr9G8sE2cOwTdYqS4SN/KdElfT6RIznO8
rH5bZqrl+PVytTrYGBdDgQ0XnVhCArkKLdKLcptvFbTdp85coZ3SMn2WD4KGDFwEtvXhxVG3HkJf
sAMQGF9DQ5fccA6PhGSH3zmApOleUdYiCkkBv1bVvVmjlWbmc2Y/WedjgNUU6FtkmQ6yAKDQBFno
zqJGEDKrbp5X8R2el7oQZf0BNmnaI3654esJ42/D61VnH46rfUNnpgE2hoesiJsadxNM4Zi/gqOL
LYm6JQZY+Y5wty5jxSYTWCJUs/ZjXB1zCy8/oWiM2xACiJKTDQMKyg39tcbXiLW6jpcxoUzTRRsg
Cc2FeZBMA5JOHtxB1VDbl89e+8fJc148y7g+0iK1xyJTEJL0nmjTzCwepIRKvvGsrqvmHwlvgMGm
90aL7nQw+BaHZz8Wi0JyZbyYZ8NUXpRDQdMTqdtABCPaX5LVPmCMpoYCnTkQop41kdeH4MpjpIx9
6Wl3WrmkuQe0mdZnSccl9G2+IiyoCPKGFP7t83kcnqaVJ5dPvMZol/5SijFeltDO8pgLgpWPf9Mj
gcoO7NMUCVUV/1Yg0pa5OrAMjIXFzYb11ZYwW0hDSE5/mwbaqpp2E8HdT6icF1xLR6MRyzjn8zeU
oxn4gTjiUcEIxZOEVPd+V50+iM6aEVh/zJnkPlmfMVP8qjQpJhLCIxJZT0BpA6lchpwF0klU9HAA
yXPKtUWRTqml66l0sacg9HIz5/NFBEvWrI+NtXVZUCyZjoXhXuEGpatiQxSMfCUt2CZeTbW5TzkN
XxbksFT3u/V84zDUneR9qy/G50iXVonGMtBFdMJwL2XwAwv/wvxoFnjy/2B7IxltIZ38WfvprDaM
A4JX4n8rpHdO/6GgFBd4SvTKa4FIkpx2bancak1m41HZZz2IehOmsXvFdpKd8CUUHLo6AFCc/CIl
DHQvA61QfF46m8s7lmOBswqTU8h1PLjhs2QfoZCYGqWpqGv3Rss1NzQHF0a5r2n9KL9vjr28B0R0
LHVpmZ4IJOpncYDK8dhe8aXXeqc6gpMFOrCSU72LjvvM6fHh3bCJTvHuabgrJx3VJSuVSyPQ6z4/
oHdIUWeYJDVYeo0OAut5ZXjInMAuV4jKlqh3CA86CsYesxTpTfmYI9OnFKgA2bCtSRIRY1efI6/R
8D1VUnyguY6Nt6Xe+UhwTf2Ii9KfkFHVNJOea2DEHkj8OGaaOGLd8KRC1YM7TYr59YZUn3mPrpjY
fI6LZPQfok9zlxEp7db+wAKUCU4TsG0ewOzfBGrzIjCX9laJUIjREuyWSzkN2I1tWCLW6a+cBCaI
pTPQjffBPDXbRfrJkPblbYdayx91PD5kND1YW6hDPZYtSjusR9K48aS39g46yWhxhpY1sFYHhkPZ
wdZulNpAHnCR1JBSs1Vg3eNPS5PXez8/tR4Jfyn1S4pP/fe5JgkdoWZDAi2tvPTMZ8f5fhNSCbu3
QW5RNT6w4XU8VG4OHIOyKvrsDHguBMBnSb9Kda4eAQwN/WtbmWp8gnB+Pqvx1Hl2r/AJVV8XXUzk
OXPBhOYhYvSGLIq8I6V5t3YWpWPaSyyKdro/q1L5OwV+I63Y528TwRTU+moTTR1QfV2cW1AOfdJt
6A4EFkylgSkx8qcuzCiHYmapunDxIhJuAw6+QgJOD+MEdcgXgccA/kBXTYTw0mboOsnlL77mVESm
wD+aCy9tf84sYxwYiEHGf+TnpvgXgVhxJ+sbMMX3a2lskZjpMvhdRm7xO2KQX5/Ji2ErcbeE1FuD
1cpqjURGa3KFstInp5zsy2iFFmQsbjLWZkhQ4zgbIZH3IDbTN9KTvpX/CgJYbsUpJnVhNCLGSWBN
FveqWOq59Byy4ivT18/WmUFrnRbLd1zfTaPeUGH+0hCxXRe3SnMm+RYvzdGmpfFUz9G4daO3X5pm
pDpxm+5I5Znk7Ch7Iv2kQ2UZmFZQbKDP2HUVgx1B0z8oeTiHyw3WxplaACU8zlDnG4DZh4yp08Wp
UjW+L8vHYb3pYILOIZwp0+nvigYJK1HCYQKfJW+TS7DrrOCAaHQOjTYEoMC+MLqwCCad8m0AIEpm
hLqda1wo1qNyq2hSdv0+LaqNtMJhtKGcRZXwDP4modGxRecjJQqcQeMVyWulik9VIX/lYH5yjN5x
MIDxXARazeFShJ3mqdqntOGFzLAepFZ29r0ka1Ll9uarhyQ6+Aih0x/8w4F/oGRJWVkvbOmP9Wp+
VM+MeZzpJ+G2mw2F3u76CEVZyZY95SwMxWhMIcQHfFk0ZhvR0umi2nopc5GnWOkIuM3Jr5MCSWEL
KeVAFyVrr96XM4Ndq/hp9qW89HngIL9mAC8MPPw0dxy3im/kNwCbXv4wUHV4vMDSTxgBP7SkVBZ9
oQpQo6Prm2sNncmJuuxz508qWTLjwyNJyBwhMC9PtuE7Gu3vx6hDnxVa8AP0ZgZv3xnHDQN8KXqo
GLLXDChsawuXPmuMk1+30a8j5fSHvl4hIJAigkkxuB9GG+rvC1ewOQoXGVYharjoQyQb23OzBCzP
jprIjf78/GkgdMErI0B+o51EAu5p7CBrFQwcY2bgePOBi03/DzDM2XlaqFNowh9wDzT7OVHJ4brX
/O7XImoviyqOI0XVWlFltYCopLpqCcl5mMtJui3O168KctTplT8VA8Im06T7gM3+nCb5YDveFW9+
xd+8itYVtd5MtC/L2zpLHWihkqHpi4+GUxtixGJFmyZrlEPfYtVWSSjmT1q93cQCx1T47z30kAUD
AU7p+DnICZYJK3+1Sf6OhA4bOGeGThOLjsJy+WHSFUV/Ni/+3IdE9B/pgBcZQEnyqc2vzBd084Va
huUvct7aGHWEdtdKHifrL7NtjEw15tu+1Da1AQ1AcGBGE1C5PrOt65u/bRVpH4vlDJFLhFnDdL+J
zLhP5lQf/B7ovoc+Ws5hFdbMWvUB2/NnqoKgroii3m6WaFD4wlSvokVTD5Glwm/jX13hPUU1VNna
lIb1pA5ZXmCM+CpGwsBwaBB4RJNOaOiBsURF3hu+Ut2j3tDWwJjgkmXLeiMDxCQEYVsf9quQ/5Or
q8M4WPhEVrHhXBfc4W+wbjxQa+8ujvTDl8P75QpG5qMXM+UeFPi+zO+fvFbZkfRteS5Hstdrrt69
Lkli1UuQ15L8rJ9VF+zmcNUEMuKJc130eRve0xGavpxwDVbTXbnOm3nnhqSJNuaJJuxFa+DjXuav
ACBjnAvreitnXrvgH1dKYOyt6UKUIZ7IguATnHThYKZtwyanhHe0WNTRPXrOZcLaea30i6rQKCKF
wCyw8MM+rX4RmNyZP+ntXHYKXKPiE7VwOv9l6Lws86QHfhXAg7Skt9ewc+UZIxhk7cg+ZJdsWc6T
pULrzTSJfKYdf9hBfouV1UNrApQ1pupMPX+6sezUmVXwul9yrP4Q1O3THvOiIkQ3ncJ+eeICnubY
rx0wCZ9zimxQ6tPsAAhbqGAyi7+wDdqfvOKx24sHZZSSW6ONAZckHBhEonr7HV5RTsLMS/q/0KmI
ss0HfoC16K+6lmLagY7rvydur7ZVcAh3/y2zH27dUI56T1DaLd1DG640WB2ooR+2MJDJJCDtapCw
An6x0Z5K3FhXv24Sg9t6Cxd7r8ApjXLsxMwykP8fdzquXiaOGd4d0rfs+Y6qhhlzCi/kP+D7MIBJ
MOb3RLScVp9EWFSbxah6K8bI5VOk82C/e+zpXxWyvtL1pS8tTtKH3nzsBjetfDEjgoewHF7S92Of
Ak1I1IFNO9mczyGF8/4B8BKkSOrgW+Z9YC/V7zGxS+Fr/IYsZ/jcyAoYPRg5t8ejnGYrFn+EdC3d
k6T0+cYoKhyhqiH+aEgDLMDmvqlaQ7o/04qex6EAY4BMMJP8gDjWXgEV2UtQbJTAZ6TNIRaQYhHJ
+kG7jYUVStFbnbpvLNqKUcIlQ7wvTj8uUxorEz+7AFFbarQbFp2TI/wHYvw2wi4rDy28f0EYqC/M
4rIMzDFMR8bpR1khHccBmRpA5F6ivfQNEUXiv3C9YWTm2OY2xyq2bvgKF10B5EC6YgSoCeL5FqaG
hmY+pBZ2W/ZHjxPyDe770QrHb8DsSOfXU6ZYbFhCN0vFzFIs4KnwA7nhvd5Okc/3sa5o3xPY8P8E
dPqi7uifTYU76rho+LGTDIGZ6cvT9V17D/1uxRifRsHmyQ+6k4lxXO3/KMnac8wcP8Rxe/WdstGl
7mACmx58NqEantdoDpDlUnM7BJYLcZ8CJCNGH1EuA7DLtZ+vLqetXVpPPCNBwABD8p4bDDI8B1+i
JvVeL1OnBBY4QQfWS84yXiNbv/4W119GWxYbEqG1cUaFX5JnTRTAPqHxm75mCBmpccmR1zuMBUpf
QfmSY3Ml3YhYEGhe5Pf09v8Wh0VFvBPNpy2kwd30EEMD6wZTZb/exRLQ3rwt+qI3vvjeiyRkfKib
uHR2PFS0kDZBRIViO9ZdEeOoXergp7z+IJlYpMFZ75RWkl/JXJUr1YhiCnoyMWtxLmkVSF0EGCvO
QLejMUBn/N8e0JR489z4ZuvhMT+bq6EqcfivNkH89ra/EcaW77GNuUktFGXBYb/k3pIQIHGhwXWk
J741ReAs9qpVIBfv/NiLFFaWW09Ewv74cegqF+eYa0VXlWlZjEl2hI2G0eRiZBwMMMyRlXsayw0m
IO1SuER/8njZS3YN2EatHCBuSRFKxtvqwQJk/CyYCOTz5rLJcvKdJl/8p7j+5AolPXiPpk10iKp2
ZjIGtdRHFJJwIp0sJnbTJQPzBkOOim06NcvXPRUmS6ciVGO5wGLrMhBhCVZWShYSb9Wi4DQmo3mr
f8pDskqNee0zt04YZxHSMgdkaZOkB2mQnQkbvSw5EmzHkTKaPsr+TTInRub2QJNUntUj/ono5vEC
qdmIgTSWtXrq3ItG5GcLcYlcNPbqBFR7YmCFxRukPdfKuFRSPJKnfYpFE0id892GVlR+E3VWoiws
YkJ7LBymcYdoqvK0EjoNAUUL5Y8N1dEORuGY4pqSz6JVxbbqTj3Jdc0arBkcDM0ZwI+7W6koY+s6
eyAlC8EUj0G43tOJDmaKTVH89g+TjTZkE5+TChyl038upwT0cmrD8FJbaLafJmTVy2f3jiXt53MX
y+zgLnRIictVoU5c0y6w7O/5k13Ror74i5tYxvAbYvPOiI+XUOSeFEkhg+XrqfMXNEO/WMy+Lsvw
zpsn4mFcImOyRHNtePrulc9RAAUlqGGUm9AOtZuefDEWw2rCsraTl6t5fltQQiZITtmgaqS3R3zr
GER3uh0QZNJAAZ08Ht32KbHToKaeChb16zkQg4ZH2ie69qgWmjmntJvAdeNvwDiUmp9EIffw/M/P
Kz1GRm4F3P6ZJW9G+0TkCo7IPsfEIji7U5NE2LkgyLgqd20a1+mrC1sv8fWIv7fv3C7Rc9fR+WQ6
rpP+nzVUxFojpZVVbQHU4is/DZGcBvM7lbmCMLmFbjO7P6iEqAKRk5ccAFUbyDajyiBijVRCPcX/
HkEYg77R9pfFu+Aji/wVRXnAzSCTpyC2lP9ryMQS67mpVyDAZQTYOb9M1QzKQlh6yGXWz8G1Mnwe
HNLa/JvlSK7PxJvXnBiRSGtAViOI9VO1bBSClcANbySu7uDA2yrnv6sCkwmGlCENidKMisZskf+P
T2lvNCv40L9PxHqwR8Mv/I7G2IHRnZFdUoECZIAkvxHl6BzaWVWjvJJBRmbvQq0K8Pd6UzlyQ6Q7
pnxpEN7ng7iPUYtstVAo3WjhwKQRBMzj11Fo+rgsxY3JQZ/+ogKP6LoSUJTANAyAp9Vske5FJ1JK
XGFy06uHFWypq2sxx+6hdMTXsHCrjMaQqgQ2PS6bX4Vha5PyNudwaKjbuA6Ow/qRs/aCBrE6dDuA
8vz46zn9FPbIkpG/eaw+5J3rOc6o7KnVj1EYV30jPNUHotN3rkk9N8GPorcg1OVCWzQiPVqrRueU
9Bbt+7jetB5GRpbTlYfXDFzSI1Z2/2T/h3QNM/X77IlNyyH+rE4er5kKxD1XpmkejWtnKD6wCVy6
IQi31CSTJV2HK3IxGqYSuQ3La6XaI7y5WTGbqCJxJHCtMQ1YQlFU/VhOSCAcQ4t6INCEAdsiv7oz
D8Tg8BU0NE8txkLnXm5kP8eDYNPhMYP8PUakb4d6Shh5eQaAOKINBA9sGpdO6nmycU/FDEU2PL8y
tky+9SotHW0bcNXWnEda674Eq+F1xzMkIC6ZMZV+W9JMc7cU1EBvqYIyQrvakOWjZgA+fppLNaI8
pzSC1rdlvxm2eF4AOBO9Y7TWNGkHtYGcXERpjIMozRsHT+Ez4zLBxSHoAp2od3VwIU8iSA6+oHIe
Q8IneN4vAD8P8TrkdeUCAJW6+GiEmde5FVjVKs9A/SshOUSbroggpHvf/HmmW0A16wEs57hGzzs0
+gVLcdtk4/1eHeyBzDkEdOUAmtc8W5C2r/HcYnQABVwcDdE5YzaB+wIs2S6dHzjaCieptneCQTlT
GkcrFZhbK9smc5QtGJ8sQ+CH27voKvVFB3VsaYGrj3g8XFw/JNsOp2lW5ipzTLjgHSC9t57cRJQw
AkcrdjrI5F53lpOpHgIgV42D+gi4ZymceRBYanUy79cf1SggoX7scvELlYemjoL+MAoh/ruzQBZ3
xGWAZ2XTFQL4xoQ4VVGp6lim2bcLdUXxC5q5FSen0hg/tqV22SoCLcNAdrqRfYiLmBmJacawP2ct
21MvMrvw70XraIsjzQ1epeI2AL9HCEBvpApT0GhCHj/hzzAMkiBZSmzJwYVhdMERCQIlH5PfsjaO
KCVqkEwB0OuLE2DZ4T1/qG8UF8ZAJ+EZTKlLeeWTXSBQDU63MtgjuutLnZuzSlD6N1TUHpOA5f82
B5BPaBhMWWZxZnRdkMW1DarfZ775EBwi4SPTvkGVEVMapUfwaZaYu6QvfOJk9UknkjIdX28cfGA0
qjUiP9K8PYr57iSfQAmnF0yhYiKSj+HClX4x1TuJzc+qnKrsi8P6C+MMvQxVzwmVE+puvOYrT4yB
eVmhL6AaQayy+kvac9XeTOGyYls7LLjEL31ncjGYZmNU/3gjqR5B/S7amqHrGleI2bFzPPLAE8Uu
JS7eCjNRwhXaTJ9c8A5rF91QllGlb/kRaOblQziaFn88A72g9pKlXf1iRSSzsfvVSZ+NFC45dAxt
fqydaBE7cjXLvf9e77hiWFAmN9HvsKrVTHHQnPg/bz5mW+X6Uoq1qpnvRhDDsgPmz5p+c6JB+UAR
cTZexLbxO24M0Mer2OkPteu4EQrI3aYIe0BW/iurV7Oun8CrjyWqrdOG1EwC1kd3m08/wBMewXGQ
bNaXDI0LuWirxl8Sv/3Vi1y6uBGXoDcKY8Oq9DPszwjKijXV0KBmkBtoYdZi/lawu1c+sSKamfNm
gSbTKPHNpWsjfB+j6haC/bgfwP2npKVfKr7ARucdQwxMZhjI2H3Sh4qHIXGKdRatfQ/EidaNLLk7
nxsHZEgTVVlhHIvgsJ/xqvjKCcs92eFoIYDEooGZM6R9PInqNo7E3AzELMgvbDp95Z45cwUZldB2
kdhjZzechrfdZZ23Nwn41KUY2rgi020thlkV2glAcfcJI80PacPA8kjd8SbTu0EKBiU3xmc0LVFw
ujX6TOD3km6WiLDk38co4Vs1sOSQzhCZbwxeZ/oMfI6wPf04vc3jkP8JCdOZBk0ODc+WjHUaAGTV
hOgTJin0zPdOsiyjKpEu31UUy8guRPGeel9iLq8Ck9S+2Es6UQ+yjV8Sc+IfVIRuibX3BvjcBlQl
yaDojAbyNVxYKDL95Nyw+jqQGdvNjSa0tbRDYZX69uk1Q3hvUQOVhN0sUU/BM+oEHZuCde9jf8/e
j08i4CP1qKHZH7tldSN336EuApgCiF+cj9aU4uMKWbBQVREXAF0atFqi/j3A5wEE2GKW/inGGWV/
Pza0Ryz/yuwrhPiHtRv2FLFM4KLUHdOCGBCA1k3GqntjgpoxaqsVCSmdrCxNTIpvWi1Lojco9JP8
WpcuN0cj0Yc6Wn+mcaq6OdV+Gc69t3Jy6cfKdHLIg8J7OvMxlca8GfAo/Yw/jdEa0h2KSF9du19C
WVoVI7f5k2YszKzh/U2bcfodt6zxnRhnl2bnAbKdUeJqcIoqpXcGTasl8u2bEnD85uie+AA9Oihm
o32f79k8xtWduAOQa57oq8/B0Ldj2ec/pAqVhWfcBU/lLHdCv/+usTmWTSjfgTzw7EFkRcINtgYY
OkCtJ7SVZFnDg7IINZXjM5k9g+5exYQR3pW9l+66VifaRX6OnftwIKt/xGmVL5ST2ittq7akrVms
AMs1qSwZPa8Y6IDfwvuT4DkwBZoDDyfRaa2AHzG5x0Q1TucAay0X3fVu9XM74ja+oUJfMtF3g7ro
cLXEdLfF7pQHeyATM9vBv0AigzDb+tnrfCcffCGwpg95Yy6PXGIH/CSf5f7V8BgAUnCj5PM1t7W7
HyDLJ8amvjht1mukaCi/+iso0sF2C1B9EkS0mS1hXMNRLuDXllpB4roPy/gL2R/yepooNhsCCowd
Pr7SAt58nW559avBa+0sFGyH/1nQhmoc+5WrkwP0ezQKvIR0bCGkzQOPsY7cXopsI55YBO7IeCQo
tXV2abAiTpxKnHvd6493KbeXPoLTQ/rlGFN4l3XQ4E9PoaWz/apUkKAMyf6JDsVmzfmTAONeenSx
T4+32e8P3Wa57yhxnfJOWegRECG+XAZWpyUjkw6hKg+2+KzfjuZzTKnCZPEjCFqL53t01Ql5o+/l
hBpDnpGdfPswrSW3lyNq3+XdzcSB57FSdc9HZCRM1BaM4n5kdNC9aRvaggx7OhY5Bpv0TCkQWq/F
q/M0/yzAsnue75lqq+KdJCSvu2L+HMMvh93HOAIMVoxuuxmj9Qc7ufPgIjgPOgboT/lrkqiFAXUG
NnhrL5AlEjCUFSaDJGO/P0fsdO7E0wyzbk5KNfzpFk6yhVYRBGcTPSFsr+56wCzteil6sOOJ4LIF
1bsjuG/irJTgJFEuvbXgv5JT4pNDvdHNRkd5EtzU8TEBpsqLBtJptTqXwn3LhyQNcypEGH0YsjTu
I7Dbq0ZF6Un4bVlahSE6cqsCsM/GotBrEziUjIfKTJ1cIf6VfyyjpiMRkbitFlRPn2Y7oUw8gRyq
Dd3InLNSIHM4x1VIK9ahEo+JpbcL5gchD4CGUxdzJDS0Q74TmoolayZw3Df0DzGTQKBRcbl1Dfyq
AA7VDu9Hcwp7HYJSj26VABmnGxiVvwR//tUSq1aJHgeE0k2G5MH6sN6wvtZ5hzIksEVdCGV9LwKE
rxO3sCl4TcLh+5z/ikbB4bMT/JU6ovvRZi42TabiEVC1Pdgd7NhsbYRX2YDaPj7A/oJSRtHdfdKs
QqrBIzJa++KDKQEkq/kUzPtUhidzea3xuwM6x40uZ2AyJBZXUhd0LrcrOC5us9yw7eFlkwKYXUlp
Y7vnxHrhahUZftHSO1ODmK5UAnqMOPZRmVPhvAhoM4/nNii9j+1TN8v75qLlL8fspK8sPOc8PH2N
tQ/6kbbH2g/8b7puxSzVh5D6bgjHw9unBAVhAIYQRQhEv/FLSmOExov0141N7XNmpax6vfBKo8SW
724sWsE+q9Pryp4jO480axA1aT914TEENS9OfNLLNb9Tp1KDo3tvIFXxw4X1R6lxG1z886EILMgR
aVBZmfu2y9xlPyysXkPFUg1HnZMyQSQC/UPzJc7es3FMKD2c6L17ucffoqWUkmiOcRxszW/2Nitq
fIqSALdqTAzsZ3q/Nw6xeD0zD8qx3DCOaLYaXoJPDDB/bHy6+Sf4Au3JWNDsLUTZTg/Sfruw8+dz
ei/f23lu4+B4SCIV1OA/0WtJ7ofvgY0RMFfg5InoWYzhR8/fNyDdIO6k9rL8HDop68v4LdeiTpKo
S1MNtZQPDRrj0GeAfHzrBnGuYvREf4Ul65d+PpPhL12zUHkrv5abwC95FgImiDv5jVZdaNbvnH10
e3t2VbVPHAtaNczTZHX7s5GNKqUiGrU8hg6SftCY34wOXGmTnMfxK97825DUQ1gsmySCzy379FZl
EOJOPDd/WqUe6sbMBtMbpHLZt5z7FONOZle2KGM42P+Gh+KP+Up+/AghAaCaqhYD9UwUuC4dWERA
OhHGcJNSVpQixA4KUFnyh2h6qlvdocp5Kz83+QKevuvR6XdGQ9jsWB4AYFHFjQnjfVTbdvdUQWpp
wjCYOAI6njIkiAwdfLPyIqNdSmorssBDKRDMDC6AL2aedMjvf5L/gO4ZavUpHxpOrbdCWbbWdw6I
/Y7SpjN+koS5UoE4mDudDfrKCFkbvlPtvPsalGRFgnjjbsQmbriczJg3DKs+90De20QMmgWzwnvF
cX08Ii7nrtLfv/EeAgJ5nSSsKylaWmS+dAc5LzH0OTV5kgk9xuuUcUbyKU7bXGyN182BW5jZzQN/
IoOGPfgzz4o5U1O7wEkl7Bq3H+UDGyR9MmBtmIGea0h+4UTWIEAIjQ+xdYC4U0Kfu3DMhG7QIGa2
cAim8VXq2sjTN2azLe14e5u+FrJFJ0pGofGwuffXgOh72UFlHQD/AGIts5oQ/hLkOBfZgQ17XGm3
8uT4xUAyzDJcOnWDl4wqoWCoM3yN4Bd8V54rKNoSnMdy1RFJKkVLartygeItF7kIFItICNrKG9rP
ELcYDbkzaj6R3Eh9jOylMDGzQSPD7AIQyVpXRQpVbaO+jmgWnHiTDa37vOwNrkTuFvsfI11sZh04
s4sm+Pb0TPL/ekSEzK6inJa+69bV7GrWoLZHRZVEkwCTDu1plyhtXb/VuILj+ckPnRjjGwF21qda
a3AnS/8mDLis2Fa9pZcwP4uUkp1PCE/8YFTscT3lYjszWUjTvVTqcScJ/QwPi8XmCTjZRHShXQoE
S0fn6ug8H/LEwY4GMnx3AUfIVRXOwNZFU6uAxfJfRnTc7JJZO4e8dflyvOX8lJn2QggI7T+1nPCD
rTGqLgPLhxm6dISKQOQ9rgp/TUla0Swd9zPcq/yJXXcTqLhmOVhipiaJRHHB68HldNlG9cZ0zPWq
XU19DQ8x8e6jBnoBz5RuUnFJ8ttKGtIitTC1Vi6A5LVERwGnemRqgrGQhtxqZPrcE2Q5Qdb1ACmI
ImooCrmR1auDIDQZx4nXnMWs/xiqHXZZHWOxBOxHi3lyLm3bVheDI9vAl40db07tVT04hvSxjYMR
K5J4ot6SsmGWGum9k8sRw6zWxEBjCEssN9oZ1x7HvGcN5MFuQKj7niV8bDErXhoT07wvKY//O6/X
OEQQl0wAJXfqX+lkF1nT40aGuMDj0BoA20TUuZN6amGMpPiYGFCzZOXujeVgFg+cKsYoZRe1uI8E
mU0I6xGhc5afMHorX+LH565RrXCeBXWj6n+UaaO2aQBoVpUHGRZLKh7aC+dAXepkABe2lB+TS9sC
rNb0SbNtOFNUBdVZOnF4O1kI61+DckY7TAZsZ5jr24shmq8CVPZW5yp7OEWpq5Hbu6/BMmExG2pH
8qdhzgnSofk47n63csabUBbZcytWBYXfmJCqoSGBIsas3wDF8OMJW9ayrTdbK5BhKmwgXGM8t0uP
1o2KglJE6IqK6uxVr/osPNAeQ4vKamldYl/1NF6/zuaOTE9P5wg7fPUuA3HBXyn3t1UFxrRXubkw
ELgU31lD5GPqfXVi2Phetp8B43yNL0DsauWc2vkPksIa7zgCNaSR8+sDuaOEGOSBkthc610r5IKd
qy3feV/5127OVuNQ1Ych2nxP4yNS47ggDz9pZzev6VmeaH0dsHZ2jdBN/9x6dagO2i3N0d/SHeHX
UTrjUj2P2FZ6fZm3cQg1NHb0LL2JBcdpz9grCM1IdCOggbkK7mSl14uJMcR2GOehH1Z0sZ0Wvnnk
5tmdUyoG/IpVuzKWlsLsgwjHqa+u2ehaTqAPiZ2iKne4gWQT9dYJc/KxbSqDBgy+0UaNH/XJHlMk
A+2ceWX55B1Tqz3PWR3KlgkUNVDTLpxbZz8ZXzUc7/hZWfnOY5/YLjEPHyKOzDPGj2r4bWETU/UN
sLzUnqw4HJ+UumZjYXbM7aHEq00w+kg0YmV88DNpdMdufC0Vmj7tKOnLoIKOw+NAgk2JjViwYUyl
VmUWE//oK3UWg5rODyRXJUyu1xKC8Zww3REhbDestPDKY/eCjWU3uebWUQpNxpELuzE+w5bVv0Wd
nLRlzOTyaGBxpDvMpBZ1V9Kv//yd5/rntHcz+0lXpUBMjJcHEqrxVrqf/s2f2xqumUSRArd0mkx1
afGCCwr9yf4BIyzDBaSm64T9YnPLdZZc76Ty1I51P6A5eoua4RK3Vk0nKuYFdZfDYZ5gYoCBLwjn
cPvNez9I9xLkILbAyOZ2PZQshCs+FXsWm8PYwz78H3JaSSFbZI/llu6Is21LMLMGaGKc563+RW2s
VkxWShneYUsckHWpKU83HRmQMdiiZ5tRCRJk0p9JFuein7iy6X1+gpe/bhi4WmoAKjalmm957K4R
8I27ctNKnfAyQMnA9lq4Fx5J7ED/uUhiZfFUxyHnV6wFS9w9bcN1EM3jXtUpIuH7R/bawbj7RzdF
OvHhj+Ca9SI5TmIE7u+Q8OVGtGJ1m8CByPLlalIR/RB+BqPG8BuSzCCSbrPBMVZuqhYbOfFh/mJL
0UVXLSu8eT7f7DqRllR38W6CebfRkkfIFvmqBwKNkGRE4eAdl65wj1I1sFf1DX9iHYWetlsPRszZ
1MxanwBfQ+WZj5EI8KjOHFNicLLKVtdRbzrOgblik1L6fc431mIbrJS4IDZArk83xz1pIDNb8n1m
nZTnbIKHOBtbDoLJ1vF0RjGk+zTbbJLB70ilPFz2Yi+0zVVePLcC7jSPSEykrgpPA1LFCb4WtSlh
PvK9adYbcw/cLUNhGur1j4J7BXMufFGrfn5Fn7aql/E26aOoSpaUixp24PGYXWfyH9NyyoW5QXMa
wDQfMQSV4ebJMv+X2RnaDWwv3gipz4lDMZjYxMqS8RjN0Jf2zYH5s/sS3GAbfWT/xQuUZXBJuhPD
HF6R5ZGB7OZMpQG/TIKuEHE6LwawV/botzXEHJG2bAYGSYhgU1pA0OWtaO5FPUEY7C6XaaaV/o4y
fK08D0xza1pISI0LSzzbTECoVHZFmfpLSS+z88hMl7zFlf9HPN8ig7ENOp5b5lywXbS8KELY0VHc
JSo9JeKj1XYN06kv+a7Are5H1SAG1A2oHYrbNUCMP9Q3c6cGQ53B1LblwTnDLGcNC5XK5rsbQUfI
PDL1bty5hf/sqgldbG6uEZyQgSU0aRWRFRosehF8FFL6zIoCqiL8vCB6eD5l2h95m2srvBXi7xru
edTwVa9iqr9qYBEDnok0oGOvyswxoVHmC0pl+9oeYg5VW+dUzDCY9bIhc4J/W55m3JRz7Orm3Pnr
5sQzGPJjyH8C4mq/APrySgSQ5Tb1isDQnh8wEIv4sfdMLMWMrrs+vUonIZ4J6u3awDljZoqfSm44
vRxnHVldsW/oiKzPCxpLVPmXMA9jpr6X4iNVI57RYs9MYyzsAjSDMqSu0U/+RwG3BJn9trF2p+Dj
N93119x56mrj/AK7VHBOV5kyem+MPHsi5kUyjFTyqjYgDIoCO17OXAcNhGioKr01r7Rk6CkYCRA1
Qx2yrTJCWXs1S75DYPSYnPz3FRpdGH3WS9JmA0Q2XQ4w5vYOzMD1paz948GcFiT/NOYpQPaie+Ir
nBIRpptamwgQzX0pDibhfRmHmqEQyRj5mymS6W2GKPuflb7zo1x4NV9fU5Oo1RmJoWNlhxYETDkZ
zjYqFM2PEkhTebuTKgjRYeNP7S6+Puk2qW9x4PLfqzSJn9hDtrUuiphVC/J6BGjoxylObRIIUB42
pc90eo7laLFfmBpc5d6mW7ENXlCsPgEGItV9ok1jt95L3leQi4kl9KrojbdRzNHWcw2aEsGsk3Wy
qF4o2IG3VtK2ERpk4DyQvytwvJPp/HMAFZJjUVl9UDnBMHCfbTAVvsPYsTya8QGS+POkWMP+UHi7
wsRGIagrafAU/ratyFjeVHsK1YJz7dwG3VUg5ROg/DQgIq04r85YNRETC5wWc9IGZmNZ8OMzCvJd
q/cTiD5APGisyWd8oO9WqzQql8F+sVYwh20S5SmCz04GWXoMHxI1/SGyQphiUkqg/X0TM9NXUYlB
VXG8vFuPHgQBjsuFh2HkODF2/nHgF1ON50WdXDA/AU/I3fGhl2VCRoZUM7fDF/WmTIH5ufbq3DnM
IbgeeaNg/y52rcxaMtog6uKcG8wcI18w/b8L5iAmPWpvzEUeggEtjDExHOf2pKag7DV+2CMQKJXm
JD1eCiU+zR1OVk4RwVJRy73kYvN6YGcSZTpq8Bzip6avJvSbGue9iSizWj7tulnDbfSWQLlA+jFN
OysDw/gJsoLGYUVAWej6BYI8C79TEI7nra0NYIe7Uyuwi0Gz0h8K2T4yfgLQ6i0pJT7pVK4Ncp2n
M0W5O6wiZiN7giaepW/vuFIg18IXZNf67DonE1M3gKVvLZVFLdxktL3a6Piq5ZW6q0r8Zea7oHVS
PPSyYYUtLthZGs0a8MhQnbUhuooicjBfdBd86JvANpH/tVZp3G+/LAi+mvSOXyHBQ32KI6/xgVJm
zGtKCGDcBTXR9Hba/WjA6hdQh6xtPco71p+U8hU1JOYNM4x4SyuxodQJr5hZB1s20HiCi15WBK+m
djp4aMSoUWqY9FKIbHBTICMMJykekuQY8jzZC709dWRGF1eXY8UtHXpNOkaEKQ/xJglw/U8bsl2s
rofxbubjvUmtSoB4QGrXqhjasIBfGIsRwYpJBBAGywxly1Md/6+PRayHrRjgSWB5Ra1MUFiF9rN2
+XIksnizLGgM/n+8UJ9CO4xbUwhmg0MfsDq8Cmj/WjimqGRWeqXhBY27Z9c7g9FYLDCbUmliG2LD
rEXijVAGoiCako9m5kKu9mcSc3LTX1YHpqzt6+HD4hn+sMEPyu/a/9B2/OcqmYpiLCWDf8b1cVjB
0QxML1KpUIybAPsn+n6c2NDw9zOl5nsv5Qksmv8uq/cg0Qsj+jdRqcCnWz9U4yyuOx027yyWp2iZ
n6PePGSBttNeC8tF5a9Y47IkDgvoXb8qz1zs4Ef2LYPlkme4QIMJy2VfbQDgvPTdqCjo7Pv8C6F6
z9a7l7jBN5sbkf9Ig0QeL9piH7fugy5+PCijPV8wYrPN75LPVuOztpC+Xt8P5pruoV0qGQOlu76U
e/NYo/G+MPgplYJ1ckVYhD9gVi8+jsxQpPRPCgVTHdA6UI4qfhXl1zhaxYMgyXIl6pAPTdhkdLgK
P6FxX4j0IEsQuFYn08/GngNbJgANRjiE2cbWjm/816qgSfNO4V/FFjGfF78kY/7bAoV2ngF3Y7RQ
2vXGxo916O4zyQjptPEuZqPRnHPOtSJhcXr9hXKG2onhJPkJNrEvSQGE17CQISquPwe0Q9dC5hdC
oek9G2zoY8AZkViyJIBt4SeZRTX2O9aIZyfh+l/1Fk6py0u1q5QnvBulfmKGmJxqGO8Q4G8IuSFi
0ad1kXXltfjT1QbZpjMePt04Q7nTiaXgozhBQ+oCZbKvGSzZSVCJF6tPPvuLB2YSEs/vhAxLRA2L
MsEYQk1noM5AvY+VZs5YWLSp4HWeaFQVmx8WLbgVv16WHOnVTUgO2xs+i3LDave6Hiwg3MFR0Z4o
K0JJG/40S9v/GhP/xWyVl+EPQiIIoYioxkoL4dLtyIDd3tTzbtXn6wZHpLtMGEyP8LEdKjWWAGIy
UqcjUv14wdLhO+jXeREQhSaWJSXnFGz9NbeplkZX13QVicq98G8AD3Qo621/Lw9S3fFCnuf62Ihf
DsoT17HARoqMVyMWVsc7rbIZv83sUVQI8g/S9PS1E/z4kmbGl/K8WrAbUo5jMSDlQtBA/rs7092w
r0TFtXruU3rtkLP5p+datTRzKB35latNjh7H7ThD1Mk94/2vfCctbk9D+V1SU5+MsAaLA0pknY12
q0zHBYq1wcLV2DtIz3QhnDMfXr4+6egl2mB0FhxN6B04+w4ZHJn+KE3frS50DjQ/wJcXUOg9tUwJ
DbXq1rTOzYgFpogQYXkTNLSuEC6wnr/S7ZnO/NruHsI5s12Xixz+6FDKaGNf6rJ1Jdrr0QiQdm8+
rw39yj7e98Qx2kZ0eqSbHLqpVsjiQkfpoIOKwMTkSF9ys0ubP2S7yVI79/SRjHufoN0CUYr+Xa+2
LJjdmGYriJvxOYX4M10NeEdMsqnfmrqAVNaBEfvXx/PeKBHXZ9rnYKN92F8LGGNF66NVAhE+w9sj
tVhaWwnlum17qaEy4vrM3nnYFBYN9PLt181t8kVFoNys+mvNPKrQ6LnZUT+aoNY/JcwPLrIsfd8S
EJyumSigtpUmPf1oiOdmYRSMLF6d0CnFP7AWOFGb8x8BCcDSc9CbZ+bGlZLLnZUokd8zvBuZ/BC1
KPlv4BC03fFKJ4sJM2pvdxD52mSKQNB45QBfBB2lqNbgowscyi9XWW6NtF0QViQFZHKNE02q/scj
2muxQFSH14kr3VQ2tNnwtCkqgWYMMTNNBQddaE/f572RZwkrW6NF6/RqvCZGWCXPYuu8ERkPxbfv
B9RQWcWpkTxo0F8yF48kt6sUJ1a5c+gvVCwS7JVKyZ8sT/JeiR+1B6mqfFTET9QPFYt18W7pGGQB
XAP7iYue3fMGh6+xfrHOUNmyUGHQJiAOD9ZL/uPhDj1ZudC1sWbYHnIB+VPF7db9AwuLvJ7d0Em1
Iw1dwBdSJjcPRlLpcwzXPiIHM/QnyV/lX5E5y1yCOe32oh8D3+S6n3aKiI+/vjOlpmH5aV3Ll6u3
+1pJtTdEfYyEoU6BYWUUeEKDsuuE3Dr0+M3HeHUTOye4IMY1dtTnx5UQYunrtq2k4QGjOO5jJKrR
0rREnq4ztZizSNtqnQyOQu+PM7vPkoBh6xpZrXO4ou7I6ZksFe5f5rI8nPFxlT1H3dOGdXK0QApj
eRekd09TNzeTkEeO/gdlqKyronlSreXiWOKUgmdHPPfj6CwQ0BoGpzAGpEBrVJaD7OjMuSxRKDGe
ysHPw3y3OrcxaqKjQG/Og6cxnTUC00zvAPkKGSFx4RYj7dt9uC9gbgcj+b4aN3j9JBcUq6Ez324j
qURCFANcsHj4JNOaE4KUeUeQj63g1HGywjsFRdOMixzfmKxC0oKNZjicy0xirYJNFFKVK7e3sy1g
I2Qx5OBeR4bf94LEUWMIvPhvcDQSLmsGDJ41SbvL1FIm/UEqvVhawSwOj6JqD72XcphbTVSvB6Rf
THBMdA215X1DQaNwe8ro911g74eza8uvzBiBCh3KpgagFvYrU+3MojiTDGKt/Q7Juh6/heaUKMLD
iGAruGiY8jQvz0Rj7CZYybv05Z7zyJdZ08rRnb3ws1uO99/pcTZwFCTwaDk21gotSxOJqhyz/6Yd
oh30lwY8f97t1FfOLj/qlJK/z3ttQFI1RAGATfvt4Nc2yBkWxT3Xq8dwaHC3TV9Ek4cP0hLVNqB+
+P7eyJO7OoTlUoLW/sQR1LN2AN6fUnqp/JkJQyu9d1bemG/Nc4GuDOWR9+oaEy6cJDa8rRbHHNM9
M7M6VjGogmNa7JXvyMr1pEJ6mjnxJ6weWru+CIYLw+2keR9nHqYefVKpW6roxDg4nBj3VGgQcUJA
ZGtrW6wD4EJEE1X99z7nrmiewwy+poqBPodMkwU7y8bGiFeWR9J6QbgJyur6pz1NMiGJ/qjzlUxl
PRYL6OUzMGfnrgOdvMnkZ3eMq40TiQJlv9nsKjSCsWgJwvrFutFG0P2l0AgmdzTigfs7NZl4dj5j
O6u8Ph2u7f910j0tNhjyYZYa4uV8tTYGhbCCXTOnaFav3fSxpruwwFHVkCskQwUK6hv3zkFthB2j
BBXJuXiyPnqgEjTIvGqw+BJfGBYyGEnbHtEJeD3onaofHYDuCiCu6bXIjsNxsFNvVGkFGcy6KcbL
qvyXo9VXBwlEmJtEjb3edkbE6d8I2Pc0wMJz2tOm/9gjYQ+t+Y3kXfrAJJXZeDH7GgKCWLsxfakW
l0+KzasomceXEU/AjGjRmruow12wphIefsewLqU7OGtzcKlzD+AZMn+0hN8/gi9Q7UGD7B3GD4Ug
1x8zg2YlgWY0kAr0CipsE1VhEKieFSGdT9r+/iC2YSAWMY9o8Upy2hUhoMvG91vn0i52TnN0wOtb
nCPaXNH44uwAQC3kMqCM0L7NZGvsUXx1KbprZg2WVKsAcfqPoNvIHwVT68fFcWCXdSXm2hUy1nvE
zJx6l6g/b5ItO+bLu3nz74iCI8p4K+o/TtOhPLkxO0ohPax8PqT6owyI7kSmsRK0ZdaDXuv3QEen
BPMzd5ulR6hwxzi1BTH2Keb7sdKGSEQtwnK9r0yIlDyNQlwoZOPPz4ITnFmyffitQ3ezeojUmbJz
QsEczpdehGNrQHEeiTE5IvBOv8De+kHmH+5eaWz/Guzy4M6y1ybVPg4d7z84zanvMLJ7yt7ld6tl
AY7BMNxBTJDBTjZrXZ4iSf8q6cp4jYv5unKjxN6Ew7sQTylsAVwc3fNBEO5+F3Jtkoqy90PBch5F
A6h3v4eFR8aF4SQ2ePHR4KVvbymlisWEi9c+7jbanVrMqenrIqsmKHlYuweoFxJhS/7/ZchK8WA0
hS/q/DQcL6FUC8obBf/2lAA+Ls9xzDq3cJtB/LxLIdNSjkOa6rCt5iR8XViiTxIZBkB5OFjrG0Zs
unv5RpXHsK8yjNx4I189BnGQxvKNpAppwkpglmI9/duejhQiF+KHwcAatco1s5Iy+Zgo5SOLcolx
2hu3kcvOcZYpwAwjU0ALfo0jv7VbpNwFbc4U9h4AraM1zgW+ZUIdl+f1iEwIttVlDr+BhgmlbHdN
JFzNxslV3ZToKz2WLaaRGAcahGxv4SOj6l5NnxElCCDWgNgJ3oLQiSnHulQADPBK27Kxi5cEVdId
W0vciowhKLHuJrTGa25HQA3AXuA2oDZnJaNHFmATjwxDl7pKeuyhYB3K1ZStfLXx9u4mVLMZaYAD
3FlgR9UL2l5EkR+Q2r0MG0bR1M/PWQ2VS/ARWssLM7V52d56vcqBrfKCYwSNysfjm7wdCNv2BJt3
s/aj7/qVXP2qzd1oG51GN36PB/r0DgwbnYWE00XcJH4nT+FwTnfaIR+LSUwf5CoZGF0KSc5gDWfT
5f9hqfYHfGyHPKOuksaTi3YMSjf77Rgu5ma3yZIw0V7tlh+bK3Ct3vrSLATQIgsxvkB1fn5M3e+t
V9HhIwexPZCMbaemQQmZw90UO8qbI4Et0N3mtoBkh6ZXwmrdrPt7Pj/iCvBlI6gQ3IwyhoY/jteI
B5RkalW7HAH/++uiW4ThhmzsoAXPZ5HTS7Xm3N5y13WMGzEOm3eFP8s1uF924ARmwP/+CAoyARDv
oPJbuLaOZfoLOSo1S+pyBU5oRIm8DqQy0ziwEJF+JgwOUh6UXrymWC1Uk6cn4YsLdST8c5M30gUG
eKRElJnxu2PWCuBA85IQfX5BEdLO6Kp/WqZA3Ly36LA+ljMp70Xv+zB5r9/0C5WcVdfapQpl/ACz
LCSEl519GFpuYgiOugnam7bCnenIn17HBIEWfXWT+7+XFfdhHbItQyiCdkspjBF7yoVYoWd3zYqd
C8rdrWzULVL1FjvbDVawU6AUlhEd36AZPJ6Wy7A0DPbZyhlQS39zM5KoDOT71po7FhG1chAuZCP/
zIeEv8SO6OYwAieJwe49rEwdCjNnSD2cBQByWGjV2KRgrwiQNqhawRDLQ+N8LLujdHWUOFPVDmVP
asFySnTKjkUDeY5SnkDN7jkcUfpFy32tXq3o4fWF2PHJ/HTjg2+Vq4bDCCE7r+Tiib3nsND8Spp8
/lP66A/oSzBUuFXJz8SlQHwJGGNXzPVlNGcVnV4NDcFWEFfg3IrIP6jQjGs5UQ/Gc0i5vuY1XHEp
jE/vG4BUSQ4NDvda/Zk7Rgy5/RROpZ4M/ixDqVGMx8ECKvmAQc+R9zCrGlhhzf90WOfC0QcVo6OT
v345KFF+FZGlIkdpzkk1DPwTpa7x9NB1W/kRn51EGaRl7XbisQoWAroe5aLtW5U7Z3vQZWN9TohR
Ott3NnYsa242uSAfXhvASNCGyTbD4W/un/Fqy47qN6u8PQlCsSO0pT2G9qDkO9UL4P7ATfIkyyXq
QK3/TEoz5p9ptUTCxMatynw3O31Xn1qlFElv2Eh4b8CGFHot7VvnOXs0fiHdJM9SW1ZxvGf1YBFZ
bZyypNQcDzP58uv1QYEKXC206dk1pf6k4cLvQCC5q4hk1YqK78G4HRX4aoYW+2Gtm5qgCdn/HkDG
g5P4QEVN6caarOpQwkE5mM95zWPF6gGNOCU0ENK0XumdkkN3sCd+Jb3xnswfiWVFn+BY2ShkLunL
hmvkrg2ArJe9poZfng4GvEzTIRaevkqXD4Y/kwFkrTXwYy5eMjp5QYkeHy4kfOOSKuAeKtq7oICY
msqaJhZ0AtT5r8l1t+7owtpIUQRB+OPRhTIC2DSxJoUDji3SSs3jy4o5B+eLi2Bn5ej2VLfa58X6
pEqm67htclDOdjRyeL5IF07OAipa3jHiUU5EEcOrQQnIqfPzPRC6d7qdAmXGbqQCBfZ/1v5EHQjZ
720oXlKXtguvsTD1VlsXhfXV6vz+Ae09eDcPnx4lyhVM3D1MCkc1bTcWpSjhrLy+0UACCgLPJUHT
wuArrEXNZidGnCMemQiRjZFZSa92ilrK/Mr39DXO+spYvsM1ihC9j8ZAqizYBhtCfdVaqRoAckQc
dUeJuFf7ImrP0tcPmljFBG5fRBV20qHN/PNIqyboBvo45qRpfXGrz6klJPw2C6icNcFsVzb1OcPU
o3ik7QtSDYcnjlW4XeCk7fdNvt4tES17cv32QeMQ0PETkW+D69cUwksBXo/EB0/Z0tnDCu080rmD
WD63Pef+IzN57+Ylqjltu2S0YY+v5szlduQrHXjpIqP5gOYWDfPEzvFqotz5RWZNdKgdSHExAeHj
zPzMwwasj2rZgfUW+T/czE8Ikdv/U7WSgJbCGnytEgO7wFHJpJ+1qu5mqggIvViANAe91rnipMoA
NUX16y1gw3nDxTZ96UZN9id6UMTkQr0ArRJw0kxj4oyWK0BaeOVFZCWgll1akSUriqt281lYocAc
g+F0zpGnM8qWAfwZarXatb7dlWzYcGoB/TUY5CBS17vWVrusJvjBCGDKwG2iVmFKRJHfKOnr48Ro
Ogd2XCYBwZwWRb2KUsgMf/XosXAXVGcg5JSR8W1Y3sl3ZPxQG2zP+n4okkdVPlk6G1dj7Lm6DH+c
HrHy+6MZ996WpEtitkdj/Kx6HmGwZoKuaNaFNgQ0vaoDy73h+vLNNXQq9uI5IjDtgXrn8YuIvP6K
MYcpyJPNa4u3OVDFLkaRnygxwL8pIGtBemvy0m6CKO6NeNMbPAqXYCVZH5n8ED21XY+Usop+uPUc
qd95w6Ww1r16RA/pUjeIyESdAnoRz8zG+NLtuJVur2WKRokixUXU85Mu3rXcraLQRkPcOCz50VLx
hbPJ1omspXLRRfb4ezmfk8sqlCUyPj7cu50664ugaiuHo9TrjiXOZq9SKXV6HdcfSdt7RBEDSMVp
9n0+c6G/gCFBuA1YOmpPoQnIg22mMeN/YDqOtC9jHlqW0yTuK740AYsNmCXfurUIAeYJyOOKbe2H
M+6iAC5Wlf+umJCiab+CvOU3gTDJm2ley8wOCjLBNiLBtTJYwQepJQCaZdBiHHMu3Lm000TxEM3a
uNTsqlqvKiBvMQgJevJuzdzhphfSHrWyhol2KVFFeWgxueDviGQMF4QF9LMVpai95WjXFMDdwu86
4125/etcBi1B9X0N66Ck2ApgqMENdnhNEbfNiMeishIWC14bt2K50HDALEMSFNd3p8Ksl+fJ+OuW
Q7Sf8DxsL3PdbXYsmwr7m6hR6R9ihkgeFT44GnqsyTKr+PA0eFpitR/7iYIzqBr99QIfOM8vwrEO
yf6FsU6RQpF8disOiSkvWogbOCCU4DUBtpQfusI69puFT0dzVaC6agOdxkfPlSPySO5enmiJf8f1
C17NlERKFZqzUdoHcOB8RPaZLlOiUJWyxtFroSmRvBhCqTKRoqTHWXGywyj2rzyeKTWEAiB3k2VZ
tYairihQgysMVYoZd8rDqPdzaBKqeHy9z/EtEQbMUUoCtez0/jTfK9gcoINuZm/8MQ8qOdqWEd0t
T03JLQXRt3BwAIiR2AC5fiUxGMTQTP8rgqLJ2gDIDPHHeczD6udB1OsqENssJE9wISfqSs90R0Ov
j4PtfuBfv3u4jCAUZndF0iksGrfKVZLPuuiG1b4F2lIIdfICk1+wIxtt+GMl+XkO39wFHsN1fq3r
3dLkkyKvsvS070CzOYvP5/nfjOGVuqoXHtKwWp/SxThhy1OgJ4rH9JLzAaU+YgGOpprIyNjODpsT
ii1z9gWRNoJUDqAGeCkqI7s/LPIVQkihoI2AFXjX2NZcbOE3X9J4NOxuINuzpi/hL0wAKqwRMsYu
zPQfq2Ym0I3CEzhKGyUh+pudWDGAWdV4C5kqNe9DtNSWhMRMnRuJSiC0LTDtt+hOFUzJzh7hNP+P
JzFcpKgqJ2wBLm/Bqqule5rtpxwMKG/G4Vz3gkqH57oVgL9m0EiH+LR5VgzC9x9EeUeIx3cYr2ko
y9MoW/UPyBANBMbDZ0PKZgjX6bDxNPKZwXxmXQ4kTS2DQimz+Bqq2rtZT8pqlIWPsiNHwCb0hlrT
CJjpGNweuwpHTR0rKrC4oMhbpqPymgyDVkaChyHp7DlVhiRAb9UW+Nw8VWQ8O18e1A46oryjAqiB
+3rHoRXCj/ebjE0kZcSb4S9G72G533yOTgkQgKSD7gKNj9CsJJPk6G7/AxxzZAiuvZDQ6WHJegPC
J5qZoUMbuZLmp11EiOhRkQhiGXK0B3Nc9GO3mcZyGQY2JBxVTBH8F76sthPLrnRZo60WGmR0Hzsd
2Wt8tleZyZjMw4+8haoUB4k0sBnR2mwguegLrJOjWCP8mblXBKDGU3YwjO1kiPxMMrCBob8BBUNt
GBB2ruVp5xkMyjC+g90RjOJ6yU68Ljm30/KWrrzzgeQ5oTCplbHd7lJ0d5fc4zbzsFheKdFkTtul
XzbuI37s6XctQL8zMTvsnKiq6POQf8iSKKzQkts3jW90ArRR9TSDnDygyhZHuS+5hGSz8djVhbih
PqF+x889zVW2KQYXhphfFzqF40qshYwfJyT/YQWN361YI3N2Z46G8X4Ggr/nxk+EvZsY6M5Hs0cX
a6DGDoO72F6Y3hqAEJqDB6+lsOBr2LcfRW9W2bvXUmpmH0Wh4SNEkBsEePcuBq3ytb3UABfp3kw8
xnhQllx4zg53joRpEMy8JFeJ6Vz8G3L+90oH/nrqqqvKbI2xbHFaEejR5TdM+Wxe02Uk6CC4kx7w
xEIWZ8HO98pD9Iy0FPPdvYET/RfxTbnNv3Dbdoif79kuTjlt8VnZh5Yz4pwuNSaGenqF110nFxxd
Xya39cJ6WUciPqVJSuoGLNAPikQLmW0ouqk0/PXExlczpeIHVz9y2/fSxwOp/9wt+5cJ4L7QZr99
Q3I1KwF534T3eynbC0uZRPdDSHJU+YzmOWArD9I1ljEKqQ0CK1ukwQLX+nW5ftnCCbHJphDVVMGn
7HpJ1keYKB/cQ8f+8khug5/SIZtA5nkVccI0ETPOcIsy5N+P24Xwj94AFrNZmi84e8AGnmWAycjj
Stm72bgZbjqNMS+yBOfH/yN9ZpA6ADLQTlxhzl2kneQXv3sSH8QM4TCzrdd+sRE0bo/QOBAiklq2
J7THkS/koMTpmNAbuM0jxJeCYsCKMAeRXAwX1IAAvh1lgT5mUGMMV/YuqahI0abcmNeSfUcUXFL5
F+1FsoBNFbLOVT71HK2tn7HyDzmILCS7Qz2knkRv5c2APwgxVvmQ+MbSIwAxJ2wcXIKLNEamKTyN
ut+prOlPT+6u389wYQOSHNyvP1wFKFB1e89sLExmN8O+HiFpAVuJFslI84fqlYir/I1WQ+ZqMZiy
kLAx+0GIoOOjBKvXE3T8fDB5Tn+wRQML4OR6woEJcrobVshJJYZOL2EknleNiZQOQyeCfPY6eDqT
z7tcP7cOqg+8r47wHJ/WUVzMooAQuocBQVF774XVQ1fAVDrvpRUss70DeJE+k3uefSN3vTiIaLw+
VK6VoPkNIClycomRhV+EuU811T33T4bFKwd+i002XneiWn9cMTybAGe0DH/s77zFnxk8i5z7P6vD
WsTM+VIf7BJQ5OcpjJo9JtvnE/T8+3NXQJU2LK0NhCuqWMPseR4us+48kdSnOlhiOpbvCm1NiXM/
jGL+D2b16JLkZVDR/6R8hSh7XsjrvjpuOIqB2qs7l3MJZRras8r67ZtsMnXsCamUujfKx1C/qiko
mYYatoJFEjXFHO4ARDDUL5m/KKeiEJkbJHtQa+NHBsxjM7ItiGjnqKC8kUlWJ9Z5gBQuseSvxEkH
4SruL5RDZR/wIYi7tCHiQCeW7LOvOp346UdTwY+znSeecSyMtXIbh/UZuPOFAafHe7PqeQe4P7Y+
mU3GwDEnEU8coh6BZaJn5vvwAiuZrHyb7zctNz9mwHd4VHrfLGnBDFPP0gR6qHLhG+MvcWQ7TdE4
K/GS8AOr7jJuMm5IFdoPNpoN8fJtdixMTMuBoDmn8Ig1Jt1R6rc1Yz9/f4WHLZ6rzjQp1MFuUDqK
N6OMqZ3HWE+JZkF3/jrca2I1+tjscG4jxjxhqbEe+Y4NDJkQ80/WG4ctM33kzbs9x6ql0mIJzYRp
8Jrpp2WwjvrzgurBUzyVjN5gvhVteTKgy71GkBPGUhOdocuMZuOJaHpRWYN5K3mHApp4FkEAEZy8
U94oPXj6Ws7FTPSRkMP7RFINyM++mTcW0qRtebvak9vNc08TG9I+P2NmYcBSb/tDDsrp7UkeCqmg
1WAiYfMS4nF9w6B318gyT881x662M6Gh0te8LalISZZrrPOsd8IjJIZVIAHk32q6YTZXt2ICWAqW
o2tNpLg+ZgCl71/sG/l4CIDWg89VRrnigoTzpQ1ssQMk3XIQo9IeVRels+s8E71koji8lD8Q4o+c
wQSW80QwYCrcNN7axuqD51NxXMxFgysSOqswtqa4M8eckgFzbQO6x/0l2l2IhpBirM0UX4M0IN6o
5elKfpxKVvgJTE37814jta+gihFeIZc3RVmnx1hyZ/v9c+HOrLpSLLAtQWdMeuuUMhBWw4chlazx
rPvg/mtTS4do7ioAfg0bIIoqwiFcQmRuMgHJUVuYMtMEiSiv2WU6XJ1DzBhK37FjWqmk0N50iT/m
pYfJv90dkHmECPyPrn59G0z+X5C5LaMJVoY6TVqr/alNXD/R66RCDzkKZgP063qAzmLRVk4znEkD
ItT+XsZAR6oQC+hgIJ3/4aXnq+nB3ulzqWIL2AC6DPNBrIf/CFB+WtX3xfVBqlucnvGbvJeE+xYM
5XgQQT88EFQTi+StdqljeOwpdClzCSYjF1vvT8uq9Pq4j31j5fiCq9oBSRQmkpYGbprofvz8DzM9
CcEp8VLQl43zDPavjavJHVu1Q2muCborItentR3lsRcpHLCRxhQ2SXOX5oRqycc4R7SQtOgLHy/Q
xtcplZ0LKMaPd21Pen318RFlrclGtiqnPH8Hn/RFfIWevHIHZc2kOe9yKLg+4czRf0exwE9V5HTw
XZJfq67dm7MZvSs81WZvKvAe2A1ZTBxW8CrKtG/kQK6kDKnO3+e0IR/pCgPLAwg4YrkJmBE4FT8u
tNP6glo5AV0aIiI0hz9Ew+Ro6FIPb8A6cQ1OtutxXKek7/tg8QtAJ35d4JiC5dsw08NSMJEgVwFz
knM5fGzdIKXMoKuZmUSSSKU+2AZ7+Q2dNtHBaa3AEudLFoEQ58qXIvWd5Vg8F5eBL+IIAG7AKoqt
18RPBTxe60tTOOaXX2w85/PJC7knBNoHuW6LwK7+n71tfbe6kPsWaEkBy3msEfrH1pdNpm70QXKP
n/0mCzOaq/4SwrevGM9eYfAvr9BFNpdKORA8z/cmL9aIzLD5qGatYbT92i5b7fBSA2rcza8ffNKc
be2mjxD67XY80U0xH1IgvXhDJHvfJyzgbw4L2/zMnhGrkFu+WbFUFwqulx3x1qdnVil0CbSkzO5g
Fd6Sq4R+tSaSMcuF5nPAy/VSi2pFl9NDlSRZCl4JnVBxHfq4NpngEu+qD8NTlBbKF9LGSW4zrMne
J08hiS9kqM2gzK7QCh4Qb3cwy2Mx3IvsJSRFE/SCIxtMBYyYBt3PRLK8LE8jIuIa6hq9SlgH6mPP
+WpzSIw808SSFr0ZqM6+4XQkpk3WXsg8HFKWD7KueQzcbZ7JrOyy+bVC0tUqx/i3u8CfFVt1cRs6
i9fhKEQJ/pde24MgttFSjeP11CbM879MHPs9rZv7Ot8KyRadPE4P0NPpRrC8csK1Vj0nFnI/in12
3hQMY2KpngvGcSVJT899j4EpsCUBXmte1CXp41tPkB4V9A2ZEhIMYPtTDcmt4XXgiJzz/RVJJMIn
x/Ta8NqL6gIRqUfC7vP0/GVL9G1fekzQ9nQDrOfL1GWKcdtW9FcxK/UJjfASM0hd1ZRgDHnPzqR+
WxkZvXl2+mNor2INLWpVHlBmyDHBEZPsIP0oZI2dC9mw5+zajYrErP5JIQlVgFeFppxPHOtfZWZs
g2JO7WftmUmFeI4WbUCOzZZv43mTHAfgHMqlGWrNdL9lLdD9OWcynKxIgEOoBtQHH1AUgfqkkYVT
e6eOubS3FR+rbpLAwh1FcaMsKGv/7Dtgf1sJnyOGMky752nQxzKAcjS8pADgJJ3ES8O9TehI58O4
om4eWw4NMwM8QTGUlQ9jHclfrH0nZP3OWXz+sEzyBsA50pLQNDlaiwTx2t3mCc1g1eeXFqCAMsI/
KcA+wCaZ3af7oPMkZtnNh83K/wi6FtnmzgPhirqu6N2YnWRf9nEThEujt2rI25xt0VtiRQ8DJs3B
I98LVkkHCICO40XzM1vwEbf4WIu3xUk0BeqBSLorUo5cpNctw4utx7Vqy+tKRsYX4O5QBZXQuyWv
eOvxHgb/JPx+RU5AzgwDnkn4cZ0Mk0zqCdIrh76bbLCrMXa/VhEpLtMXBG1aexph3KLfu+Yxllpc
QbM3gKEcI9mVWbrXfTga8CuzIU62oXOnHOgvZg/7MxsPTAsFtEteC+w4km7NzUY9Gf0+naDmG6a0
Q4EKrPqTSCfZWioTkPtlESWRZJoreRcqZ2AtFek2bwl0GAS3K+Npdngg0DL4OXKX1GBloJf7FaRt
yJ3LUrGtqHvXSJ/xmFHKbNCgnzF5knkToTS+gGr0xubPkhcTszXGJpvqsmuxmCGJY7HFrywmFpzM
s1hXkQtFcoS0q+u46h/Cccg3KjJqmv26w0mOlkA99xd0cuxJaVd5LeAFM0g8k+LOnpGP2/UiEuJH
MtBW90vsFrXRrq5jTPxuSGpmlM0w25jU9HmB3KAkiNEcU5lymL0o/ZN3w8Ob5Wngx4vdN1Tn5Eot
26IONFTAboktbE3qj5zIU38TqRelLv7cWjWSbK/XU0qCJ8x1KqwkC14ZYp8N2pm4JCz6IsefPW7E
uCESuLxrJO8Wm2s67+Hgd/Ql9XJSqzMfW+Sbc8/f8/3OaB5l8yLBzog7Wn0mPSzB+fEGjOhK1PVd
zED3MhY5WGUaeSa/rQtUyf8CpxzpAVOosCxLGSDTa/Cna1aPc/suEXvN+csydVySgzzw9Po3oSMy
GjIWSeR2wVU9C6IvBnptEZ7bGETrVWAzsI/3bkz2mQ2QvfW0XJWtho0ahkIPYTVLirwcUCnZeGix
AQxWtAxG7xb2ZfaI7PMP0vD1Tf71vJ+iw7eSAgC0t4n5yP8mI2QRgoO6AUwYcb6to70e5YcTXjJD
wqnXwlphw8D6+QorFOU1UTqLFxQe1WJc2a1M1UgMluYTIbp+M1HAiQSRtAwQPKk4x59tkJzYVAbf
hY26BYltFWkdvm4XqMlOpstprel6bU53dh2DWuwXhW6w9nS+rv+B27O49i+LgEWCg7/J4c1EtsHf
GENheq1/2n0bCCCsox6div20YKnScUK28er1SRp0sH0sA0V8CHMJrQk1PKfr1ZToIkP8kOWmH9fA
tLX0UO+vxMjoxyLkydD+8MpVnifX/eNEO6efoGy5ybunyW8XFjiRPIkiPaR8+lZn0em4FlQnBTQQ
En1YoMR5HaCE5ZyDHwPe4bZTKvGuvujuIE4eXBpwfLDbwt/tAl9ABWld11/PUIIgFUFXz7cxdc1j
ctOIktQbAGTfxqWasSxT6dAtlhZu6UIhB7rgYhfRWok6bfVug/ACViuQd2BS/RL7eZJ8jTZE1AFe
bG9ZgReQZKkPDtHrVdV1XY/0vGfLVhSZ3LmvOKvVsNsbr6/EL2nqVjjrijeGO4zr85qlaTCL/HcH
Ki3BL2kSzCXipDbw8tXNPl6jSEQHO/ErhD8gBuF3uIdX+dkvPl5LgqdSvijxONI4mniTfP8yGNVF
h1rcW4aq5ZDPZBFCC9dHJmaG2Drn/ti+KTfdR/Xj6ZrDrutgp4VQdIG0TPs5DZ+GZerFkZg+Tvwd
/QNsEXO7ryCzh7wAQpL+5pJM5meJhAIK7WlhHogsy46PHRPlPYk6Pxsm2ggUK6crz1V2IbRCLYja
LFsreNndDIpvDYxlp+uutD7yXIgQnHwhwsixvreVLwnO7ppjXONdLN6wjJMluFCGUwb7qDn0vjpX
+UUJm4froXKJJyeyP8CFi4jJO53mtLXsJxmxwaRHuWl8xXSuWaABkUcfiQmURFynHyvu+vqDiwdg
r9K/BlReCpHl1ZZOwdmun7SOqTdVQOKyufOdldxTlSVeNwkVbaokDKBzgWQWgKn7P8MfXsvvr9Wa
+QQITwFzyzRcvEoHsYut6vFJ66kGGHDR2lrY/H6+GjcGr2uuTMcJQAGkEqPM1IGQdrYcAGE9haBl
TsfeNP0sGfP0+1Qw8rdmRSLFLdx2AD8gds3Z5QyJ/HNG9mzrFhKG6ZH/Aa2fTyHmvmCC1K3ZvFvx
AqvEGOc4wWgeQ1ufBYCMnxkNIRisLly9VPFOQ3SSDRDn4BuSQ8goZCV22lavD5by3gSnLKymJxKp
4Fd8zmm0dnhX1Mr6MimXFYw6w61+LoWl1V0hXyq6klU7dhx0BUCUsYJu8gvLUtkxQ+RkxV6juTSF
NGm52CrbsNkT1H3Utpw8Xp5/Z0/zfuU2MiaQVeyPZprCqJQZIyntAvENrFWMeGR+Ry9oSPXnqs0u
4ZShz3UjE9dRPWTHZARvH4UsDKzOnfWA4iWeEEAxilhHZR5dz2ASwAQLeojqzkQNlf42m31bLel2
CzITDKcCtsCqWmfM8LG9kQptB6Egv1BaPqcRnCfhp6QzBmUNkQHL0lsU25y2rY9RpElR7nyaM2Iq
jpoju8HPqZq0fkotoxGMr+5HHOMd51xCiVdKaVDrw1dsDIcDoZ3oyLRQJDW+bmk+CGq2K1ZmD8jb
NtseQpKwqJcM+uawghOqjs6YcfCYFgANh7T1SE0zOk2qClnicqAReFGn2TOjMR9ojalpYusfYTXK
9s2z93oVWNf14hl35KiuJGjJ9bhkCaUH9NzNFkrqEzldlyH51sWjhv78qRTuXom31XAAzcsaPVgA
m68FamgnYIEbH67UdoLGukYYCJIrYTQBd8zdEMGagw9n8UVoKtfAZKnz5Bv51HmEWC68v4u7MAVJ
Hm/jU7xLN1ZHNMAfxsLjeHyGZO3zaz5JifLXYl24klkLVuHdDCamxzkZ5HgRgJT2owie8pdUXuls
tOcd8ezbk0qDsrIlQlz7XMov+NHFQv3EVBq/OL0kBKzQ6prOiLPFE2l31RnXMeCGXpJc/c254wF1
cB3sjHD2XPdtNAZC9T0nmyox5wQkUYPrB8U9x6JmvqFk6zQAuJTNPtzQbvRq9v7OFvozdJIpjjZM
edsaNRASXXeDzw++pMnz2WL5xyz/lbbtNt6ggIX6MpvL4ZsuwjW/ktyD8iea4U0hj1ja4eRIJYEu
lXcujjYjsNaGeXspW1aRIskGOCTqYYRQC5Kc9PxD8Zuwsj6jPvq6EnPZqTQEgcXTM7XYRhzt+fUA
Rcq8bR0KzaqpNLKa31BP56q+/FPNdlUhj1v17S5YTt0B5VwklDf+x44I2obzv85LNQhkpOpl0br/
yMKLH1F5Nh05MYQHossn8zsZ/lrCWqSBG3hGLCCCINd+Zfg4gcnhdefRbvJUGoW+DTLaxzz7IYMs
w5WhVJtd1hoQcnRdZxVvGLXcgDQvhE+d0OnNbp6zmkOXgJ93Md0dVP12vFzogRNxI3apdXbifoH0
vbEQbvKc5dg30XymQWldqJ2wSlaqX/yh2hLouPK6m2VxatXHbqgdpgfpDqsUlX+wICc7z7c/LKP7
9zmZuRoNkPo8zlnqwB6apo6t2SCbNl5u/cIrBBnyApIrePJ8yl1hJCnp5JjrA0ejlkyg7gQZI5Xe
FXorX0s4GzMW5CyKOvMqJQ8/MvaoTZ47cbPLLDvIwHBSyNKO8vbPvs0KwRpZIHN/ywi2Vem3qM+s
ZSGzNJVDAHj59K8vLtviNlF5qsT2A6IsFVOPwLS1Wooh/XTdFK8tRIqUmXGPOpPu91JnKPklZlyK
qcDV3qT7EPb19kBrPLojPf8uzcU7U4DE2Sg6c8LdamNzjhQD2k8r9ikDuabinqunBlu8bwJjHSAA
gn1XxKV1+Uv86uFXNC0lWBdotsKUHDRuwwRK0uKrVGZP2fAwVhBYNy32jMDOMASiYNVqond4f+1J
Y16zFq5u7xu4YUpXjyi+8fTiYbvDJTAHo8pd6n7j2935K/zS6PO1cyeZkYeadWBHU7EM4ffLiq2i
5u3dM7RT0Q3VQkIh+wdloWYclfWZ5RGxWR8lFVe3Zo9E7OjdzzYxywJdkvqrCWthU+8jEedsHvQT
Ho0eBhcH8GVwjczj8lxYVOP6fq/OFLEZkd3nfr+6PeeTm31OjKO8el867pW4klxgVqdhUaeKkzeP
ACxYiJj6gz2MKmsemt4s7uIgAWncCSNT7aWhazowmsLX5QMacZeBkVzmO+YqmwbsP5Fu22LiM8LF
K+GnK7hdW2kFHOA25OtgmS0gYKNNrA4vPljL2CDxI+kmiFMgEf8hA7klVa9moMpzzioT68Col5J8
jvmDaWxYe7EqA0xfvoxtB+sY2HC7195NNdbl1dKTujaBjTow6VC1aOY4gMmerG+Alpz5JwVxbSGX
6svYrbrGMDRNkrjDlxgiI3TeVASBZz4YVceDGZMhdjBljL/MlJPJrQxQcoSAlCYphQeRCIWiZ83d
ySzpBSa6JtkSrVW5Y/5osmflqsdONEos2zERlcumFEjoartahfVp95SG1fqdXTAsjAcqBDqt10S4
mJW7HATe4SMQ7OeOGzpp5/1eGzjD5IT7vWbyigOhhVFj+tA+ay6NdWNMZskaEVN/CQKC92QQZDKN
ZPOqZRhGBq6crBVgXgabSAziLEKgNOm/kXBuqK7d/FQOnxjPYHPkiXzVqCA+SgERYx4JwYhZ+egZ
1b+NkGzUCn3m8w1HWdP90mC0omE4Jbyj1YaCzyRUDmLoJg8ZIyM17mIJ94jrm0xvcIUTO6VofhTp
Dl/lvOwYBr5WA4YShk/Lvw92Ua6yWE7CETeYxyjdpOq/Vhs5Vg29C8z55PaKNXZUL2R3+743/m8K
Fg3NXBpxEZwBZEYoIGm5MOyeg0TFsTcMRY6uFoT0FQzu6KDGiAgCD+DJw2N1GDsdBYO0QXVEY5ud
0ZOD7XxWoDlhkhsCfHbbcurJ6tcoFLyFHVQUj/p1Lqb6YBpOjMbKQoC2k08fVYtRhAH6i5cNCkAJ
kmNRrxjQXl1QYsiIByNvreqncDZt3iAWEmkzinX1qxQKXNuuatfCPdyX8dv84npwgMOUTTfKV2J7
wBfVUsNfoDXTf3oRWBbMJdyj81JPKVTniMM57oANRiuJw+EhyejYQWKTAJs/7obC1uqFTANdj+Mf
SinC+HPCZLNEa1vSa9jy6LkFuyRz32fhosRjyi1Zl3D2dgrr0RlyZ7syDxHC9eyiFtzHR3Hc+/Zu
MJ0eHARmmSxnuvcakzuhlGRGIDMXJhaGqGhvKfrl0lCggAixkv4PcEShDsmavZLnqEiL5FtixKSb
4hr1tgSuq8nEtju7HY5Skxv5DvBspPs4JjFUwdxpCmPMN01Exl7uolETh9CaEvJ2P/v+7La3PGna
YNLKxwdsyejEDBiv+x+8sW/M804/1CsIBAQfDrNdh1sqZ9F38+zRys80JlP9pmfYfiygzt4dIBzB
SpR9IXhHIuDeC+UfgVyoLZjPZBeLT8FiZHp2LzjU+wzpi3BjO7gi8GeC4kYuDLOAGaDCK3GIAm4l
8wUYz0s3v3DInArsWdivL6TiQwG94RgXfj1FlNgJ2KCj1opYqOHJfUyYPCzaGibFm+e+z+JgyNdM
VCN/e/CRwAbCmwPYn/fnXBovrgVGxbAZAdu3xAqRG8GYgI6W5OBtcEcUHe2GIeVJNMshVpDbySnS
WSNJ2hYJ2y10RcVw2QtxJB00QVcBahqiJmI8uoJEzCQhZyJSgYkKKbaZoLxxQ4ZfuDX/wyV8vhTC
xFIAxucR4oB+9uyj1SArswy4UW53cs4Op4p2F7TIMbVjUDk8HhPDdCQgBDrK9BF4F4EjUtfpK3S3
rJX1wLTcDe+Bq1tn+wITpfNbGeGwLH/0SD6SXNYX8K9qwgBh2MNMFE37jS0C/IkHOKP9a8NxTZ0O
8/iKtDExxXJ+NOTVf+SYzmTX5hGjdm0gmNPTm2YYCvmQsmRpKv9tss4iTxEelIeMXTQ51rc94F0h
WZZynVufiBbovphDWhv6EYxUaWfvlsaz2BBKmjZuMln2anckxcYDO/zhyiEDDLP//yvlYm1R1Lel
4bDBmsd5NMBlKCyBWNhMBT50pUHa9jpdQD9uJyamv415jTpwdV/GsVCx1j7pWc/AsVG1cDNEh/EK
WNGYsY60cJ1jOr3oybx+ClGwlj4Mof1nXHcECDwnwTSDme3bWAPAC7eaVDD3X4HPjEAP2LXA3UCI
yY8loVhZseJ1jrvpBbqXXiOA2y5v29zG/+IllNplXKjvcTIf8EfphCkq/iF48EAerwxsufNyGxSm
JnD2RlKdIse7SW6ABv+SMqEnr1uetvvobmaLnsPsQi/FMPj1hVKQGmaOSuBjs1PD69l/2GQvH9Qw
+rcu5DaiX2JQeTRU/y7KBXUuYAvNNlAC3eDkhu2aAzSRXeN+j+AzrQY9H7ayRWUs45EJHtji/m0j
q57NlJMB4rCTJmEGKSl85emYYu4D4AoBk3bXyreAFXe1Okl1rVwnYg3UP5uJIgu5m6Fmdi0S2Ti0
xGuvsBndkUX7oqdG9aeaIqY7tAftCCy2cg2xp02IY/Qqo8X5r9O5uTkewZb9VDRerS/igrrscK3q
A5eF0sGnNiYOjYeEDSLyKjD9ogOahiDFsaT/WckTb6PKioGUn8zSpOPiIpnz2xAd54kUJ/hFusF0
BPWegRWyfkoUSfMYcM+sLAol0nQAtLCG3b4IxUcPwPzzYTM4Etp8ZJ2pi2a+ixs49LAh7wJP81b/
3u0FjYzu0Q/IUQfAhmpeQQC0miDYK5RQWdVRWp+6MmhMwgDGUPf8C1MV0PsPfuza2tmaKh96jdcP
V+3VPS6UPD7xaWOdBCUSlmc4eWcrMk2P3bZxrKw0Gm9S3+I5L5BQQjZdAALKS/cqrB4P8XrUAuuW
NLI87hCYbcxm9hf5PG9bS/k0i2xc8tz2+Ad6bs0QFD+AKlyjNPzsQmrPmEc0SCKVZKFwHQn5usvb
d2B88IBo7Ym2GXlRg9fgQrw88vmkaplLLuyQdN6PT1Y/DVesn3nWqydluI++V/az8/eYf6Vce2rb
ufhQqFee1Dl62vzlYIjj9wvRfwnOm6KR0xPLAmpTT6xbnr3Cro95msMliWRpudg8I+4MEc9LWeIS
t4HSLpVhPs8l7cJqc5oou0GDy/UGNlQtw89wKNeAmzl1kfvxrsbWIBBUIDDlYKIiVrwEGEUoQ9mN
rAW6F87ji3ZFoXmdBwBrpcNMzpSosuRcFEBVwAGWH9GRdxkh8Q0gB2X2QVy2Dg+nFTkptScgb0CU
fBTPtd7mbBpy4qL94IKHawNbh7K/2izYUI1m8VxOVvv+9kID9+bKmFTnAfvWZmGsplmOJqcVegzV
bGss01ALfODLUesOIm1AnbPcAbrX2TsGPIMa3KqWt323ws7FheDVaiB/9oJiDs09EQDmshMUzk0g
o09x4m/b/gHbKtJVjB96Oay10f8JSfc8RbLKg0HExUYUCjgWWhUpjss2ujoXHCjOOECUlIJnrkx5
xfouQcS82vz5tOW+sMt59a0vc46AWBTC/6Xz4GUQXFPImUV/G/zl8joKfffWbDjIS5YtdUPajrNz
p5EUO3cQR4FkfGK3yIL14UKxYJMGashr9SNad9J+7ABRDo13UahuS0EcV6XabllAZgVeS/Zyog0T
Y5HE4uGQ4Ou5lEUFybpLPz0jhJldEeLfOy7Nj7bK2qlJpiChEGvBR4O45i4NBapa28JCcLAu/lxf
8njlJJ3+0BnJs9VimqErQ1FfSdXVGkfdtl08vlZl/uUv5jxZHEfrhnANAiPwrtJJ57ZEFTksG6VG
iHh3rl7yBmFckF84eAzSZv83Ysa61wKYjFXjwCEPsOzuaYj0WCZT+0A7swCgqKBRZe9VWMu9VI4q
KTGx7frQ3zypruiplkEPmK5MiztOF1S5ykbE8AjZlr9/aCwT6LKjv3Ou2YtsBUVJeM5eqnnBpDcz
ME2hZwI9wddAYDRhmQuByspsmOwG7g4e+UV0iNJ9yGWdXG9cVA60M/6jKkbDBzHAYK0TuGRb7QNe
qo9LTHhbGPxjcE8UMunYFBbOJsKJ3xEgtR7I3FGk4VvwoOOI52LFDT7xEuIK4etab8QfXkZ6STB1
lV3sCpd8poUx6YwUOGx61huZZhFYb430JRABghkBB185Tfn8mEB8KUutTIMsXoinZofYgjq6Fewl
jjK/bmT8+bFokUO7VwbXZMCbKw0+e7VpOdeAUlBkNS0leY8M+7VfMcEmoKOUBdlcuObm6CjrFAyI
EokRNEBvVoYpblFtPQPsp0ZhyKWmNisWite7jWHDVODCy47faRdfqnuRnXoFV72L9aM1yj032cFW
HEJ5+S86mBiG9iemll9fryO/P9ujMxOkhQOcbj8DfAhh/vxu0+5OBhrUQgRTkrmzxRMBKdrUogMZ
QwutiUCC34oV1SRwi0arbQjj1ZD4euPkDDc2D9gJ1Fsjoz3DXl9fvyrqfCSHQGQRy4cLZsfLGQdb
IACntc3NHMTMmaoeRyWa8aHBvv0T2J+BQShT0mlIjhxPOc9u4ybQEz23JbdmOJCWXLpFW/FG4AST
prPoeRE9GhQbJ2/v1kJfslLyW45ljFEdLzMaHDF8Iqmj9AlZRi6XeC4NN4VfmyXyHzVK2LupNXba
xtumN8XaSVsSG3i/AXJ8VgZtLXOcH+QGUTjiZB7XNR0RP+w6StCA2oC5dup9H94fCcwhXIPPk9l8
6CaHUcMUh7jbj6LvmB5/9gvaAmNdUmIX+VyyoseK7SOw/7Eis2HsXFWutJvMlGEnFR1bmOfkqHsR
DqhwaNtexOb3XPeRYFjC4i1dc0F2fwOTDa9wbMe6xeFZJjPU3zfBuxrq8wYFKH1MMMYuBhf7NGwf
beI1+HRqzV4OCWK2Wdzd2I+uhbPMYzmQ8Ao0FQNImWRxk7N42sHcTdNTzoE3f3arMlc/IB9qfsMq
kSEH1rBPNCPYIKJFFeucLMya/Es35tHaDofKMcNzF04RkTWnAJrRsxwXCMGK9pxnJkHTTfrEdvau
n4LmI0IfORXuLo3MujrzJtAfjfRTtwMehY6riGNfkBUh+FurnPTUf9KyuWyxtoPcbR3ejVivkxH8
NRl3j22D85Vijp05e0qzGEydpK+fzJekuJcEqPSDxXESvg9lp5U4eMuBtVO+xa1/GMtvfM6aKttX
CTi+xky8HhDu54zAd9pRh/xCU7hK9kZbUsvDB8bFsVEtWRtnXtud6y+N9Oe/ZoUtmWTKW/1A+1hh
BrtNxyB+Dy1eHEjEZWOHLZjIexXx+zLFzjneAXsNutW0kSJK3TMAAYExFgpl2DitaNvU0Wo3salS
c1jHw8FGNeO/t6q+DgpH6rfauoTcIBfYlFqRO+stHRouGZdb90yWccTlGV/QVSvpj/FQb9e1sQJv
mK/qlYTRoNsRh5w/uohXOsisEzuxgvsdPu0v3+pOcJVsnysiPtq3/hByAnPdBoKy1QCnC5R96wK+
EnQHCtlez57YTBW9u0/nAR+kPiXcQaTI+OJTrDaohgwa7w0Eo66xwkpo3Yosyd/8+z3tixw5OtMA
5VFsM5Q9SGrNzVCeJRr3kPmXnDo5mbCS54x0EKOLC5B/IuYO2sulmxouKpHEBLbTLyx+0rGucJ/a
5VnOJxsBfAUfZ9wZmqQ9dREjU6QhhAqeyv165YmlYbIB+COt8tGOHu1XJD7ZnUI1DBvLVhnRULzt
2AoaRa2rVSTnpObpPll9qhCOwSqg063q2lJsGH95KV+3wf3dWsCuwS89E++mQWzQrTgBXLVJDoLS
WXaaok4wJcaPEkGPMkAYeGqrohzli+OOBEfkbhWgrU6p9HUVemNIPCmQU4goyFW1byEYnJGEXg+Q
zXMkfLwaSm1q03grWyJzDTbu7ZaJR9TaXVr/XczKQJHjU3mL4fccC90a0GxBq05uy985X5prtS8/
zPYD1izc1hOuoyz9aUpKasY1I1il3zmKaPmyemqicu3VBn5P4eMZbkHRWXHVmcb0xz/8Tub/DJDF
ppzDQqFNLu3DzBaDwCi7qQTZgpf+xVrQShKSY2Ate0Y9JZT53LkHw6rqWuLet+nYeGu/yz4lPYZU
axkughbiO2wUN3bNUQ8etYw2YQZkVKlymgxgflZLkZjnPJsk2bKrVoRXOCRyZHum2h6NLAIBNIfb
lBxKE80CzrxkGtjSUU2sQ4WlhAFGRc4bEt6DJu52F8mU9JBhlnpC4BiL3mBZdYv0e0lfJP3K3iUx
vza8O2OQkRjCZdEdtcqJuDOPqIHbaHKFuiaRltS9MSbZQFeJEluZTf/fhbwV8yYc0rJrel3ifGYx
ElYaHciHpcTJe67gCiUuI0MV0vR5WCvWn22WULt/MyjeF4kIEsJ0/MWWkkxxUaVOR+yv+c9RT5sS
U8XK7p2ntis8IiR7wB2EvFZlipV8+f0mQHCdsPU6t+B0RDm+z2o/oATrVzTXxsR23y2FoQZzox/j
97SZ543+RE5kE1kg0BoAuIo1Rx0GgjlPV8dGAoQRp9OYSC/FnJtupkp8nHw3qFXSl4gTQDe8g1oX
CEYyDDIcXY4AmOMrq0afne9eFYojxtxmpbktjuoT71uFELRBWV5JbCtPqD0a9sgbIrlq8ib3sIDK
2mH5e8UmSrAskDJylBBXuNnAok01tW93oMtxc246GKiKkYAioGZtRGmAVTejYctDtHjZ6OBb92OJ
W2OPAnURd3wScmL5y4nFcw4yl2xLqSik++32ib6xaqsY4WmvMCFLnoXhU7o6wWxmxP2s+hoXGb17
N5aqvxZCaEZpHPYYgOgLyBRBlS2yQxUsVs9LcRSA6n8W3slDea9iikLCMBHAW+XymDfUGoRXsmAn
u5yctsBckpt1++wtr47y8M1OOTUMxjmM3PWaxZwWmqjsX84rAs7BPfmyKrXMdgNHlZatmJ+oFIgI
OqlKENHu4YbZi4xobc3E5t6LSqtNcl7PrAYGY/CAbA0ODfmI9rfws16Wjf6K5A9R/G7GfUCThUk8
EozexPsKY52UjsMOhi38uS+I7TVjez2W+i/kfRCXaQTkqCTKxaU3LIc1OMMBfWx5Co96RhJ1kQ2G
GNlAcgo2vWISggEW9ttbpgwVZoayD7EBeWw8ydJ3hRChLq7ulO/vHTIJuEcfB5MM/Oh2djEcFP9Y
aE55hG0THWO740yziIxxq4095gmDG5yeqW+GY4ZG8V0pZQzFPAK37GKDAixjFCKG3WUlB4INzCMx
VpiQhrnHHmRRPDMz/B2P3/nHim9nE8VUhyk/cE7Jb4knjV8zykfpSZY85Fo6dHCiMQetAJj5ExTO
6t5vUkrKH7+2GUgat9OtUWk2CnaUb/DRsFu6tVW8dGcSxCT5MXBpWX3u3tFT6jjPLegFcWB26tlO
hNL7N68qUaain1eylHJQVjeu7kLxGZ6BwjZ9LCKq5kXauMkXKwjRn07I66XVepxHbbGjnHcWeBvY
zrOWIFlIK0hvW817xYL79I97kzUfgGfuBocrRpl4LAY0jgqR8Ys4wOkUXuDOEIX+gtJQm+xOQFyo
gjjUsfQMbwGzF9jhHBJNFMElD1yADCtAgcMBEyKiJ6ETt4TMBK7drcYiTFVh3OrR4WbifIrOD6cY
qlYUSbOLN7occYYdrBDt19UOrFKtCs0ebVusy9F1LHlhQMyHENpjlwGksltbVhDp677uTJR2JoBD
+vtMYu57tZKBmpjuXclxiBUAKOHXwuPvjK0YHziUL0JqQE0Ey3mvXT75Dg7xrvO+xKNfw+QFN0rQ
K5X5W2X2Gv2j/KoSsWuowCXhRSTAcgwMCShSOh4iaIDOkf4t/luM1vO8BIEh8/cteKE/PLwVsHme
X/iyXIlC/JLNpZkNm42UUj7wHM9F/wQxbmuxivMRNJa4TfXch2Ev+lwCeqBBMkYxjNBtWHOa0wVQ
K37QmQC6+mpUtfI0gtk0i4RusXgtdjJmkDheSNbRtto+f99VBcBPmKRqbJhDlMwAVIYuUjU6m1BM
WziBBp/9EqJCZ6mNslo6dTaiEr7VILh+7BeMgfuTjLAz89xAUI8GfwIIscnPA/A36Whes9eLbg55
LzBEtYw1aySVofwDgcC8bb+bpjXUXunLvPzAlwvs0f8mRhMXG5voyB2MUCKfT7Tcy+TwlgNRNmvk
KdJ3vWpCT7LD5VushNvOAApv51tBxEuM2nxRFySGBwcZGOgQgdUCkgrsNwT8d2pbL1bQDXKYilKI
lBY9vVYj2GImInBEX94/hX1ui3ePlEaVglHbNCAdswvibtj15Hl+EkR4x6DiTDfeFB1PilrtHOg9
E+LB5Ne0uDTj5UWyQ/70re2tIqBaVocToO0ufySC8OmbEXduPBfzsBwChhfO3p0uiyD0vox9Px3s
t4vwq1ejaYyitN6ucDo7jwoZcgmCtfs64h0SQyncZxVCcA/2lspwGeVGtpolz2UcSmKTFYOz9lv+
hgg9f8wLuUmCIwND4SWfX3Wre5UXkkEklXAHUoHwOJBaqYnxLMKXUjiEv7in6g2l668IGfQRyVNv
AGhrMKR3/uImUSTVMiiV+/PmplIe8htzd84FKrfo8ZtFOPDYNagmV6EJulnI5l87CJpbAb0nDbYq
9zzf1oPPmkaZtESmt06OH4+VaxBBqM6ugAHMBnjNOpK/M3BFGIW0PFc6l9/Y4adhHfs/Yr20W8xM
LP9UWjsyNXcVyJ/oEyX4MuI/7m7PhI841g4SITVn2A7FqVwP+hSjiWi+CupI69HG5pdVp4+r4xxC
pwmr0T0EB1+9gf1rp2+eiodUuT2Af3Xj07DsFZUsR5ICuCp8cD7ia+jDFcOqi2WWCh8BTukzTxnr
xEJmrt6SI0yVM5Cheg6bNSf7luXtwss3ClJLTRU7JHAS7OGqRtWvbsxeehi3VDNEHOz9RX1FOIuD
6DFWzBvPJfdACG8BY0gWVl61iGi0ajceKM2dDPTTsXe0AROgpSU9NRNydfrj2d1CeuwSJdM+jXBV
KGdXWSYVXCkf0lPKPyJGffWLf1m2cR4NCM7RpjL1IeocfUAbATLYD79S4B9dmEF2Hmfwvy0sRNu+
IbNtuKOIhYLBzxuNHhSNj31BvxiLOcI9FyN1OtUx4Qn0tL4Dq3SfAZq9klDdxmbzP7/HNHGSJaA4
fbZPxA3sRvc6fTonJ4O81fKCsJtgM76uDguaFcsqlou6YLv7xuqml6Ii8JfNVBUWdNQyWg+vov/4
0owyZUFH+jn24sqNXq8LctQAMSAS6/fnKjWOk0eElq8rgB3/Okv2v3WnqUPzNZaq3/qy2fnJbZJv
qCVkGCuZLxq3qZRuz7d90tsNBMxP+cCk1rynEesUw8WhPWvIUVpzz6fJnSfKIh5/tVIY+0k4+5CL
rHgroiUILeLFo4dZtu1BB4vYniKhbnlXaTNqgztFXv4DEQ2gC8/PZkWacOcsk7r93FK+mJjJb4zd
ZznZ/TSIdsHmq0GtWIeTfxrRdOFwaJAb2y6rrQ6+3LKRMOeIRBQNlVEpOSMCuTgGl3claHLIQK4k
r3Gh63VzXcwU3gX9QF9ey+TClfnP5X0JBcjS9Hl2kkq2uIKuc6TAb/93Z3o4UDUyYv5cBTEGLyjN
sMpe6QK5/1ROAGwoHhqctgTYKZc7tfQ4fvonN4rsif9P75YzpRigSDjooI892DFIMTOwgxo9NSr4
kja/szuWAIOXx0QhZx1v42Gmw8ghjSFpzvrWriqB4bXJ3i+fsOGBnbefxVKdMu7qhwddJcGse3RX
pZgq6KIItc/HqjPfjm/nU3dhDuZhjH48BsPCIViMWIDI2yQsETLVsFD3ow8ADNaElzxWxK+mYFmd
4kWuWbt2zzmkrydbzOQPAJxXsIgS0oLcL43DhjSbKTzOFLaRWctoEI0e3xTqDjHGVbUDBEbwJoep
jMOMIAGXrvFJPlzC9c2oqSO0R7AozggMqY7cf8ep1BKpSrDv1P7iS5W0BeO4RTn/6yM5kVVj45zp
rxriNR085gFHWZP6MrrcXPVzWhTPsLQXovsVKNrcn1v5T74bxlP8aIAlDu6kWanZ0JE/9xHymFOH
relJeuEUHZothc3FUApeo5Npd/f6EFbrH6ZEGKSAf7qJqRndPasF1D30xAo95bv0odt3hzL6eUKI
U0q8iy+p0RafaXhYOTB0MH0D1cqJSKjBvDhQ/g8YfTx1jB+Zb5MEPlukJGnE2JPBKJWjcKkNZXgn
ocZkFvkc/yD6S8rmf2HCJQpWxQqrgI+G0iU+xwC5dxNDcA1gqWXrc7wXxAn/awszC88ExfniETh4
RrQggnerLfiurK2nRIQctVTLSgzesCDv5h4IbCi8s0uxSYWh+bespbyFhLOaL+/fHdn2s6c2x5hH
ptD3izKLW6R9uRGNtKIHln4Q4b1nc0lCPeOaRiSbE1hVTqKJuHH9wxaVII84GYpEXCx2wIt831TZ
rJVYeh5uNJL53xnCPZYtIqKYzmK9op8mwIWbF+rHQQpcI5+1dZrQcnRCTaa2JYICIW7CzHZ3OCZb
LrX4Wtth+VhDb3C1vm3XvtP4QFNrWDOkP/PP1V567e7R2BYquSyGhxu0TBTKUASvDES8DxjgLgkk
04aNfI7NwNTP06EKpnH1C48Ghw5TD1q1RZyC/w+qhwu0ii/Dch7w14ZaQ0Nc2pssDoI21wbn1yaB
UwzBV7kVLYgivhBO7PF/zejpk4lXaDlaayLUo2zIgunDQi9F2rO2+84M/nd3rg8CoXci2bLXqBte
zX0lt0w2ZRQIVLuoww4VDlLYnWT8a2FaCdYwt10VBg0FUbHzZaOprWqz4zRGOwE7cUheNTUs6IxD
xsXmtyVTEFp/jwg32Zn5/tzdiMx5YEIIUR2vFzpOvEvv8v/YeakLAi5e8jrqydft4vLRVne++BUa
QFpZ7gjfU82TI13tZwWvReRZH+Hvqdr8LiFgPDnhrYJRD83gGOwvSvghrvQrhPYN1Jq7y3joUciM
yHBrv2D+G8pB7NZCtNB/BIYAUYyTaD5Oxx0E/s3E6fwK9woFswYYbAzLfn8jOA8zXF8Cb4qvYCiv
4pZnrOlsdLzWEIRS/JSh3tK3HR1iVHxou6qH+oe7EO9IBCCG30MI/sOwgJxh+d3JmzZaKg8TIkcr
bqr1cAR+hEA2iDsVp5Htovp9RaTdIQBU2ztAt2m6RI3HePSM9jh1j9P8MU5QVQT7lvS90ZLYPTiL
iBQWQPVWPdE4WjgwHoijlEgZBBUR70dqGQE42IUdj5RgkK0IsppTnzWFvPsfrF+YTmPaM+A4cl9U
Ur+zsq4ar4dxSApTszwMGlZeLNprsD70kYEmuev3dGD1FNTSAyYkB3AVZanILqYvd0QaY8vwZT+8
PEVcq15FmQcmcAu94pDvjSHIqpb3BqXpKJscJXX8MKtRzh+jTlJSomJG1VpiscqPmSM8g46o6VEJ
hfSaKhehpeRjraEd0sqKqDsD0LviR9LVkZ2mecwgOtjVDNBkIjIwH0WMi1ksHWIdXZGm7jAjVeBd
f1GFw5e2vaY2eJ/KnvR0lGE3LxvOA5DcgrI05alNdau26ofm/NpNu+WlgVwUsGw4OXH4ZfBbIkwq
niWKMc08OPAxEx9H3levZeQK23r01TJGlh+gFa2u2K5Uj7ide+rK/8H23W3k+l7l0OwL8qinVRwG
g/awopnqs6VhP23zQ/MQ8DT3jMki2NjHSqcQJuE0MIRsZhJ2p6Qxkh/FTm2o5vqKtliB
`protect end_protected
