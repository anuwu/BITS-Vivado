`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ay83AUpql8IXjVPYcDPto0irEAk3jafaCXcP6KIQNpP1g2NRPF/2/jSTFn+D2wOi6J7f1rZs9vsP
46j7ooq8OQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cBdSm2HcUM1IChVOKHkRJNUocglDuDJSFxYlgtLiOwZHhsfPwquUtQDg5m3+7UHB9KsDE+lsX2K8
xD653VvfGyVusStMqlvTiGailRNCMoET8Vqb5+EMWZDjsah3R8OqMlduI/uK0oXVO3ZdHR8tVO+y
OFmuMg6h/oWeWTVs9sk=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
boswFhIjuW3JrpRcNOhZfpm1XDgdd8OMyWaFbWmG0yR8eGpODhEXr1Up/HEpR+Bt7BnQQ3YSB4/0
bBa/PznXzObsSKwrxzJGHewuQhbnfvw8DcjNlM0XnW9wZcC56ui9+Azt1X/PHtz5xcaiIg26uMNh
5quyt5G7wBvPX7i7dtXVY3UjcKKa8rItkWdJl/s3rsL6xv7SBTERGEn2IB7QVvVRZizhdin6Intq
gUKQebQCJ/V7ytfrfVs4uE3UrQOZD6aWVcrky8PNaMFBNsFGQZ8P4ibR7frajP7ANPv5egT0gp/w
sRxPMaKn1SM6Pc3/XA+syCPQ5aNshwmjO4aqvA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aV121xtU0Gz/9vBJBesdl2ebJ5C7vVKA5VC9dkXufCT2XRyecXYuPD11eqDp5b22Euqvht9bLb7a
Y3c8IE8mTGhBgpgMo5V1X1kPXMRomXG2HXYRo8NRsKeIIGLBgAGNYtYSGFXCj47SEpYLFZmgGVIv
rqMOFeXoB2g153yJ//3Btb5hejVkMgvrCeeFbzG77iHTfsD1MX2moqxm5YquVRyk44ctqFvAiHou
cqOLt95c5h9FL68hEJZ1926og/mYX0s2sdasy+TjEcNuAg1zSggJFmPBkwz59BNFa9eSyRZGOPYi
M1rCGju6Ii6/IiIrSIDYxDOhR7SBx5h+n9UG8w==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GMdD9bcV09glvUrA6wL4i3UtwZYmjlGSqXrRhqV4p1va8zfjBeL6jDLuyL9V1PgeFs4wrzLN4jTM
H6DVgJ0diW92fz6VhvWraRVpHUg854lOi3hCBBSTI72zX9AJgs2Ty2H4VBLenIdhZ2cLnZPAwDjg
AZqCBiQ2rIagPrVigvTTqErxy25jemkSvsasjgmhlPwCYXeGvaAkIuiCaulTjPotxEnk7XK72DzQ
i5LG3ijsiUWhm7840nHR5iG3LP0HCcgw1Ou1E7fvHPmjGBBJs6+53yh7VdYZAn6i7zBlLW+tG97o
DRtO/sNA+hXfp4YK4axcF7XPkoFQ19LdmwR5BA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bEjTFKHXA0gQCUWeKSbS2CaEpDRPTIiHg1FKlh80/QPF/hSlP6x9xe0Pq/myQetv5XqsgeQEJ92/
UjMdse8Hg+I10nCskIP1eqLY4U6Hr3EFT2wUBknnJUMdrctNkDCHmBgpssH9AXWQPYHf2/W3bWmc
20W61ePZCdPdlmDP78A=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZH8MXw2hh/beP6qBcaURW/8Os5PV4Fl+6TNk/SgLTWs4GNrNVURrkcdmtKF8E51TvbX/Q/iyNw3M
GzkyOHLfeCJJ3KGt2/wXkIfYiyE6mqp4S0LI+Tyaf5rFcBcgJfBKn74DUmxdZGX6FX6ACt65sTSJ
Oki9/ElsOGRaeHRTuscVjGw61sX/ZDNfRAjeF5ZhSpR2ORHLLy/y4XF44x95o4SK5vVOtNjiJVzi
DC9skLIwL4rQMuTV+cN/587xdqvmMVsVQZzguMbRAsd7+Dqf00L6jP7l/aqrXPL7qVLFZGha93BA
aQc5hLquIf797wDYhhZ9tF8nL1P0oqlBp5mhbw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fkZOJxfDoliI1UzcEwBQDgn1GAAuHqa7R92GpHJzI+jrkcu9kTKarddPR3BPozG+6peBUbORZKSa
kNu65cB8ufh4VXBVx77J06xSSrzIlWsMZgomw2IOSky5BSir5F/bQa2RxunHreXVxEz51PwsXSLM
SulDW/xonyCF8+09ZQEC/CCCZ2d8dRm4Un5tEcy58MH8dUTB4fdonhn9C7yTLnCKYtdF7l9GH/9k
hn2BTJ4BHYlDjn+7d/+vSh9k319vgeEVFNBG5oMnLhCLeAaCW76TqjKNGzKS3pCgpsZa6lO/emmY
aPOA/yaow9Su4vVxs+ZqRFVKK2sj+jadfAajdQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60576)
`protect data_block
bjpsDRwyZzqTLbg8dTGn9iR6QzurylEWIullL+gZB0JWZtwokxYL/SKEXHqCfkksVeG69MGOTM6K
5uQhR3DuKXLeR/VPEKwollwZEVJlQseohBBSHJdw959LJdCmsubaQjGMTJNvTwVsiyM19npH8E5J
ruCfi/IcHVjdWSTywsZTJBqSHcunv4nemlEcB+a3Jh6uvqzMroCM+6UBrGDeucRUJP0Qm6YiWhi4
5PHOfB4jtPJ1UFBo2gTgvM/SfQJJvwJCFQJxyMjfkSwHpIkMZ3KgB0Wz7JfFa+YEuMZsFcd8hk1O
12fMoLRSLJ1fRCQNkpAUz4UKQC+ioIHMXj/y9q9JiFmXitb6qHrbgNr40AYzzbqROUBRyKZBRrQZ
q+gVObPDVAHKy8iDovrmLdOt1/b5IXr0aVMrQpoa101ISyhTgIU1O8VKfrmMb43cEW9zNQw/5klD
q2zQ601SjnqUJesDTlsNcOaj/VGv0M3yZhvGgdCTgr1EenwVqik8jgLh4GMiXBef8zg/ZhTLFvoj
SytufKu+zU/tZLQ+avg5Dz51F7XeiZL137lP4XdeTuAgXqEbT0bO0oPthHnGhT8UzPAvbhqQveQN
DCRiWfRnoZGJBBSSYtXwvHrR4kr/cCGvj+qosYMe08MJAafR2s0dTtrh1Pi2kY3Bit8HuTCikzFH
ITsiLG7x5buhZapDRG7bup/jU++V28LfkWl7u6QM4dEWM4cdtXlgErOPlsiKPoxNpmB3tT3qxi3b
6wXlPtwbfbhHiVwxH8FI/z+mbFB1au0VEFoJIBMmF+apRfRRIjyJs+eeRhE0ZoRhihTQ0qvFRUFh
J+i26iIPa0eERHPIKrBpvlFd94HUfxwG1xpMLcs1t5a8NqvMUPjC7bBt5FlIF+mrwG+q5rc0ulLQ
h3v0wbLRcULU/nhyyjo9AM8pZQs4baCBfuwo3i/3dyHxw6gZFgFfyi6w2DXlNb+Mo1Ukuhf53pB6
5CxLBZX/hiNS0KsFTlIQeFB3J4GJR+Wn7BF6NwQefRYhfegP15KMunu55MeemBdEc4CbKvTWnvls
lsYOPkn0CBWvzit1YRsRww8lEQp4a5F8Ioc8pGJFtHGAAOTvm0ytoEFgbJ5BfihuZUG72bmWy4+H
vnfMzdhCedEQB05MxH4y9v7KV70U9sCvR6llbperuGwjta+5PlRmB1/LuE8dhzIvrVrBn3vAOvdB
0onQSe1ikD60pTIQ7Ylb3nR38OZhoCG24heZsWoXkuUS5VXveAS5RzyHZ7evKOzRSCe9rWiqKcGA
2FEd86P1KWw+Fce9otZ/M7oZAq1MqTvwyBBS0HC7qpdPLJrsEkJv9Alg9gaouGrOvJYGIqSFmoVw
wom7bLbwDJ4TZT1dfRrJx3LYpc1UAyYiCk92ED1JClDv/dthA6Qus0XhnWr0fLS9mpZz2aKoefwQ
RmdLlXRUNYqrFemHFOz8TVGY08vTrdzn+g9095iJyYaGIkcX6nGnMfhxKf7NaD3Gq68HRTquXnUB
6ddnQjz6e5OUSflgZhouE7wzk2HtZE6HYeET9kJVxadSN4n7wLDAor2xPNE8m7kxAG/FbEzR7h55
qR4Vxu61Yl5mYveLGFYlt6TKLBitxD78Mlp2tdFgWBGkcJLVizz5rqqGdrsY/CJ8nra6ALxPH2Tm
cO8xKZ3WBxdO3MEJfI73ZQ3u4qgT8VU1B2W82R6X8lx+1gLZNrBO8o2ED5XNbE65kkc+Q/dEF6Jg
39vyf9gwLz4XZiiGtwP2wFuiBS0Cb52e9ZxDO1haDKyNJ77DUepear2oqzGJVwoGIk/bmb3uQ5+u
pp9xuTbZbAjg0kY9szDYC2PeCJ2EoweQn9GzhXw+GEPgWWsOYzKrxMrahZahxZDBgw9tml+uMRuB
6HuE19tc0U4ZvrY3qBfhd942zJCstuUfRnfkNW4HOzzOXBE9i0ilXm7miCBDJAytqg5ftvrzqcKo
8gvE/1Scrb53X1Q3mhz4dyIz1iU7AFhVkYftgW3nKfhfo8MmNFBIeW+dQ/wMME4QjCcEO/geh5dM
kB6WjprQn2VJ4w6fv9K7fDB1l6MGtFgdrndAG86EkUlPZ69/PprMFLXeUT7f7JlzICRpbLGTR26L
kOYlq8vADSp2ORSyuQdBqHXy4iFk5BhajE/B6CUr7Y6jmQRqthVpjPlsMNJholKuS5X4ysj5TzOv
+jJXnGc7v3zl3guarmuRX1Sqtu0L/yyx6K/yNP8jIUT67J7p4mlWHFcPlIHYImLS4J4YAU8Z6VGF
8Ut5as0QgGfvN67xNoT5KhuFJWqjqv2s2SEZgDSrPgq0s8BIymYv+niJUMx89UW4izyhlc4wPOBc
Q7W0ew7XDIbSSBFQr18SEE1+0Br5r5r0pnHJ72qH2fPC2TmFyiIrE2/Qju0q61iN/YsILbbiIwfC
3H5xhBd84DF/htHh7qNph5X3qgJ3fzJfQYls/P8HDfrMp09pYy87ahZxJONiVWBdCTlqwrV/zxcH
rdrZaYdIHTl7ihrjoIMCJXs+/7CzQgzUZ7wdcsk/s4Wx8l0GGfDveh1o0k73idp8BhsfWZqyB133
jdcfTBwPG5mnRAyCW34RiMQ993QdUrtzzcN6PNwVB/1xs7hKQ0xI9GWLVZCcCKnUvM0vrTBg3bXh
UjzuAZ8GvSTbyGpUMfgnKGoJl1yEnoxQ2bY/UCCdeYVnzB14bJtojsDJkDxLBONqYHELSXhujoAa
aOBpZ7ug0epY0EgmTH6BB8Zm2FY3hbzCTSx6+1nJ+MqH+O+Sb3UX5k5RrL43U/DXVsl3CxxcKVpP
JMcEW81t/EkMN4RmornnT1JLmnydA0UUrwl+toViBvy44XK41AsEL2ZE2CMyv/nurpRSLj1hHJpl
pVEjfke0EdWF8klmCbnBeSaMupwRTTK5wb/ldlojDVTFdS6BB4RAxyW9x/BizgqNA+qtTbudxDpl
PvrSmpPPI4ii3SeDGJbZLLTi2Q60QFvb+SL5b6lONPFcu+JtJPdZvYHxXX0d/jZdiaJS5rX5Ke7A
IUtB0HVWYI33MJbC/eVSktYKtPobuT9t5uucDjM/qcDQfos6qpHbSSPHF0r4OkYVbLnOwljM4UxC
aqaCIPzvhztq3LS4lFZNumg5suC00kw2Mu1S+l8z5bjQwUkAITBZBQUAB6uQSryImTrrL+4Xbp8r
7MWU/ikmi0NPT+a8Mb17u8RdDMmUEigPv4JdMnkOkb/Xy/HbejOjc/1DP9QfpiCcL9QRjbqhAAI3
zO48je9sKQ4IjkBR7AP1I67dvGUsPlREhquzae78HXzCen1sYI6vRDeP3CSksK59EQ/49erjZF6r
gKzmkIAeL+AUjJCJO1jsWReADhi6Te6LXj3VbU1CtDpNVlmWDUGfu7LI1U/1ovt7LSox8D0xMLXY
81JVHYa2zO6O7EwVElggbl64ucr8qTxbl4bk+5YMNziJ6RRFFyu/8Ry5dmJIH2RF1tMYAMiJ6YTV
/oxOH0KwN28RsIdVkzsDbxfcUSkgjDSD4IEnstTNQpwv7nNMJdzuqSvlfKwinOwOxlnEkx8zmQuN
d08dS2bfpvrqUqDtmyYkJNj2uZa7lAdA8u1ZLTDp+iNNYLHWJeA+GPGxiNGbQYVvhlZSThjNSg7a
e+D6KDoSO2+2WnrqrkJWZG9qoKQ3N9uzAumGM5+wi0RqAMPeZKa/RBF08GOatu06l+4J4Tg2tGsS
s4T5MQzRcr9/BLJYlsbwVLGJoItV6k0wMDiZ3dUiq75BvW+QbJ7XlhhMsRRdrO/2sMhZcMtZgVbn
It1g+MJLiWL9RycEEvLWUcu+GzduSaAhXdCKX1+/oOEEQrO7oIM6VRJCJ6JyOSSp0HUcsctIBSL9
HWXR4XF5dItaQnKUsZj+vCW/xwuWN/PRRt91kUwZw5FEQ2vNuj3zU1p3h+tDFCs2o/lYOf1X7VtF
GSk/v+JV0TclFT7cWji+Pe+iXaIvvj3KPiRKRfZ7kllTGdcFkklLIASf0RrFpobvsWQ+nPGGlUeG
RqoxcX/l4vGq1/+mW0/bbcq3cDl9Ld/Qh7XV0hILTXgLp0Rb4iK+XU0LHrgUYWinGXYr7GMV1tUb
3eezirRGMa88eiGOlEnoWeBfa+9qVS4aPg0UCYPFbmtHV+1++0pZ0KGYn063VOdykj4O0rBqQ/Sw
sy0pDLlptDhHWReQHkCapcS1fF3B/gJmV42UKdIti5jbnpiz8zfrf6Tfthif+uTgDcVjb2GI40ag
5IQt/O4qogSXEsFTCV2dQDczl0D0w5KhPAv7e5SiSpm6jV47W2Xc6UJ8zoRcRgC0djh+754ufU8R
EWkOy/iWEgeWiDqeQkGwEYRs0M9VHIYl3v2FEIthr3PLt+EdMgR2HZlIF5OcI/92hCPDdhZ5b5dv
uxT0dGIpRO8uGeCwTg7lo/r5+aTlsX7NuQPYl1tNyuApM30e+ZD7qrfjYDSfT42NOlcXRuD/owdc
hEjyTR6VlBWJtrkX8rCQaQ0sq87AlTXqJdXSIVYZy3ZRjz8PHYeJ0oxgxMpgvRhHTfQQ+4B0dafL
7oaulu/vDMSJPpZVrk3KwJ7D/fBjwwgU41svKbYfQdLvNqXuwDE8dLDGL5O4K6jj/uWKnTpFr3pU
l86pwA2Uz3Kizh7W0++d9aPiR69Ki2h0ce3Lc9m4Ll1izLGqzSEXawcgrw68j10MFZFDhZc0Tqu0
kYZsRS1XWNC+GtcG3ChexpaWMYV2yGXZcpW1mGhWqVByJuPcbOPmogT+1XsQWS67KBUc9sg3apCY
ZEENSKk3J8MiUEQP3T7H3rg/k47z/R+fWECgKiM3zuQ409KC5xii214jxXMRIPdE5+oIjZbaLYRg
CGnybXYrkjOtrmkgBc7a7bGsSDfUvDtbwqg08j7Tn7V74jAEh9fPn0x9eRRek3/L95ezcD0k3SOk
/BI2xk+lL1iOTgjrUO3LeRLqXKjxBcyA7iMFejkl13ccUnOyXtNn5FLhcvR//UOUhRn3weTHkL8R
LPgKxSsqt4nl3+PeasxICvP7LTpzSqkxTuy36JyxwXOVukTHqgaartX4M9HErsZ8/rtP1KP15/Uc
GUb5NLVWh8PGkw0OWkyvZKiYP/HQ7TublsjNfUS+f/sPdN3FklcANRZ7AhlHFkr60IMMXnETMIDf
BmT3lPOED1Flz0q7fu6I39MpPEvNowZKw6P/BSOw12zYoltQBQ4bG+Myw0CqAT3jB3s+s8u/QaAu
oMx/8FB/dovanTneQUlDWnf7AwYMW+LZqShvx7Cq7x3Cz79UybdBd/etffNf9uYeLEGqZswmybtX
9r5kyHWFpSiw+R41Al+xjSUi1TgHrNehZPyxdgD2cVigdp675/ERPmCD34A0as7wktFUJf7fJe0X
2ZLaUhlsAjBrd3iAuHip5m/WAWFbRYnVN5ZdGknkO3IoJVpxTYW9ctZ6YFBvn7nBLMZHeRRAdlYy
5HyN24JkBCTDTFAAkoYNJw0TUfvAZ6k9pRU4TpHuIYcnNCHKB3ZsdgAB8KlHW0s+HX3fAK8IE6cS
g86VLZS1xnAUuj09xq9JpzuThZbinfU0J/hnkx9eyPrACMzhhkkOWfC58nJo8UNjy/dxOjgdt55x
u5ZPuaNCKcVA6lbTvGZboKibTRvdiWGp/LAqQY1TKKr/iegvHlAMZhjMiz5tUcd27QdnvTDFaCD0
aJ2/jyK2zXuwBVZ+UtFptyOkY7dk//gchOLy9WCIUjP4x6gxR/hI1oLM8i5lnajUrxpPNZjbRlo2
KZ5+DghjXi3X+25EtB5gdntQ56joHVRfHjWn9F/rRyXl424YsbyiBzDDzC7TueRNZPbKEsxCGuIz
XpMx0YW0y7SjzM6rz1W/IaunU2wBnudwyH/jwdSV9Xq/eOjwyvZ6b7D+NgIRnqWQdJ2jcbLWWBw5
hkphg7jFjc91xXDXm8G7WbCtcTPua5cUjX3dfjhaIfu2XuXBxExppYtlz+vscbw/CFKbE9Vpik0s
0Rpeu8VmNsohToI0wAdGXZ7IOSfDazuue9dSl0JAozRtFqC+bd3wHNOLoEL/xZutLU4wstIgt9fW
Q5nYr5cXI/IOZdwWS/9VidoNHxPHGaaP584X7X2dbuiWvpglp9ikWTUsksK/3q6Q05c2fPxzAJY3
XpkRdWZS5ktmhtIAP08YkmwgZxXDdt3YkrgWZ/buT7MFyOACMwqNSfx+FbmUAcTxoV9Hf729V4v+
RA0ToKN1h4/Ey3Fo9wor2fanSG1wHcw8uC/qZxrInGuuaZO1izlPeLOIq3lFKSRAyEgs8Elq6Ygq
AISTqIcQRonYKWfL+CEVKFShEHFkR4bkAAqgDbJmcNNVALuzP/Fs10jFSL0x1O/kpRvW9FkIiCgj
RV/MQ1FFcaFVQ8u6eIgdik+PHKxvMj8qPw2NT6+6TlxyrrBDF+vW6Xqu4ABDjpPVZLd9GStScsXj
9AM8OvOHMWI486bixMvyDwIrZJoLXywnYuALo37lcD4ZgrD/BbFQ+sjAGe4bajzULzgr6FUW9zQj
3u8c7Ca1y+/uvw42p/ZWk2SKOUQUA/OoMZrmCNEe57u9llcwE/4w+MI2eddKUO10EtU2xIYa3RJX
NvOcAmJIzeX4gaWGNRoXn6zPEbUgSm+RMyDK200QgtEwJk6gzPrTUvWkc0/qhPJTtyFGpY6efOG+
3MQGL9dGi0yljZZDvU8luslendMtzV9vQcyJ4GjAOVJW7ng7KP2G6RFGL/hd3xjarxnrTA7O46nQ
9B17ONQR49Fn4Sjeb4UDdO0xM1tIaANpdJJHyxjUPf/RtRaoqOKXkuRKFWGl86m1QX2LgsUp6/hV
ZF2AGv3u22Ywrj/PNMy7N7xEJglJnsxTDW3guzhi7wFJh/LiOwwhfVWzGy19Pjei7w+QTlHL3feE
527TXUa/j9h+v80Ih3fCgRtY0nWQbw+uOt9bksY6fj2CuxEfgQvRk6p4XZo5bRKjwJMz7f4oTZD3
9fRu91fhi/lE9Rtpjr0BMu9lGRRS/jmqQhEDm0BwSRyV4ez496wUZmEoIRyRY7vTEKm4yBRNGS8x
NtLy4SHb07tqc8Pq5JohLj+igTFrmebHcw4ldvTx1aTumqWqB952NkfEU7p2RacsjsSPwb3OyK4v
aWbrVjeXqB9f4UxY7vFqdbwRdgrBvlyG1b3/s/BUdsklWrYGHvunom3Hlv0CSdDEXM6UMB/z3dFi
rg6rVlo+raqicCpdB4qioMYW8NYlR8SzvIdAfVaksxHVLHwRZlX9d9hQvESp2QxG2bB+yDSQy+tp
O0cwl4CnvnQZlXkMjzxwv99MyCQwv4Ex5AxHuNjQMbRUoeMKPHbKroFdkMeeZ75NBqFXDqGzr5XB
Gy665+YRaeCJ/u7FdjsVAtq99kkrzl5pQTXW0QjYciy0lQKYG9nzT44wlHp61j2Y4zLdAa4vDzpB
MEc4MdlHNNKW8jCvhKcLg2QQgSaQUpMfSOi/1rA9FeGzFkRMPEBuiatrb0kDHwMwYqjKNfsDyJqj
s8LS60iHVaVWnVxXoo5OqadbTbMzkwq4S1qyK8DTW6F8IvFIvRdXz8bkqZCKtJLPuKO9g+zcKm+t
a41OKwlZVnXwHKcDH9JwQ+wxsFgNblU6pqUMvCDQGCIKMpOVCEOwP6+IcaJ2nhX8JJPdB/uHhEPP
GkrIa2n+6HIhkbLYhKbSOchIMOz149LE/VtDIc2N5D/3tBWVq4eCGzI/EIPf841wBBEA7ItjYOob
qpK06xO2bvLMehzG50jnatWTuGiSM91vCsP+PZqRTt6vTu5EyuzE7XQ1LfcV4Xptvh8siM1ZbY9C
SJFodtKM4xkqZ5j6fPNZYpyQpATvH2qMf3wJM8J1mR8nCHFv9VGHj9qpmRsf7enyT5GaJpeCWqMC
dKqp6dkC2jW0BGKPO1TMV9bpfWMmLUXDs1+wr1f3Ew6lHJjwOPMqUuLp/GKhCsEhXngs67B1Uour
bvavsnNDEw1UUzmchukdEr49y7KAa6X5Oo9j7oiOYSyvqDCJUNCR65SlVqefWkcXXbSTuyP0VyyB
GoWTiVfjhHctjvVcuG0wTApBdfmf35SF4k82V3p3qTziFU8GLqhKbtvjKAb2200mzLWrFYUq88Yy
P1dE7om63y0nU5AA/asw5CQrhDfGjdaG95I9/wCBQH1pI4zY/RWiojD89aMRMAGhxUzbRIUOQWVV
WPJdlFvmsH3zNoPAIOnzvF5MkEQQyWBRXPh4qOxtd6Og3tbMl83re7JdySKA7/iSYqScV3d0M0XQ
57FQxU38C4ekFOOAiDwiN9EMr/NievIrcG87/A2HiDOUrf0Uru5j79W/JJBN9qT2YY2puSNuXzj5
d9s6a76dAxOudTQC+ggVD3PnAjP1YrA+dtb0YHJvLm2JpiSdh05fQU6uglR2nxA2aEv664kmKzpl
dB/lD18w8H6dCpvPKxTxpqYqiMH/zoHycjyCSKqg7+eD7ilcj/r0N+IDirV0Oq1Q9IkGkvnrQPak
pt7dYg2asvu5JqgMgDVNLTCwKLCcO2zJlNN2PN+pNZm3LJybdTb5Kqv/sZkuzeUaUWEL/pgUtk4Q
tGaNcaQ4GElnwDqYh37GkLvInUZHElz8M0u7ajUlfC+/5AZuSd0Q+zcZY4XQq7ZU9qvUC3xhSjDU
c5zIgZIhCglzo2JgxGV1U30cnlNQjAS1N2H0L2b/GLo97p8D9BfuXZOKI5upoGggSKpT/Uxk+lj+
jh6EFia61bn6OKSKxLUkQYQ1JUXntTr+XuH1s2KGn+jt28WPkSxRkA86N68b+jqWXjVaXsmeFCCg
e2p/dLKs1/JnxcIHQdQSvxdOQTxCSi+m75YdabN9joIKKSywB6rpmpRIFjZFRLscxnDEQmRrvXAi
L4sNG5+pGBkovctJUqgfBZUMXUne96c4DTFlXVu1GU8p4S9QkkDvb/7JOAt0Xv0u93rFoqpWnePd
WnRzWjUf9IwaYzoa5dj55TBW6JjzJ6e96L27lNPqNYOXLLn0u4Jy45sTtMXjmJsvC8nSsP52rjpe
2EJ63exHbjDLV4whgeRnMgbydY7glnqgzenBiE/4Au2TXTe7Mu6xxoq++fwrYBkEp7s/xnv1J2Jx
0u1QMD3hnsLybRMLCMTlYxwmN5JBv3Byz64l1II/tDwQWkR8h1WPGQ2q3N0h5XHirqm59KI68Jpe
p7Iq5BxFzN7wU7QCAnaVUI7WI0KDDzcmnfSxsWUZBYeL36s11z6Bu+OEn1+gMW8lbUnhiyDbNYQ3
MKrraufzcS0+38KPX6WjhAfCgoDAHJNfKG584dOhYTd1eyjaoOAdkymOxiNqQygDGKt+llVzip9V
UnnXUZgQsqQYLrSq4MaNawnlJEMTZ+3uROttx8aG1kiX38/4Eth7GzHB6MZFWCFu38MkK+Lh6sgQ
AvaBjEExNUydfFmbEZdrtz6NXKntUkKL3CYPyBoAIhUNgO7tV9X1tuKZ5NKzj5t13ok0Qnf3dkLH
7LH9PXqu/EIdapRZbNq3CXlo6vIk2pldS5vzJukmgAS5sKiuphRdiRcCtr4s8ankAVNMYHsArsKv
zWA/4ZswJsXuujOn27GY9HHNcvQK3JIpPD8gbUZDiummySKVKYBNZZlITBvBnGuCSa4EvoUVkTWA
4BTLySlfuSmGYkKVaX11jgjaPiB7FnXuCDqjcpEFMIME7YcjQEspVRFcZa87tK3MIY8k+ja7pQyw
TStmRPt9jBp5Ma2ApDu5+9KGAOweXV+2L0YDYds/wiEjmHWEw6f8In66a5XVJIipfh6bCTTirAO+
5WyBxnXA7Gy0El/Ck0boOIMK1bP837GOHP1nfvFzCzZOJzEjjb+yumbcjOsEkibqtOTtgKNqJM1/
sifwFeo+2exFbKiDmTZL+0OSFDNp3xTkqMsPbNuwUJWPgVU7NqkPSis1YDmuYfsE7U0pByf1CRRz
57dGoWi6rr6bwQWEn07kUye+5knbgYsFbMq9iEu6igucO7JDq0UHvgxcO17JoQYGqg7Icg7RuI4Q
lkH/YP9vfzxNLGg61YJj7ajUqlol9DD7XJLbECR+9uGg1osseldU4wXjQAEAkEbmPP+NwG7fIaqO
EUShuLBE+6dLkeRd4jyIisE5s8vEwPYeXKuvitBkQ3YHwAY3vYz8iWXG9n47ED/ElaZMF3JHrYmW
fe69at3kjcrZIkqK1OZwFhegKetaNKsppMr/8zkqVIX2N+4XWlMEfjk5XTDE0dtjjBDP4u7Th6aB
FY+vU4xkBwO2Vgrba7Gi0lO2x6XLDQ4oQjCa6ig+iUZOwWIzUNdfv0Mh+P0JFgVqWGv8HRD/xWEq
B086HaJoZBvjEyWLgu5Wc4C6Tkk3wmSazhpxAynw5fqu2LKOvQ0dPAasofSV3KtY6dKk9g9LhKTL
lsqjXZjAb1GIepJo4sZEjwhqaXoxMhTYB2UbUojRNv2GzkUXaO88GZ8ZFVpai0q+Jrgul22/TP14
KSYRNi0K/eRsASR8kcNjoXLzP0kmg+er9KOGMlGNrpIC3Ir/LWsyO6HgOrmRvkfX6W0EJFgaMqji
iPG2cpvu2ZL/ggDembCPcDUPTMDMALXP6bRzF47f6S8EFBWvWoc21nwenFlD+1j8JYu8llzhUsLM
YR9kTWLovhfzjySYYSiu634f4Sm1vMYQgmWUkuifmEcE3Iqt4K8qJqF0E+OMxcNGHWo5J+HOVgMc
W/Khwew7mb+tgfrRWV4GfJo64/JbPyHTDhJdDhfA0kWZ+6oxqjdlboWtlQKkq9FE3MUwNaq4jWVz
loNHAmSZ/7pAyoIvX265Dt3kweg6E59BG34TYcf/YOmVd8fCvyfJksVFfPRo5Rnvf9bMYNbTwHwe
/aWKG8glL1BQt4b+nFaHMtkggq5iQefluHjDJQz2WZtK5KxtCfHJrimzdRVRN40ln7XDcaUg369r
eYijd4v0SuFDD5Niv2qK4oLPJQiIBYwEyHFwfZOoz1TUjORalVrNJrq6kPz/ZM91GT5Nz9bQm5oS
TXTH9st9cm02ROERknACv4CaC6M7d24eQEUDhjJgUVQQCo5OYiZJJzqg+yJqdvmRR6ytn5cI7X4P
tXduVXF4IyIXd8MDlBVPZjjPZpfrr1npv7sIlhff+j60RqthHzIu7PNOjR9HZSDcLTMtqD2M2thw
LkpD2woq898bRd9HfJahqNJuXyiHIfVBi/eCxfzY+DV5ecb8r1VJX0xnaH1S7RlOHBDx+/ctrUpn
DrOZoYtDw3CmdD+k9rAMOy1Ktft4muOtIy4CFM7x6RADQ/Ef7FGppGr+5ozRAcowICDCciDOSUhC
V1A5DvlU/rANq3c0Er4EheOeL8Lexfnzat7n32CtxrN3hyj2sXXZt8gEg8OpEJKzgWBuSwHzWhE3
tmwjoWByME0ZLBVj8cPiBjo577kjMfsg+UXP8QV70xaAU02cPIOppw13gpmp0J7P8B11R3idjNTp
RUBGfWfJtbMYg/7Nl7Vip8jy3Z0QevKJd1pswN7GTopTm2/dbyKFJP9aVFS5R5JtphyreJV2fQWY
ZCCB+0M/3s1ZjMNTZCIhnkOoahFFaeq9z+4uTubJhIsvyvDeZ5tELXwagYS/iuReoeLLgEvUqAZ1
cgfs7hAdIya6qPW4vuqMM4ob1UxhDIN7+th+pij30jiei0e4B1YVeDw79KXoP03DY2wj1h56Br/n
c9O+8AqlwqdNuE0O0kGi/iG5xpSGZl0zW+x4UbPAy7iPVealqkQ6RouOh5OfVYhoHecS9XSsdmWT
A+BGXc2uU6LAOvj6J1MjLjOaV0aEqW735S76A+acw9r4Qj9dg9WfwZ8Cs+7QglVoA4vpfiC3C14M
EVxTT+SFNbncSjwakAbZgOc6XJvU/OmD/GaBluXDOijiBrLUxsgGhfd42oIK6D9JkbZ4YOiZf1YB
TIokMkdr16TDJerFpDuNKdzZWIRD1aOZJByPuIJPBjSnzbskJNL9G7gkEZu7ohUrxyKmGd8cA9n/
9vnlbm0u4cpljSoiKPjRYukAdjtyEbusIIM9yaBRYkA5spZrPCF3HZ7fMO2YDMH9RRuiBrGHRXRn
T2bsyus1lElpMYOI9whW9ciB7TQlbo3PyVBcHDWq1FjXwyylnL8S3XTs8sBg2hxGfTfG6B2MWrT3
r7XqBIsFHKnqgSHPGec6RpAlZmuNKfrR9LjmbeE0aUaXUvY/vZzmsJOQIRCSnwXg926V8msI4aww
FWPo/lHE4xmzyLh3QxNIHnEMavCQnj5j669hPVJvHjVJxFy9dcx7f02KOV/oERx5NJasbotedXoa
JVYR/6sEv0qaek0ewRnTba5ViIRlzNISro8J0mKOJi8rYtNZMlu35q3p0eimtb3UtRLXKSA1/PD3
ocx5qNoxDTsX/1FsIxsRoZ3eVEWNi2l5ES+3CoG/O5rveqKw+PTrkSI8CcIarzfEb4q9HCnVYgLt
InTJdx1Oc+elH+wfcprwkyOrNtyakxJq/TaqdYIIBBPFYb6LVvscVIXQ1jYozYSZoqG+L46wxKpj
dyTC1DbF8CUTvqfjycEoRt9pLadCRDxPMF5fCZmysf4pM5mOAw+FWGA2c96SVVa7vg8ELdtPkrcH
XP0web89eN422UFZQ0g4qg/L+aw4IzHUz+iTIbZ2LZru/sngGeZeK8yiOGm4TWHHQXWxMOH1X8Hg
WO4CrI0S7XDchLczM4MtS1b/itWy7nwfoT+NzXCdbveBweSYJMsI669j0BjFotMpHHvFWsptXt5x
N6YDFYnWzJ9VWaUpGw48piwOhcoiEhcEWPIU2ilevgO/6yMIwsgvTShnUi3I7CTbFLo1AWH76WBA
S8FlCmAtX4kc363j8W3RUYVFpOslZNvlsEc6886favElBAccByWU0cTcMFePIHYQGnV4R24N6JSu
PFyTrxPyyWcbMsO9eGRIFVTjWqOQW9Jgt0O3m6gSSLYbc1fBg/FXJWmBJXGdUhhkBnISitdMJjuj
HdH1mEO0LUWCWKnucN931g1rp2c3Ae8bsDIBzWVsTb4BDbLJrN8MQuzt9Rig/0WVkAQ7pru8h8wI
+MjEGA3b5Pg4DzBEA2FdoqfArPz+rvFOpI6s7Hg6QDRrUcFk38N0i5yRDjCYllNB4kmdHsR6vyLF
9XqEGaSmeWWEIkWlRARnu3WVOzzAWbsfkC5luFXRIw13o2NlIafy/kpnBfT+mCKYXahbsfFmQnSU
he6+MhU1Oxni0q47WWw5ofdPMUaIu4rLoHKk7YzkTgg2IMEfmYJzhyJzvp1P07sUV6FyZoOTCqaj
widDQn9YU7Zzmtek4tQTZO5eTmJAQPnMUuc1cIiEXb8YQ4CUTplzQM3ypFR0rgjGq9znU5wXef4f
zNtpwfyCYsIpwCily/LXxBfXAAG6MwaBw1xkDdjShF56W9R5oa2Gnpafp00XgzayaAj426ghO5ly
UOF3F5itHiMZSCNkfl+Yt8c2IS90QMhdjmRnmt8s27p/cstGrBTuEkCAa1GMfANIlYW5XJoGVdxE
v8W1MedUYmnkDWY4xF0koBWe2sarHMq/o82HwtgROygdn/GoDeQs1Lg0LAsyrpRvtGryj3HVSyvw
Jf3nimOqE9oyfve7Lg9TbSqQJ+9qgKRQt4Q9GlmU5Jra/n3CrS03oj/EHXdwAgHFarOvv0LE3MSv
M2yyTiZWo4vL720NH72z3zDuu0ou9vK8BTuSAlWml3rt0x+Z9LWhc5yml0J18SFxCIcIrKIPj+Zy
IFTjlJZ4o4fKeYDcI9i9Y+rp7gYJm0p7de6D6jRsDXtyaFZSimRnikcgD4RYJ+QlVNFfxsvtwAv8
/pAl69o+9L3bNKi+9k8tuPN8PSiZBZtONlyezz/M/9u2O5RB+aIT5ovY797DNBGLDbaiGWz3h7aZ
57xBU09R2zgBYcv7Epp48+5qbcxcp/FK0QDD0vIxPutqo9h2N3S2JDWuWVLoZrDM9a09P5ri8SCj
FBOmi24PGFz7uwl+fqU+aNBzsORIn5cx0OKOmluHCyKJs7BKD23pjVzBC2WMksdTUEsR5uMxPFhU
V8BWAu2axXimsYT80xB8cEgPbhIJJvQjN/AXzVDlJR4Tjiug5X4/FJc15ys9ElhpVKDkMBh8z2Q5
u0+VrlBjma9AbVF93pXpZpIPToWcmfqFH1zhjQ8dwx0GMT5nySgPdETRZ0rKQxtWpI/K6UFEvf3z
IbY/hRFYZNhQ39Mumt9TR1tg+6yJbIr4vpKYQVY915E1P2yOeQHobeOFFMV3M1fcX3irklFlNuee
bCdZiLkULUJV8NYKu5NTA5EQHRQIyzHbSsfv1Hb6Q8PK9QaYYZ4YBfq82/jRYKIa7YWwnFOJSOTH
uRMnmtns0kV7LSZe/tALP0sDLSSZUEvzmgP5+cnTNfPWxZh7HNFdcbLU+XBFvipYBy8ld84zB/ji
GdST8/KzfydBVEWuHzzALZaM1NdAUZ4QkPSYVemXR0E/U2mHXEE5UJ35tyR+4j5gvO2CPjBvomBl
KvXLvhyWSl+HpJ/XDdDHl1nvstaqwEldAHM7kLpwJirSlodc9FrLwdp0Ap3+6OfBScOHzlWhMVL4
4JPYrB0zl+AP3cnBNE5k9Mmdf0PXupq4WEfn6fJtTONfa1RNqDQ+4P6DmuXA8ctRwFPsdjiYS60p
vYwKjidvFB/iLi+8tZxRj50CnafoNwKmdfCFSXyly64Zzjf+aO4f6FsrSuAth9kTtJJnhxgAS2tV
Szuyce6z6X8wAMOygcvnnpeYJ/+7mZEx97wi3Q6iz9j2u2Y1TS+WB8y/JO8ozKudlefIeBrHDFfe
6q4gHVNo5Q1eCpc5TjT4jZ5qKKgcCcHvxzNcXncsO9BEOjiLq3NuJk9GluiU3nnJVPPVndyXRWoN
x+EQXjykuU7jTtCtt1qEFMl/XqhBmU0nnXujwROX15fzSqzbuPUjxb7o07X/PAVq5ILrai5eV1Oj
vfNtpSy23crSIVM1n+umqlkwsJK1ds9ekLodThxA47kqxRohwUZ9qgS0SNBvsGZ16hN7ltmmJD4b
iCCWygxfzHffG6o6TfyrwH6oi1gz0L4xsnHZrCHUkqVt45YOKgjRzACP7DsbJAhNiscGv5GaQdjD
0Des/o2U+9OibXJV7/unz9uhlQxRbpy1IFq+oABkZaHKRwypsh5JsPFNTVU+JiKqRII4l7/kts5+
znnu3IucPCt1S6qy0zE4KmP1WWzzEZ+PooEdRTsry16wl4yujlSL+cvYl58xTz5az+B0Dk4fxJlb
1axaXWM3JFfvPfCg8LQLy1JYJKbysWCKMW2Yw0KxTeMwsjTmRpXOSopxFG6Jj3evEYkE/SHBn7Kv
MSrqaLvWddcXb+bW2b81JyZUtXQ9OOJiwTOW9QaowrrO0TfwS6SwdulwsxQ5WMUuyceobT7K8/Cg
DanEfKtrhSl4+BAG4xYe2Tyen1Tb47URkd1AtSGHe3hSyhS6yq6BV59VSn8UsGPMFS9KnO48ArNf
XJzNZmfPjuY3GBNGR/EBUOv9fvGc8dzb+yNCJRnLcM6SZVxDZ6FGJ2JcD7c0qaOLrvdceSjGPfQk
ZXQQDZ5beDHHWlLA+uxO+OX96gDq5vDaKoVczD/IilqZgIb8kqSE4xZ8iDqvGogAb9/11SygFZ/t
eRG1YJ4HIgtQl8GUr73ZEyOEMUi51pFYDbT0BogM37XQxv/QytCL/d2DldKT3EPaap/qUwNTl+eA
E41WYtbsOq6qX1Dj6ALlJBoT4F0IqYbNET2z9ARa60oHVesHMFjAbc0KeyVdYzbMotgR1FX926Gl
0YUWohXOVo1hyzXFP23pxo2XtW+Bfqa0JB8cPM6bZ6odpxuuw8Xerfj9mv5Ho0QPqZKwOw8caQxw
HmPwW7zx6rHxhYZn02nsdRhLpebeszXxTKwL0GwPDAGJOb16KrhTWiWkSIZEyIfajnFxmlXZIiPv
Gg0uTKyMptNeVLxje01PCIIoATdJ70Jz3+8AG8AYk9XoxoGvsASGg+CUa4FdT2R/GokdHmqevEjN
ZNqh166W9VhlifwGG8JjB6SsMe8NgT0tEYIjpDcag45NI4yVxJOa0nyy7AwxPSOfwXAtIsH/mN2U
JTGzKZqjeUoZerrHQDG3EKch4Z847SD4ACL22itUZIE9O9Ygk40pAPaVIapG5g3n57EpHpZ6O4QK
f/0HrHG+3T1zBzBEYdVdOH6emoPFaDs9KOcB5WIRFtFzURZOQi57FMreSc6e8Vz9SrPA+i2ath7I
kFv78c0OcWHDf+FiQyGgFLNkQy7glwfIUmWCHn0RdgXUfA7xvNg8b2WIHjXWvwYaPZvlYepw9XVC
6mIRrqXhaxabsbMXylqjMi7FGIQs1PCrPFyVWa1mXCAPFki9pAqsUROV2VQHcSw7UxbHLx5E5fxw
g1iJH5aBbIkqxqI0C/KHRMj/J2BJeU8JRr0aiamS3401gud5THatMj7bXE0fi6nfvzohIL1ArtLH
4swhAScrhT/XGQb52AF3x0lle29B/Cf/i7vk3of9W+gtWEYEXxRjAZfjkQVDi9a0Unh7vzZQ7Ork
cnxYzCGvrjkOJpRocS5XrmYKG2OVKML8P86oRB1p0woxkDlLaZZfX/QeGPckBTj8fAaa8yWvswef
e177/y5KH3ba3eZXV85oIGOzITOEjMHYkGVwmvB600j4Y/AwLFx69X02BzBgejJiXTWijk06hdjL
Vx/dlb022zDt24LtJ94QCMwS3wl/BB8kXuvCnDSJ2ilUkxxTgTYa+cjwVoQsI4hK/ZQrlKJC8e8D
pjZHuOXdrcusbWfVSfC3dq5+ZtOJy8y/ms66Vsp2zVUrVTbDx9u5kB1sBkh5cqyM6OcbJtWqiNAV
YueF640aGIL9P8RO0UzzxwSbhO3nNJp8jVkbfBL/PDzejePTBHoRDhWY+eGJbLbG6Y1NCq+BWDjy
l6CR7e58YqPLhMqgxUERhBUHpzAZ5RkQJJqGE/0G1jO5a91PapGZJ8aAIW9RRc/vg1i1RuC7PxnE
onossDzegfNwG52yHxBIGfjaiFtWeGMTapeRnQn5wl8QBT5o9mLhUyexmY4Mcb2IiirYo2A6Tz+T
4v6Y6/B3cMFPDop4pJzKG68mQ9YMdv0o0HXswECHhXOeBVXPBYWBXPMXnvKKQC5zDUMaBwL5DVoW
8qrH13lXw71tSYL8sclIvgCNNgchu8bqUQMfzRRQHT6wFjup+voP35OSqS8f7sm75Sh/585dHZSZ
rhVZHZvbweDtwxEQVOQ6q4XbUv5vURr8d2IXZUghuf/ZRQeQDAaj36SPrYwd2VMe5F2r4ABJJ7+f
SROckjrhYDBDB2um/yVqxcY88oM1PqjvDF/f60Vu5OOp5p1omcA6DmDc09xHW7HKJUAoqmZ3uH6h
kVCyHLULTLQOUz0H+lCtz2569ypjJ0H83xnSSeLtxyhVE6PZX0rTpRXvCkIZTmhUOPnZCUo3rvxw
XEEhv47sb832fzigh7kJZ02Ns609bpxSwjd5BIygYh7fL6rdjsW5kKPcHc1Zpd3USAjRNkfYun+U
wLoe/zG7ra7mLQj6a0L42UC6yJlbgPSLc8Uw5p/gFc/VOvwI1ZNLn70MwEERN1gtAHcSCaWIBQyk
yh70rshm6vJxBjYZgZVMQ7UqUppkBAaLFardCWdIaHBCl6Gw6f8Ck5JdNRbeZd7oB32W90toBJh0
p6dQm0hvuv2+Y8XoxfrU3S3luckqRbaCnsS50VYu4Bnss9b+9aHQhYTguEnEs1yUKcHfKIIgwlqw
y6pFWCD3IjuhiYwOtKGv3dEFngdTF1koc9s3uaCD2boBHIE6LAWvBCQIIq/Jf4sUGBxCyisr1+/S
tIixzlMYdQ5jYJjgao4XxrMkTSq8ztB6gNLGvOEto+/D0dTiuVfssScq+oUEWNUH1Vlns91Tpojq
4EdkYpzgedgzirZqLiv/tlnpvaFTWc8CWLe9ki5mayxM/hymVVVZ3NtXWHe4VbMjKBmlSioAGs4Z
uDiei2nY7C9jStOnTfkcdWpkxnFTdJMGBntTUEWbY++oOGF5gqV1Jj7DHyLCk7kRovNWCIaYfdHK
3NdWjBW7+3tc9/yk1acq7BQSZRhP6tmJFTiHVurQrYGmV5omc0Iq/bnSFSeMg57TqIWHx+E/VLpS
JcD5Dp1zBPrzz5ZldIUOMQK4gSLU42+zUbOxLLRSlUIBrFliF8gNea/+62ECtXGKkM7rrjiiLzle
CJVibq47Ol+pAM5faqm4hJ/aFW1hrHlBETlxqrzd0XkDrDe5t1jzUE9phLUShz2qmdKY6JbfCaJ0
gssnQTF4vtnDHfFZdP2J99rDIE+3HEJxSns8myfSOng2L5xxyb3CCa6akBn/iULdGyzZVOWpFVZt
qVr+Rto6EmDMcCGOMKehYizPNIbntVX3k7fSeUXAd0zb+hLHhSwgF3aKtazfM0tH6eRG7TjJdmrE
MaygvyXH+1c+OxV7rg88Ki3n8Sp8NAiZqoZKgdIiW3m3bl4RrMWbSVG9/MnauitpuNciu5wJy6Tb
TgmGp8iZLTljojaampisHSmmBROjzwmqRTAefSQxdkoL2M1DgyAQpghoPR3IXUDYoiL6FU3h+lJB
whfmc1InjFUjLUKZsmApISbcxEf6gzSnXJZDw+1xzBYtq+cQs4lhIAHRqXVB+17iiSz5p7Sq2Y3x
5d8nbGB1LUdxPHQysJq8L0CJZjSeRX3RlMqg4jXcfdsivqQw2+pj0sQxNuLLeS82575+Emxy/Twb
uDBVIcLM+kyPVbUv70FH3vp8ZpQ5I5Ofoln2xK8GbbpRaM0Aw82su7l5UcsBiN05oijZXKzAT7lU
/BYgVX51HsfN2utTheQMZi1H9D6ql4byqSRQL9WRV8bIrSIdvBI+XtfU38nJO89SABBZkIVCtfB1
jrdNdUJBaHkzqNyRY1s3b2dshCHifNtwzJQdTP6LvFuheU1W5WnQHhMO0Lkr++uf8cP14yul72N9
6hV0zJDpG5fEyglP/70EGaL+zKY3C4njbwMLqdSYbUo8KZjeodzoAhwX5ft+UZzNyK9AnFP5iPt5
Ua2VNLBeZGDjUwr8y+zqCEBLXAu4MauBgGAVJaBR6k8DlYIsgsVRxzKLlMY/Cef4CcesJdiDPAxl
/nzCm2PYVb/q/Vi2aWuYQh3QhWlOu+MAeUVO5O34rny6XQPKbpKObrFNVkki6Uo/jv82U8hFU+rT
GWtEgKNKbENvDIpadmOVQAGbuj3LNWCxa3AD5FfdZ8nh4KvTFbQK4rI6/UEzkMUsV4E8qUzZzpX/
PG6lPHG/oeoHV4LYccY54Iq5bXD1kN0BM26ej2A3NdaCm+QLBkNQRnxeOMcrflxfYBkz6OnupOX5
mxN3fUU4Y9DqiLfUBHQtA4DndTF0Jp3EcRb7eEQ9K19sCBx6AMgBhUKffIeTUKDtVr2TXWUJrys5
ugYio9JMBshgaIF9wxYjoUQcTV7nnDgwnOal4z/n/1CfQAUwlrSw2fVLqg36qag5+GPsmRYyQruA
k5nsBCU7Gugyba1Q2NwBnaTOay94GeOIJZY/CxhIBt//FZNAIUWohwBcChP+y3jJizoS+pcn1aWQ
Z1wIZ6wem4kZpWz7acsvIXh4w/R6AX9qoGApRvT1iT3wA11mOf/BzRWBTCFBgR+OF3KbcIfVBAPE
b1Ju7xYQkUrYau4BXbkK3pcr+GIezuKYnggFaRf3AsItHTho+7zld14LHQ4gK4dy5PjgITAnwPN+
mi22WuTd12sHZ9Hixi0mnAQR+bAgotLO4caQJM+0wiYc5paJc1NmXegJ6yHL7vkz6siuu8WWYCJg
PRAg756ZwOJharL67y0brRCWY/9A/rNtrKDxlK2UNnzI69ukWz/5LoUWHDYTbTcIuloOFosV4z4t
PNRlEtYpIljSdxvRCrXKXoZXWfEzX5tJAm1QFDGlDkY7Bnw1pOy//I1Kj3QlpjylWfLqcJRMdyXC
SD24Utc07Pa7JFdxDJOxEFCm/Od3fGQckt2gq+1g0NJ9yGzOEx+1zFNSGQyHzsYOLXauDWumVBH6
2EZ9IEvGImYcK2RVIeQpQKAn5vCixkttfpug9r6NRzDR1AfgXZpxiLISudGmZ6tqZsKTS8Q0QbK2
hiDH+1fujtWGojRW0IZvEHuxPSiBMsa40HPiEzM17b3FYi6/qOe1h65FXT5128QNv6qbkI7s8+pA
3ShUUxJ4P0gQ6jIHywSvlDC8COJAexOQRgrW8SzQVxl+YO2EK1rqYaei6CVNfhZjI6F0vJRO/1RW
DbCzrCH83exHkCxsOKilLcLaWfOjRH9xmg3PK4Rw6CSMcmJlVXD875w/h3lnjhLDug9krMQhSFn6
LrXO9T0skXarIOyseYa5O+HfUdLJgzxofldGez7bC162iH81dnoFqOofagIY5foEG6F8Nw/1oYI9
8uN1yEzoqgu2DciyVDBkEP6uk1FvJmKWB9cydEOM+CS3O97YE1q/3oJRr3i/guGPbsxVvoOUXWtd
QSwFY1tSOWE8HrEP7SADLjPhZnhxg7WcUOUdZZpEYyTgcGdioq6pzy3gb4c3fHoz6IuKBxuFRSHL
oxi4fftjpg4gN13DnxO9Xi2KS+xvMfxhnl8nOffDg11Xot0kK5mDDq01XXyJQpmxcpZE/rmMFSO2
ZDzCYs7ayD9QGBdUkd5NRLVOB4oEddMUY9muNypg89cPLeTSvGC5aD+5Id9HCfXpQck0FpvWANcp
eTUbydrAzN0h9jdTQSFyugI6ukEO5bJJSofnCo2Bb5Z4wJUq6Udq/DJv2rPyF4eZwDGl3aBGei0T
+nJ3459RSkjCWXHuC9G3iW7mU+6CO/mx0qGwJdiQQQhVdcLNqBo5V94/DCpaIVOROqY3+pXFrGoQ
z5oXvai12wQHEdGcrZMinVc7O+10ayDQqhHmiZuh37S/MkfSfxDtuxkY+2ccBBg5m5poeEfImVwR
/7U+V/rTHMZNBsikpiWEceRr4fgpUs5Q4wCegOWWqDJBzz8B4B52hMGgCZ042DsZRY9oR9vk7QYV
s+3fYYGfZRFfjjoyKZngbt27vffF5dixKoLGgIYKtgLHQywsVub4Q8u3BgwrHpdzQBtU8SMiGS4/
FkAoFL4x7hrXD73twaC6DCg5hYvmBpkV22ewbCafPvBr7BlVTaE+mRI45LGe0aRc5sZkA7IVxcag
xXQSUy/ujLQH2UKuHqN1x8ph2IzE3BF1UE6RzJQLF4prS4/cPJBy2yJQXa/jDWStD9aKAL1x38rP
7Gpk7P6A9jgIDodUeonGS0R5UQbYVVqRtPenQMhaXd4WN/Q4nDBiLORsNNkM4tSGLBdlKg44Jyfr
lwqgT0p3dEfd22ths5LdlvCSqBDSr4CJ1wdoAlT57fC2G+SA9BpBKfIf1+HQ2K5H5FZGvbxUSjAx
txnhBJhMb9CZBFLduFnboCG3g3mD4xhcNBMY1Aen9oAA6GPoAJY7TJJ9rUXHCpnn4u9BkaKub0ur
EcZmrvbtpjUZ/efCSqlnqgom2liMf+N0xvqhunfEPA7uDC85jNxMDevXoTc8O06K4YQwd24hxYzN
EARM9of0ugKTNq60YHnPmvlMIhoKzqdseZdk6vVK5lgoCEZbDDkzcvfT0U3jeCjJC13+l1nDlBpt
gg3tMimbT7y/fdyO+SbuNELoL+Ry4Aba6117c9s2Ljf1pMdme/79bc3DyKe+BZSM3E/7v4dUfUO9
M/uujtOB3oIWU2+ax1vPOFVPbYG49ekcK/fp8b9Uzp7+nzvxJwiBhYa1+we6U7NguPPaVKEPr6St
j/esWLMMupoty2LCMU8eAo2YIIAG8L/lhKr3QXec68MzfOXIv+9wwKDVkDoh+nka904aQs7LF8UC
zhMvDKm3CtlqUj/ZekgtHwi1wXG8SdQr/EwAbrle/l/glcVuwYjDlLVNf2Xg3CLuyCqh0HoL/V5U
9XuoMp6kQNivaxXCaEMcUZSACBtiJgtKFpSdJblxJ3mHaDp3Wv4BFQDrAhVD2ErKVrOv7uXAv/f0
MaAH5oxvSyTfNeUE+3cHRSdqGQuI81n0ynYnC3WAs17EHRfmVXypUgB7slGz8iGVHIrT1nYruNWH
gjU5LWRHjYhYuVmWMGol6jDNaweUcaiNNvL/YMdizUBaEe12UIjprcwK3jlx72zH5iR9ewuvyGgz
OvNn4kFb2TvC5odkP7GOxgROLHkPcoRlaVcYAqKwbVgAhPSVHs8o3SKk2BzmA/A3XMoR1NIKFYX4
YCiNP2mN3dx+O/DKpr5g5vksDznQqB4SVa5Y1XWy54O6pMF0GGHfItpxe4TFb7CAV6gLhYBY4gSq
7QlLj6GWb7r92zzIah7hpKt0sYH3ta9RJf9QFKyPaz/xJWAiQCGHa4pmp+D/95kZSVx3f1j7Cqgz
RR0oUCGX9WCPp+JyeWI5eQNsBSnY3kzD5nobqobUkr/zpWrby2YJbOjv94I+VCBzZ6vBFA6XNhTl
P8t+ZgkVg53L54BzzzGK+R8O4lFKZFVe+P3c9oykt1leSAtK1MBd7tGe9VcsJXITxFp4Q31mn8aY
R9u2Xo9X9ZiXy7N+BinNuB12kFyH7weMvi1qd2m5nGKtNWUUiQIJRI3xNFIGr0/wER0x0A2M7x4C
WRt1EvyEvcUoMFuWSqUbpPcCJvPU/2xA+PomGozBVuD53U4vpG7wIvgp1AqXkoRSK6xAPc7A2uAA
J9VoOBRIGzeivu7NRKvlZxTg1o9VAOdhVvU/EUOx3MlcOIcE5XCOag85OZw4ngBFohxngszC+iEV
SoZb8ExVAeVXKVi5V7OOxvO7qUr8LxBkKb9smz7XR/WlhEF7h3XwHKZ+Mm1/cEluBBdrM+w/VB3e
Z9eKHqrHctjQfQ73yuFom6h7WGvvdEBu7vLRh7MpMf+ezSZg3l57I3fAJzZ1sEj8Fv1WcconL/3C
ISD8Xd3jo004Y4KX4Q750Fi8zgi0lk7W02YuUOyNTAw/otKf44JqWIPQ1GjhsMZ1HwQZFlEgFdnm
APu6LoFBdKaZMSDdI0ocvk3Bzg4DR/3eOPulGkklL19K3N3tNa/uxoLfewDpRCHjJ/kKBj4hI7yE
0JR08kyrMXsycZdl2pT+4qlyuoSDM21cMgb9njjrGZV86Plx9K0LdaxNyEiIg6jGU0rd2DgjcKVL
9ffd38rujVF3tU/JCanPpKBDjBiG7SzP7QbbQJ+ukUeB8QOaKM/b48zoRHYJNDWPcS0DnTjwq/8E
ixdHvpi0dUcP8Y+bNuJykurj857qwOmowVRifuQgchIt6Q2D/r13UnwPA3iatA2GiFGWP5eIEt9m
rXFrJQVayG8RrSZec2Xmn4AKQBVTp5P7ecBMLPYcaaRTwHHnQ7na7cIMQdiboV+BFj2Fu5SxSkxI
AGjX5IM6xMKcexVI/6yojbOJ2cgPRHTOK16tnjKlrfjy0k/rrqlYH4/Uez9HKTwRxS+waU76Gl+J
NiJIMFPt6ZGvh2qKektEXJS2jqYNMk3oFDeh314OP954ckIGS5ig/Gd0mxC5XnxtuaioZbOA/jW/
UOod7zT7EBI2sAm628Sdltel3dgx80iaEHKpek/URg1uIP9RZpKxOJGoDArn2oVZFp26BbFQtPTk
yCDd6uTQd43Jec2pYf86KkxovI72VYYZr1BUUnlU4Hz5DWmJe3sJ4gYKfUs5Wn1tcv/zHIxhub6w
+gFgXSxmfAktsVd3qvjmtKTny78AXyzp36nGlHMKx8ktt26r6WAvFJiR4M0mHKh6ZcfW+72cOiEs
CymO4ATB2j9IUfDKDDn8os20ymbf2pLaDD5QHI3BcfZIlr7S5OQU8L925+JOEQDW2lHirLRIgSF3
9Px1MlIdsi5aasVhUZaAj9LefoefxPfIhwyRSK5ambX3om9GtXnmjtiFUjnshAsnIO/PWYSNRn7i
7QKz92KjHFapvhZdveMt2Mms1OfTQZ8oeynhcbxfpyGgeJ6I2L/9DB8CQey/TXGHnpKOHLMoLoEG
PhlNVXySVJqMjsBk51/u9y8oSdwLjeWHl4iqrsh+97KjZlGMLi6KxDMUihisD1qJp+G33lla7LtI
wRJV4roP7U7qKZ2Rb+k9TOT/K6IID1Gq9GDBU1HJrWC1RlrysqZwhhgpRP9jS9fx+x/tosjLizqJ
cOcDmNebCUsNKogTAi2vP8SkX1y82Q0x+o20PDpIqNE+rLF9xhfEnO8SqzyUaEAbpXo81awUdLby
bnQHgmBsqMfiExejDHzUtwQL2noZ87UG8m8JD+09dBl4hy/9E9+TlLVu1sZ4gq6YyekfKnYBKUcX
+a2Z63kdpMYUwGWZrscqQvOzhRxmhkDVvQGcAkg/hJUtRmmG1pgWF0zoR67q1QRfP8N/MvLfdHxe
ZrCUTX1N0Tqn+ta45/7xJaQzNlfmDeloa8tJcOeBVmGKd82X5LWqqxdhZmaC9whlpeaQ7vFMESj7
m/8IHrs0TWeAqoPXBUL6UpzMmizTFXAtc11e0ovkEz2DYFHKpve+C1T3cVnb3fTQo2zua19WWCkP
kfLts9pgAhbzaknRfyNfay5UoG+x9nhGhJJbgHEtvr92wQTvu92DJ2YtswS8j8cRa3xpCMRXQclA
I1usf2XXAxFS17mC7esvUvBITWdwGz2deZNorxPba0MXkHrjrCZpQ6D0k7t1Rd89bm7GIqJvROro
GaVF0tCsbtFNPKmn+pgpqt0QfcDgLfkToXC2WOQ97SZzjWpXNF26b9fPwQVWAjW/snht/bUkOFDc
E6qpa9nmT+GyK5zxrrwldAgNfQ9M1s0VC/5JYzH+Q2H+U4m4VWYdO2CXzZq8yRXfysmW084agsyS
e6QivQlCO5WCFJklV9oZjBAxajzCEUEDA0jyYQa5Lz7BI3W1g1Gj1n5VcJGGaDTQF0uzSa71es+i
GbU4GgQmoo6m1hAp3eFpY+TEbPfq6b8IRnqvw9pOPml6D09N2FbbKelkgDYrQjjIDXDvxeoeiVAy
Ij0EtNhehOhgnIzaqxYtEyUlY/r/0mtzjqYbHLPF7XMHSXpXCLDwU4uxCOc/7r4BFzNcDiuL7bCD
pnuuPSjzOVjBUW+t07nSpYM5eZVL2V0wK5vOAFkuI3qaCbGuowVXWbuM3K7BIWsWCiu5MDZ953c1
mArjOyJHhpYyz88AyEHQimPF2Jfqj5zC8HY6Ugqs4oVA6nxLiZSQEj0MnnH0gx+kb+LonTKNnjMG
gzE8vCr4uRhCxSoQZV46iVcomMVMb1dQCde/SpwaykFGZ7LY/omq+QiC5glM/Go9C9CrBQDupSel
uW5qtzPGO70sYiSK3TpXjrP5V8JNVxLIxZ2tI4qYAwWsI5Qs7buDisvgBJnaC1ESajRsamqUhiNt
33pGHM9p34vM8uThOAJ7FIKxkaNbKF6WvlXQKi+38JNwcM3IvO4EARc1ZmfkhzAuEQvmCguL27HV
EGrrj4la7dbgFMzvygKJetZQEDUIrWZa8VHaxoD4JHlvY2jnh7NmLNFxa0V8tTeEdTT9YiTqVmr9
t/hR2sjTJp9iv/0n1IIoAdkvM442oNwdvs5BEWm405DZDPeWdtmxqO6x9JC3vMVBD7xW4J2UVdVd
nSaD1HG4UMoXjveReqcdY9mEtd9TJOvonqzbQFzJf4wv2o3Y+QTQhYo9b0B3/odEzUQAH1Ea7X7p
3CRj5fYnZsaAOoha6pZ+V+KrQOa4zZBL2A3QpOJX/eqI2CWbXmqk/gdZCuLf1FrVGmCfCgvcQ3M7
GxO07Llo8LncR/nN9LzEgOmw5JG41h6mIcgShlZ8lHuEA6ouQx054JIvtc3Bmtew0XkW3f1meMzT
q4bjBbUIbogshyNQ5XwlweTyyCA5/U0ABn4cvRvkwwqhXGP4czKLNb1KO1sPsPmYJH9FvGayWmy0
KDl6Jfq1tMz/RxLqMneYb/2uGrBgRv/GVMCi8RClD/3R8HCv3cC16OQo0ekF3k3GBHHjRXuZq73J
wBCLmWGkSduAP2eeWUOF2pq7cg1HN+cME4kmnqSuzv//JpGPNgEK93ZNWeuJJJn1/lcm3R8yq0N+
bgIP76W15BypA8eaRIf9MgjHIsiKquJWXldSFRBCs3H7W9QP5cssPAGMfW+KjQSKETq2gtVxV1+a
ChuwQ0XsK7QeVLDBZUR5xf9uiO6fi6Cf8BPwsUUEMXADfGEyFgz6IUaJb2ONTphYYO/ciIXpuHuA
3rnhT8kCNidZac9xZEAanOCo1pCaoFtaAZDjBeyfZj6PhIx11+QfAbeBgGNMcmwmfGE6aOc/J6sT
rifEXqFzj1ll5pTPUp3CHMJJLg732yKepeQt+pgyZASU0ZlHvfoL1mkEXSkD1cJXpTDlR0Ytp2pi
aOHK9f2JCVxxZwVEHhyaTvaESJSV/CZDL2tiOUYRHey53Q6qPFzbC4Q7Dc00C5L6VvqrDljmCTcn
diKJas6Zx2bzO3mKm4GPb9fxpOuzrvq9TSF4XE+8mS56NQCB30+nfb87uEeHKLu2LgM8nXPjA00J
WbwLnF9EiiUGbu1A5wHmUfbpERgw9XX8nO4l7IVCDwT6d++khtnwnUdjVi4cP6V06mZgv6qsEM/h
eWjK8DAFkfqNrdBohE0cT94nqdxNWdw4r3bspHQuSCPdMeiFylz0/lGahIXLkUJvDR1eTN3usM4Q
g0IXjil6i1N8TPLpMDL+EhVvHy7yqmveaael95Z5a8Wr7dOcc5peOrTvGCE+mD35e+IfsY2fSwSf
gZseYNC3GHulHoI0fMPAzEDkVqGYfABOCMjUilRQcobiAuReP89sTV7GTNeksC6BdLAmj+jaDfjF
Xi1UEhd8X5ELcjEYXdn7aSDru5/9bkFzM53FVxDPCx3H5AyXe3sTBUFu5d25ege9UunU2kqXIsJo
pXqDtoiw1GcARawlVYCDN/uW3gi6R7wvfRfdqlDUq074omYKSD/liJqwrUMvpVnJ+NQbJuWFIDVD
+buN3bsH2hv2KG1csoBhhZfZgliFB6fkCJWaL7hindkuKxlbdb68UDbI9Mc0wQkPWZ8yoXNsKb4E
Garn3Ynnh/vUEYet6KFcx5vr6SsKWIOLAjEh0kIg8n1UUH5UKqarun+p5/3hIxNtmb1K/wq4na/+
C2FIolLci/7ZI1tWnTsJ31gapELlkAajb0nUXC2FhxLTQP3BHF50clyRLQAGScA8qfRGJDWqhTp9
xucYDHz5tqYKvWiJaWlZE+OSGg8v3MyR6bFzUnfVmpgmW9Bm+JQQFP7JTz/f/3KiFU7ZTUgXZlq8
UUkL6g+htkmD9VGJKyx1c6ebWAcVCp2m3M/qdlgsycXacXd/GTtLENY6CbNALu+KM9LdtOZgdjSq
JqzegqtPQmLySf6PA3aX+fkVDxwAPs9LMNAQXe0N2MLDcO4g5PmGX8FnrsFS5WoYvdw7sdH1NCy8
zMutnl2VqsMdoxwsuuFhFPkT6orOx14LAOCW43d1AuMKd4bDRqY0jTaGsZGoZM5jc4zZpT/x2nZc
gGIUlfBgPy16PSlP69owAgRh07GNHC3epWaoB4twRL6LkZBEkZXywzmI1SXEoxe1Rp9A6t7J5FdO
/zrpfirH5+kqM0aszIvTWQlvuPUKEKKZ/u7VSroejmK3JpxKEsWXZRV8ndf2gOEIr0dJIl7CZLG3
PoBiRfgzalktprj1sizBJ7mVoa8Mp4/Lj7T9f0kl0RGt5PaiJp7d/iHD1vxxwJW6ICezHvk0MqhU
7JzAL9iUizeqt2vtd9c7jQ+C5+0gUDI1ipXqypb/D12FDvEpLyYe5ILJN0BneHKc4wXmugsdd/EQ
bL6MkhsXpnb5PvUlfU9Z+OJsGoe4SWnP7VqcwxqLlWY7I9tpit1FCeJv3KGJ8dRnj5NznHJjWB1n
oCfrAdMmkPWMpBBiz5RkRAh6dqvQCcIVb1LKsvmVgnfBzulgworrqMy9TxwkilrT53PpK35ZlUcY
tWXaOUFb7DdBdIl0I6XQUVXb7mD4ZNU7ddDB8HX0fLZS7Z4fa765FTdevGnj9buFhF0Cxwr0t9iO
XojuZf8pyutOSJSn7tNGujD8S3Jjm/R5uh2ACcPVKbv6uRAVWi+ABfJA3tNGAaTBJyl9qBwH3oww
/cAzsqrn+9Psb5fKadlmdtmjNTqBL78r0NXgLm3FO7QlHGvytlNyVQFkZaI/zgQcHv96+VEQ9CgY
6q5zTsI013AixtiZTsrrCWgtBfPeFqambpHzOVYQlh47AQ8CdC899P1vdZ3RvYB3GWLX51msV8y3
/f7owQfzvVU/7yT4SEGYOQdy2sKGPHxDgENHoIDOx8GtkhB8AFzXISnrEDfRzacDWE75mamSylQ4
UTFHiGEwO7nHh28TyOUx7QtW2be29U9wXcn6+w8LkrdegYIqyf/OijMOKwW1vtnRWJpgGjsYahYW
zLvJcbXO16VJABiCZtuRcVD7a5tCV4K8pBbXNpeMOzLPd0GOxab42+LmwtOL90V5FZVrHJGGByuI
VUoAAdKhUi3snjj7B7qqqt4sYbvYEa/dzfAsm7yAW2ngJEzUXAICB9Mksu8k25AgspINZkJZPny4
QYiuVAQ/qYSq0AqaJ3FPQquLNePy+IwnW08jGzAdJBgGtWoBs6RsU45/BQ5vTonvvpL2WBjdN+ff
AtVQC32xXcRbLfld9iEEaL8zuRUEIPZVEsTTJX3mih8ZJtFkfTeXhinJOZGaLImD/hf9JnpbE0m0
enNm6dOVtQokoZWLtTzn3XGSs5C6rqLZbZO3UvUEipzoW2tXcYgvMfapUci1ttbfiTPzONCylzsZ
SGyuoCu4AUxMP+117BZRuT7AjFVt/3H60azv9rziUlAK40PA+/2GASmRaWEXq1ThH9LQdoTIvILL
0GYn5n7HRq9+jf5mY+wCbV28EUcZTAxrivNNSJH/4YVm+J82sGeSP+6HkvGkw2XpAJnjlqqWB3Tu
A1zuBVBpVauNPXXoV1yroI8uEdA18VLbCLzNAupkRa/uKWUmVD5thFAYjga2NquIPjkBqz8qD7+U
s4Tu8EqaZFLTl2v0w+NaPpDZh4gafZ+r1o2UQmaCB2lRZTBlrrmakdYCI2gJxDqiHDTkEM+TTGeu
VJlajDUPOv+81vDRjmEDUSpTJRN8Z4MT6lfYoojvcOja0tpzwJzgqIAMJhXxoUQkrVBxeDsgF8x/
eYRb6tOIr1v2UwRb5KeyLc3NclcAEwfvadTKtoEOohdG8SEqZIjFy+Su/qaMCS1T2Gtk1aT0NHmE
FI0DeaPc8tw6lMo0AG4Z7G8koQcEcf2GHPrbQ9EcSWBu/S9c3KN9W6mBkSrtFpgFjI8AyudqHnNp
JSrvRpbwqBO8Am6nl/NpZnEaH0usXqOcKQFJtN3gTD0At1cCevMWcy/Rr916UJEoIGSfyzXhdSR/
zBkXX9cnEL4YY9MvrVF1cg4FyV0nTp3MhDT0Nwhwg8SOav9qLhP80PsNXayoA8fU+12zqI15DTyM
0yxByhcQUblA/NrzVWY70+zi9CPY4GdFFvRvaNIr5TR24vaTNZOTVcY1EOE7hsmwMR268GIPjbZv
tCrktPiaVZ1pJ8C9R36YPH/CyagnyjjwNmHvWNKIh3fmHrQzQwfDzTjUuziPTAH1H2b3eViSLxdj
X51vrVYW9RMwDU6bG2h0eTKxCmUII0tnEpbe2LbJs9G6IJA2y6uMijLrx98lUnTEZdyDHSEIGXSB
XzMFJasMZoCpBw40Ql7mnFcCi4yMuAiDoo/OLTk363Xghs2hArkQpmpH36KQL5wWXElaBOo5rBny
RZpOI39xEio0T5x+4VzfxMusUH6wIEXv5tdV9592UF8CViypaAsCgL0Ehrky/Z0GJhoUPy93AYp2
qUxOG+zGTIbHR3Uug4EZ3ZEbtexTMd0PGFP2v4hswUIoM1Szdme/hUEOPQxSr910jfwi7j69rdIq
l1u1E7bq3lJ8vmDZkANn+JMbluB+vajro/UB2zPGTS9PNBBoHQPujJQq+cLWFXgYj/FJ0VVcQKWJ
F6VWB3Cgxm5hESKTZxc8J350dciV5C5mkvhzJ0Bmyut29ZErH0OcCzl0eKvt/1xPAvvJxsrJYEYb
cTy+EGBIXlzrVmcT5FAdy4WZT+pDisxbsznU49smhsruUgJ1mPgKDlcmC3aPdFkNdVgKLfe9mQqL
GjyoEUCKw9eKNwCh/ba0qXK7Jx+/7tHtz+sKxkHeKbdgud+yzPxETPTJdahXCKLGVRMqLlbCnH4w
JoeWGgiDLU1nOfV5M88rJZuKVL13OTjKsY7hRzJv/tNbEUwujBDdd8QqvOzPig0tc8b8033l/m4p
KBFTP4CU9u1wE269kO0cnAtRMNHBjkFFZdW62VrMu/GheZRgK81k7uFX57ajX07GIouLLN9DkPY+
KPAQIB8KOhiAOrqpx18hzuRf2l1HdW0Bc0enX2vBq5bQ8KnCd6Np7Qz5rBa8vT59p9FNdobR3dkF
n4CG2SM6P0AK/4DAbgkbx7DcDxnGAUjsuuJbVdnbpPlKJ365j3d32Q0wGMFUYfD6UxgqnaDS8uXt
IFCyqxj3OEmPf7qAHDtfnIusJHEdJsbxdzB0A7Vfkb1yWkpOzndhzrR3W+pAPLlX6i2vavKGn8Px
PCc12DDRmJL2IBmSqqNZnpj6vSALD6LTsut2kQXAWUGHuk8Ys1KMPwb3Py/s4xcTyzDiGEKw5Izu
8+E3XJvXqNIkzAu/Dw2OPIK/M9LRMxwUqRhqKe+ADecdypUVH4okBUjkvpO26BUKvdGAxYDUuEnS
Xf6MdPzhHO58ApWfmgeeTXsMbX1xDjiXEPkauDlX2wmSo6MtZJwY4lVLzsw2QwEV40556XM5wwfI
JMXzcqQIlktz13YbW3it1gr5M4Teqgz1A1CyfcDlEqC0PAB2DMvKV50KZ/pQWXmAf9Du1H3rYZFb
MBpOSi+ioOHBTQimfn/f6EYBhfsr0w1mggyw86YEcNupsFOVX4aYzhYDtI9gwJF9365zRuCYUVL9
Ts4lXZLoqery4WqrpOs2dJU++gpDoI7Bt+IYQe2q32KCtrjLp6Ydzr0sXvtZXgmtvk4r+bkCL+La
RNB8t1bCPrzrmrhmrBq6oK0dLiPasNK6ncJD93zkCD3LsHHxwuMIyK/KlgH6DipagBZMfsijAd6c
yGS+HA2Ycr44hpNsgqK3DBm1zjRjpVNo7fmpI2IJxWbrG6g+UAhHhRk36Plc1oUPn6hzbbpIQzkZ
K78w7LQHXrGz8TMqcKKkpeU/WyjQCsBOeozkU80YMWYhxyKfAYGiRVYcaynHp1qdtoCFStMZz/53
NY6WkFtNJAwzQNeg/IoPTeQTp+6QD8P2E2P9ULI8qNLeHeRQqBiSHfo4Ydxw2HsC0ejQQcEzs+pl
UvO4b2v6HmtJaoDZvh4x9pA3hKRBQ6gzUShRye/PG+Pu3hz2o7euTDmGDeoYKU5yP2YzLb/wZhNu
PoT5d7aoeVRZyM9N1gK/ppVa/ijJ5rfoKdpJ2J0xdREf1LgnRtb8n588H9plt86fTyBGuDeTKlzf
j+Ho3wQA4PEh8artyuKNBdxZnE4FIh4gsoq4kNxGPadjC6Oze9NrvQSuvEjbwsEezJxkHEShndum
HI0TC45Un1XHQGLPna4Zuu72FTlcCAiD0QHUhiEwAm9KOKwhPUcjxbGbe4DrobfuBBSdZ9vj9h+j
DJqUhOQLyof7SIpCNLfuDnaZ9k2he2bj56phlH0RzUYYvxRKHw+DX3NEol46/TtYwVI64/D82og4
hi6o/aCcGKBnqLa/EMlNnr/p6WoU+uf5JxS0ufmOGBua/OjeEkSizs4GXbIKVioTO7BkZJMfjgFs
aPuDLxYU6tTfS41usbldIP0qltlwqzP0xnGNt1ihxlCyyUM+qYde6wa34dSbJZEh32i/zcWhRJq5
N/z3FILMRVDAEUr/SbnEJA47mSQ0WZNzHWY5Tae7F7DxMBxcs6zIJlDYw6obNjH99E7HyXeQE8S6
GbH6TR5esMkQsKhv8vB7874t8Ady8GBp8KIcDbBjVIQCZhvLCi/iR4DGEU9RVDZuf3ayfTEosDNE
uQ7ZTnbhiWzncmxyxVezgCzRimgsS1w+zW4DnGAuEOLn68A52tHnJBFHL2l5kaQ7/Wl4dJmwcTIE
hDkFqhkCokDruMcyinHTNVbK7Q8fpTXU5oV70ZqKVtaEyOgyLkL+zJQlnOFnCPvLfzJ589c8bdpC
0zd1TSjHUKT/N1tC3o4xRbQvt7F1GtD/cLESLpa+1PBVhfkXkhAmwoBiWta8G6ntKhSt5QP4medx
e2aoyRA2bqpRWeZcFPEdxUGbj3wr6ypXZ2Lu9w8Il8jMNvXtd60upT8ICTd2PIf9dajYxaiMxbla
br9BWbNUYaS26MzVOLZLIy2mvlsoJ92mjbJSKbWg3DhzJkIMU9AoeBpDWRhwOADupixWVyqPxvcd
WdEFZTewk4pVf9XrATVpH354YBH4WyF1EgFfon4oePpvy3LyMrKMibqYPbDJrh2tS3Ac+5QZ0MeI
mHpcqWRdDW4iyIYrKDIMJLrYv4mkpxsv2gtm5n1cFLUPzJ7RLXv5kAaQ79QsTJ1+pREOzQPJ35vz
5+k/4AAVg4hP4EOFK6nDvDMf0V2537283ctR8sTeKjA3evvTge2WJmY5Tx1NO27aVluhtmhTx9Of
avvuOpTrd4hDnQHJ71IfpIZeclww++mAPLc+a4bLb5anJCgJlvY68OrS8f3BFS6BkTBQ8BaQQo0x
5PLxssh4nU4TJdtHIw3Dld3NTMnTiAKJUdWyyg389zPOs4xiPWcfK5ecoLBJrwVgCu5f1U9btDPz
iOuPdRvr9q2P2K2tZBxXh0DYNxjRY4Vm6fubbI6BN0dxrTPM/2CA7S3yeBI9Lo/c0S3tqzS1Zl0a
2sjaDmX61Tza953WJpQNRz0URGVzcp7rYUD4cYNiHxZy5b/ppoAVUcG1ik2hJQ3Nh7Lt6rhQBoCO
Nvnf8ALVHaEHP5KQZ6ULJNXgnd76sOlWoYLkRWn9l65OhuNK3qxsqA2v1rCayfSSpfnr0aQxLZep
JiQd8uKh+rqHw87RgrXpVfAsXkhPsv9leTWboOqya5HH5dcT+z8GEHnNpxIlU+8/ick0SxYRwtz8
/LV18VhAh0BHogfT7FIMHmEFroAb5UlHK7wjJ8w2HQpOolPCl6cnN0fQmlmRSIBshopHrcZZQNTT
hmzxRW28jotMUZRcq0VlIwWLNoVjXTQIaB1NiF13kZXvWN4wAogsWQ5SjQjTsxFO9jBlv+PPUxJN
GI6pgFXNBbKD1PKmk7NBgJD3JS8FcHmVb43ivIZqpyH8Q2hA5k/RGaBogKu9XcWWcRj9cbjF+HqF
sDnv2BbTtprREwQn9FaYJpT9OHsCRA9TX4KsEIbEkQi7BbaLyAMHLNYd8dM6mZsWL4gs8DHD23kE
faZx5LyHCr/XPL9V/oXrb3LS+umX+6ip5Uvv+htJf2SRJQ30alI4nI4x3Q2quOIutdnSZH0++CPg
+j4WLNaNOc27HgvBOC69Ruj/CLTUwMI2DQep1KQiw8Pvv0jz6zFmUKz3VtozaiTjk8tHWFsrXqCs
xzN4T39hBbdY4TdkxOrjWqKhG+aRl9ubpH0Ahbyd4aLUZA0fnYGa/wc8wKDSlNK68Lx27CqCHsKS
CNj2Raz3qkmed5KAe+cA5LGVP734Z/Tj7rJDIv9ykvhsZsXb3S0KkkfLh9dTfTvW4WlU3MShW77s
t6EDRPQB2aLVdEHAsozsXkcf3P4YVvhaI/elPpvv+KP/bJdaatNpkY12s1KpFXDG552ajKObHJrs
dvQEwpReoAlLq/ppHbKYd4NMjQAzG3UPgysDLc6+cJCHAwF642eRIxhY8348C1wDEoxn7qP+JajZ
RDvr49dxlDBywIO96LJXGKGDya8NJ6EO4WZhxvwzBykasajC1gaqKbfeKEsrFZEFGgA1dUSf+SbW
L8FoCy6N5H6OwhjBVjbTyVmlQHf4am5HvOPNDmn0EY8mynkKqAlqXwHPv1DtkZf7uMYDLx9+drlc
Golp9mPnanc7X4ryddFXbRMLqE21NsDMd3sws2O6NHwsrE2tPs634TvTSck5FilSs33QZzOp2sz9
CnbeG15+8kP3DxKpbqQxiULl6LogUZpNNkMyGa2SlWxrGVpAYDzW7GSIuV7+W/xf1Ds3ejNAWzJO
cWTyzMPvH1sBj2Qo5GmQXv8APxBMdmQnIfg1b9veSE5Rt1wXdEG7wJy364LDA8cjsmFr+DiefXuZ
cnkhZTvMhMQJRtB6PtwZIQdU2fsUhsksEuQBm1SHLC10Vk+YwDwWyEbSxVWy9K2oRY/BScxlvSKw
l0LmY03z17r2IvwqEfQYnWnp+Z4JMQpIdgIT6DNQISX8SDGcAWa4DTuviHVY0Uc4d3kh9dA0ztuH
7D68oZX8bSkLGFIha9N1DmebLKKYwWecQvsv/90Z/zuar3fWBgfN/YS4OcRuGw0CwiQJXC2xoSoC
Uccu4GtdedBvFpqVRiC9vGdQojfRJdRBg8SALQakvjiiXjTFiCfK1TAOz188UDHMWGWYYidBkZTo
C4t+8RN/ccMlRgYfM7BI7PA1tjG1/NUZi+kZKRcy8KP5llZ2mEYGtWVh9/2eWo2sYRT1QGOBN8g8
EOGU3wQylMR5zCVLnUr8++Q4BmTq9sXPqcXydIPYJn7QEYiWIljXLIl/otnkOWPOec9UqLT9Z+6T
s2vR6l6ze2gWyYa7E9Tb38Zng9h7CD1GbOEG+ejf7yXosVHNFMyKmVJCexhj3bbpRo/VEj8WYMKG
TMYjLJDd4Rb9JiNwJfo8gRLbovaJivRCOej59GtuG1j1ycNlJ3oEVSDGVZJIc9mMwmibBXST4CA/
licNGp5usBxgRkSri+yFNi/iqo9Wo+MBGJ40ocDur5Xol3MJEHUCZNkl21CAJ0khGUskwUWqgYPz
Z/WOvmzF6EUHUBEyyNyL5X620tPry+EvvA0x5aklmmTQz24X6W3mezXRXmAfriPvTZRxrZBDVUtW
ADOm45nrzdVXUYmUs+m+1r7GFe7GHhLc8670Ohh2pO5V5YzWpVxfbSQIfPvHAIz1IcRBWi7/bVPL
wnvzNCZEqV4t6KW1Rq3WFkwbbApJe02SdWiVNu7q9zzA6NvOt8JqXV5PX4TM5Nq5O8xDYnzF6Bxe
AtLLH3wHADXZbq9NSHp+rR2S/WxDcnIhLFmJtJZ57LCwLgLaEp2C/Cubaw7HuT3vRp5UikQ5uhQV
dhUDLRT0ND31/VY6TyTRW8/855gXx+oK3ACLvkvdHUQfYpdSxW2C6Kmpo0Mg9ti0OGMsjvOVcclN
w6wBsYonScMUkF7EF8BNcxZrOvMWkaQECYthsDPgMcjtuoWGwJMXHVZyMUj53sadgxFj6RhFo5cU
qCLXkC8Pjdnpw12BGtSdeNysjz1jjd5I3ho2IMwJ4bx0EXpQ9o79rtOyx1oIcQgexPLF9pAYcsW1
MejGIpVJmKEUkKHk6IDryMu6LaGjQi92UoADCQ0HPn5cCC/4YzDvyAzySYxx2TtXwbXpZJlHPC5v
wlHTQbyBRA0cGu466QxIFtHfnoPh+2IPftakZFNmTPgeyYcElbKsK4PsxeNYxFIMVmKl2IPkhoDa
puf7ENvwt7gxtM7142AtOOXN0qf2l70XoJYwNDbexrIzsG5YdxB1bg577qLajlwW1mgdDIcI47Gf
vxAGHmihxqLUedvsVkJghgJ8jB4rBuDqHfkCTivI2iSkZbs3XEUKb43PjLVe2dw1bCYAAM0hwy4h
to3hMjEg3PcvOIYTfUZ/SaNM9O5K82bE1yKlzOGId2i3xViwdqsliB8xp8V/S1uXtoRBev5USZpa
7oFjK53Zv8HUu9BU5eppFyqWfL1wX2faSQ9ZfqRjBZviHSKPL5swcv2+cnTnnMZ75xVQTn31pa/t
QPlsfW4QWlS9bNSCsDPZNxc7IhWh8Cm/A1lV2urFKd8bCHBGjTWzUQfqj+LLCvcrGx92VsT4FV8p
c2nPWp9t2mxZohEccVeywVbe5wDYqMdD++MlQhun9IdYuCyChBXRRLHKmlcl2QdO8cCXRPiHhCFQ
+wPQ7u/GDJ/hKmsn5eW1+meS/8z0Muea9N8JkTU672EG//hE8nMuEfIaMBF3UU9HJm150Urz+wJP
s3d8MjGqR9xc4TLqpY7RVnLXdpTqU70Qa0bEREiaomGTQrTVcVeI9RmLYjGn9VdUAbG4u/KEo7jb
NGnUR2HJBXlwuX4wBiAstmV9c2jDZdjFWTIfBAVJdKoZqUS/DeFBv+VPZ/0NOnXJ4U2vwPXDYxjJ
h4w4E7+WjnduHupT2IsevaOcnGNcPikf1bluU3FxbDTtfiT0Ujf/p2i9wp3mZt3d4vQKSPFc0nEx
TiZY5jgxuWN98j+I0zO4lCgq9/wqJfS85Jqs1G31HCid90698xLLy4KOYPy4uSpuOn4sXOHwDUgV
n7i2x2cy70XlgVs2a+YgRxPpjKvynWXpp2KY/M8eL6Biq6/bK+ZEOpEq6wAR41hvXVpAVEb1F1Wf
e+DwNO6JrdrAOoHZRiLx/+Wl12L5roCssS6vffBxUH6AfcekG5+g1WuJBoHS0DtX1MfKJ8g77mUq
CQCpMWcalnPvamb5Vj5Xq2MaiV0dD8GG8JPbqAjqTW/H0Vribp9jMwbjORPG16ayTVfxEt78+Jr5
tT3OQ4UGcZlxHBd5pXBdlkPkqgXHPNIXzNJHuqaCIgwrsfeZQLU9st0dJmgoHsJwL1rhDcPpLWmf
XUD406r1v50Nt1dmbFzULK47Xhe06tyrY/J+H22ibzwibIm96cZgw2XpnVztrm0e+05y0nSdgJQN
sUMEqJ/04v1wDO3ath5Wc/A+pqHQzE+iWevf9udQcpSL8V8tObSfa0wf6pP1278Ub8D4Lp7dmdEG
YU+YYg5dywPp8ZE97DMIqW6nqbOf8nDEyn2u+qxyriuQ0RrebtC2KQAMAMr1/YO8Qoud4QMG/R2W
CdC/uHSDuHWRDE1HJDxyTYR4e0Or5Yq6io0v4TwIluiZH7epKhSu5ASFwU1hSs5ti75N+pwrvNpG
4biDrenZeChzDJDbMs6HD2aAA4+LZvSbCmcMoyfXvTVr3F7GvUxv2MToK5NyeHhP5zqMgwHqmwHa
5z0h3MiOI7Bfa9uYunTac16tTpTFLsncMLey/4AsVNu3/DA81lxPclnJSYQoz483B+lWct7Nkwc1
0WPQYRRlJ//ZcSUZg/wQJ2PwkdIyiEEmDCXZUtKUa7Ts8lAgCVWSTnLXzl+UYhFEXBX3AHFQPNgQ
+ia4oWXaQE0wPDFCofWDcwslx94Xvg8td4jDg6loBwo9wiHbSJ0zPBPRm7YDeA7ITI9KAOvT7NFf
Qg/cDmb2Qqc5SI8NyLTONDgFFdKBzd+an5MDxCxnF4/6xbvgaAfrUdxTYWp2JJcZ+Fl16mlqkvHq
usa5nVrC7zVYnCJTGLEhJrdi679N/z/he3Gm2ZYVm2nm2VkePbCxZLCPo0xXIeowmNr4oml02uGc
4V9HVY+tBSA9+5GVYSeoESXYf3lOFqOnrLSedIgDtG4W5+KTWot6GyWyelNOF7wAIxUmq4AEodWu
fxZn7ntQzHG2/sx2mlwDJy4BRjE/QwiErLPhmJeycFwbyp2EeSBmQ4yy8cmY6yUna1yOOU8faruS
PG56eVopuPh2UatvwyKN51O9M/ydJj34nr8X4K1ja72qro/z/1F6VvMCmFLoqRXeWk2JPenf0fLl
aiilV4xzZPU0v00+9sXUZ4M63uXSn4gc8K0X5fpcUpbLkVUVi672hZx9mw0oi2zhjtwzoYIzyjQY
TE+XvFibuogDX/Q16F07yxQPVJxFeyaVWUAyeec2Sr1bnfBBQ89LG/K76WEf7mITQWcxJ7dRyufn
w1Md2T18awEL+NFNH1ZszW5lNW8bxi1GwPzaC+4aZMxd95UcoqT/8DmwMeF9pzbsAfbEx1EossR6
i7n+BGCaalWjgbmYC2ZzaX3Jx1BbeGHK3AF9mCnXeL+YNZcygnLZ6rrO21Q0141AIlgggKHrNdV9
oSSw9boHErkI0jTKex/gsGs3R4uhofVcC14XXeYIHmZrtxy1pxOJYOP5FxPyY3eUa5QiJJc8ORwN
5s6C+jJtDDUkC12V512lcpqA5COADrtzB86rbhv/JTPXaX/w9q6hKu/4IszeinnV/33cdhZFQPdm
MQQMOWb/WfmvWHe8HbT4jRk5yMuxLCgtLDE+2qp63iwKoyIgksAg09Kp4KZ4S1njw3jzr3BEKSgo
o5G/zu5xM8qi9LqSV00wnOpzOXvhqHiQuWAsvSmlj6Tk4jzDy3Mmk0i0cfdGMhzQxHDuwNvr20xE
EiGLQh+EHxvafL0U6Zp3cm0NpF+mJIFwcGzAJ1iaTF7sauxSuquPcoRnDWABXMAB+oVIf0np7i8u
rHfKrvQfYI1LZSitgGz86uEJAnHwY6CT1Mfvay+ndXPpLQVdKn8QusaFZkKYMNrOvT8P8+ybM2qv
vWLgr4bPEbMBb9ilbV6kmZvndqiGmCAibGP9XNARth2jqSgrhfrz/RHKFE6KC28Al1zb66S/y4dd
FgMomGj5Fc4xSGwEFaE54hzn0se1oG6aXJ102VVIhLDEeuV/nFvT7tfnyTeKwHSe3Ckh6jbmt4Vr
Hus4ECfk4Hgj76qkTG5zY/uK01psu8cj+Pkvf9LIlYUAJ0PD0PRiqYnUyk0u3SPvMp3KI9X5eGvy
xDwy7BAjkhroMrTT8zlBHPlX0H2oK9hr6gkV1kxBiTo3qg1DBmDJjcsJhjWZnVSpA2awnDCDbpMf
P2nzcZsXuzmws5JM6tHryKP3vlP6p9KPBfZQ1zg4yJuwUJm1wihEzVROZKBJRtAQnOLhQpEPPoVP
Q4tBxGR9F909VH1aGGONyY2x1BEnDnxSv9WUnWNb0QDTw+8n7AsRNbQNgoLycadSJsO7m8V3tuVK
oyUUSSbkap+fRvWZTXzJ/Uc9wkrOgoo3PbBa+RYzaKxQaa60UQEc/x8U7Wj+4VQ4WqhglisWpNAl
scXBeH1qAjQD5tJ2e4d0XsVIRAeaPHI2AERvZq/J3gSt4Tc/2qr/Nw6Vue0/6/43AD6WGMiHlabe
+2i5xAEWfo/mQlQ6+HKTSKk597fkUdnzXMo4VU4lms4FR166wjBy04Oq0zviKXv7BnUY5sXEzGzd
Nnl5fha+6A6ZOPJ4EAN9+RboeRsUaYw6jVJFkJ+kSqkWBPsTNDvD2hLQu0n4uqk2GfqIzVi36hSI
nOC3xpGJHyJc/aujV1BpGCY12imt+ol2VHoU2ucV/YPh7EPWTuXTxG3zDdJGgVt9anR2WZlMGXvU
f5IfQC+2+L/68+efbsUGnWT5Yr9k6c+EUJNYi9OSqEoRcK+sAqEjD50fcestMlt9KBsrbMQKnlV8
wCUBjpEH3OZ1+fcg5v2Pbc2bC7AGipCzo0uuGNBN5fvS01jjBgkAWPwvcD+cZTyVzvlWI7VlWdin
ACdVeJPmbUvJniScYQCgSxcxrDWbv59wdkaj+e7HkfMaH5NtddqrffbeaKAmVJIGMvHzDRYkqvOM
yXKTMq5yv7uGmkC5fCu/4reoe8IOEgeYZaYsWaM0aJzRe1Mv4U/pgulsS6Oqj3mrEDioETwZZ7wS
24oQj2/l8AK3U2qrfO/JA3vRO8opJ4RYYt1/jW4rehhsVFZmrEigh1bYWhbwQ0opIC6d7iFaa9PC
142k5pekOip1TpH+HioFseyKET6pk0A+tbKubyhbZlB8y6ogtPlVdJWk3C/uJGD273+spNLM0HxA
PzMFbiHpF382xuAcnj6X46gMj5WTanAxFoejNnuG0ZKfVqLB82Tq3NYN0DOI84wLFyxCaFQsQ8qS
rksP7Bzli4N/1AVMHiaTjfCC5sN+wd/rL8H7RfAshvkzGWT3mZ1Y+JEsolOJ3V0JL9WaDkmnm8GS
jtuybU6g4A/yYTpo0uajocAJkq5+0AT9aOZ5CVGYYgi0kOwcoJNdGfuLjr76jkFjdgsum4xy7o9w
hqsxD51lEVBtAJmD275j1hs+PD58UO8tQjIiKvWPZM0tEjUejH/Yg1jOPz5PMhq5hkFW1DCM6EDk
xUtsH1ei2GgDLHY6o0qfhLHstvJCrzIjKE+GwYn0eUTVv07NgKDI2S7xSx5Ep18T+WIjVPcfcKwE
9at0csxRbhjF2lN23qqCPkQhI2y1+Vgajw7H1ZgRhvsUvEYPbHqd2FkUaMTQacIxvVtGFA7W144o
GQpjZevk4vDW5o2G8FC/XP6MG5IdsJgLlwZ2Sbip5NWPEJzu5cB3W8cn+YTpERTdoKWK1Tw/2sAL
B80iBDHcxtnsHdDnft/tVXf4nPUn6FFxmKXSQCGvWRtZ7R8WeM43LkCjQvzBngo8DJz/i7nYReow
M+Gb/K2O6eRYfLbmoy/yaJFrvbO4wwxPzCswWuaCQ/WSY5hx4NFtvj5bfk6BhvksUx+FTNdJYVdX
V9r6Au9/owV8xEJDDiZ5HZJ9Yf6KmwDcYDgLyGlt4ZifhBouBZK8dID4z+6xiyChZhr8kPtuXD1/
D8/4TkLYawafoQMwtKdspCQ9ekTYz+42UcvPXJk0YYpMwEcXT14mb0xKq76Z6EpMh0Jzoauxtofm
6fcH3goQrv/RXrL3fIzBniYxiYrOGnyECU3PTnMI7cMuzaftE5uOSMc49GKrEbuf5NpCaotcJwck
ZCt95Q2KbNZ0x7qyD0SFJ8757ithVu7vjQ1dRCuOLInc5kRpY4PFhhhGmZufjE2ThZY2d1ACdfhy
nQMk9ZgNxkBWFnm9IshZjWwV0qTZpeKpa7FlFf3UFRoR39S+TFYDStyBIiBN3vs9fHsET/9kTbNd
ARjPI2PLtyuu6C63Q/ihRnXpWacMZEKsVQf+C6Cdta0+2GYppMCtBSiRTCkYAgkKWRdx2Xi0wyOi
r5GwcQOurV3a/JuvJIB7BZF82CqeIaCJBvX0V0QfPRxpHLKMmCbJHvRf56CNSHP7C5DxEBm+9SIt
irEqGGMhjziBMwWAnocvu5NnXo5V2gN1XUbt8I7z7AqCIoPaJTEAs+Crkl2Z26hX0Pd85Y0270d8
S1MoM78X336ciYkX2gdpttLcdmgo7oCfKzlIIhFFMnod+xMMQ7jkSiroxFi5TI+g18TfIQtkJ6ke
XmbjPL3Abk72TIMir/ZEwSFz03zBU3vpiuluQO9CMtsyXOvaEXioCNqJaGzAayFULQ3nTYw2rndd
13rkr+EgEXduIgRqwqVM490jYz5iPa18JThX8XaTxirTiWJfDrSxfsI42ekCSEUpFN5oUkh0axCw
nukAfpn0dXSnO8Zv3lp8kS3x4CTs6cYIb3nNsP5z8zHqazU7sIwtR2A1mMoa6SczS3JBMHONpezu
BOqQ8SpHtSB9Wespk8Pgu26XeYSsq9RIZerrdE4Q/7M1SgxwJjzLHs0sw37PyuYgjukAgzAQ387J
ZkGZXTxjqC7CnrGv8SxCMGXRM2rCBpkCLs6+Bsg6i34yjlCqPIapZ0bDHfRuKGNmpocheHosV7fG
UGVZT1EycJsLKSpAf9v9h1Krrnzz3XUS8ebgXmtORXgxCCEhE3xp+a29m46l4CW6EBWPZRSeEXye
9VhUuwL/lY0boiFf7O9T9Q+hYID7WGycdVuHBYQrRfgNxfikTnob8Bsdgutf9G9ujRn5vKC+0IFw
+pjfnJGGLxtWMzezKiuLIO92Ts3syQPViHi/QYtoUwuNw9kYEZbuJzXE0U0Z2EatX/mxlFK5GqiU
C1sfEkFyODZEk0jXZ7n3xRXHTUEq5Ano3ZIkpkfyJSQMkios1nz8Xsbu9FeHCgr9jeyUw7RVApG0
ApVkmcoFHmB8NrDjit6sncpiUpYbWzs734Qop81w77sznV+jvz0x0vLHTBdOerqH8Fys/uW9dhsh
ReyfdYASwcNpkHdcP2S+5pgESDsEdrwvHhafGeQ1QDVVwGVyztU3GlmU3qpGs/kgzgq6S7VWwb0P
ZmH2Hmmg5LcMeF5/0uaiUF5fEGqjzRiahngQm0gy7IEHrQUHH8cRDYFQQYOFKm+5hOLD22OEA7yr
vyVTUaL1yMUP+WXPgDVGuhOThU5tkYeuurhT7UIlZtav61VBJbp1l3/YvxYt8EHCoweNBrTDL+sU
c2g1vWff3rVTojljn6iGfZptQDRqUy9jMbeV4dYNLOr4MGPf0GRoX2hnwSLzdKYlT+RfEUJlyVGL
x7YRCnAxfg1r4bbdiUbLPTWUF7+kOifTKec2zzPc7iKAqTj7vBGfV3s3nPrS1HXgzRTGTFIAV9ax
6JDC2O2yhyt2Bbd8bWfQLJDM3ZFiAzPuuYGPv2xPPmmebpDTU+hLEqZQSMnTOVQPD3PvftbyuK4w
F0jFrka3MIEV+LpKt273dy8OZouJBgMt/oNO6FL3d6CJLrHZCpSQ+ajmbiYMNsT83vxmBNt1JVrH
yNeVcfaikd31czI7OB0e3We93KadleSDsdQ4k/WTWNckQlwNcx1w2IlQUvgoDltZ84EUsAjfPxdS
hwlKimv9/VpG0YPRJ1gJHEA3bJqQhFtvsCjLbWO5Z1jQNTCmz5Yo0i3V7B3iLjYZ2/7U61GsXUF4
7AYjONzJA2gD7Zcbj3HtBV/w9nBDP5cqUiuR6GiFSnD6CPtDtGzJB/8QVfa8xswBPaU/HQYmCkFu
Zcs/W7KvPfR8sqAzJ6fFDPhMiG2BVI9qGlkIqGqVimD6jY/FFJRwa+3lUaNBn2vNAKN/o6X/ksBs
ULqR6x+qOKApqlhOMEDItv2N2GMv9QsLQ7ANpToN6IY1BlIKCjPVhPcYtdOf7Pel/ec3QtpuY5+x
1ko6G0RaLWLQUZxr8DkxgIcQXJ3nLJAluRyOhO3se69HZD/WvshLdGM3uvyjL4kCXnHsjGZE7yYF
/TYt9t9E2X7i31kAjar0M9vIFVFRLSf519x7U6ldZL1Pov/wd0+lDNp7QSX4z43mhfW7Hw0QbWH7
UA3c7HX4GJpd2yJkvfdP0gc+ytDioghrPuxNdwLW0PkJwTG8cYPpCQmFC5piYqwqTU6GbICprdgY
I4pim4CCoxWF53vkXe63pl2+92GlOdP97iHCJEkIBGd3RyTABue1kUfhTR88trP4sYBRW6QBTmJj
jEcjuSYO7Vldy0pc45z7Ff2DA6Lqt0rvxBRLpVPLISNlgjUm7NBu+kOxTLKyhGcV8Qase+j60Ec9
6aEYVUupiTMOSGD3dWC4UNvqMk+MMsJ31Jw+upqIf5RgfXO820OVdPIvZtOolStrLTdPzTbfWmj6
/ZMR1UMN6EGVs+bXtbI+9G+aHpKR1STDdlBNgQOQ92ORswjhuS37By0D42VuU6ITfy0YST0vzzIc
5zxT1C9Ciz4f/3uCKcGMjbdktw4lJic94ZPQFOJp8S4ped282+Mnwv/Sx756E3K2IRtdAB10A6vf
Ic6wAd12CjICakCio3k7WREwMy2PMuy1IGyvUfKo0i6mlAXZlzoM256sWSnyrMn/tOxo956RPkvV
a0ib3s12nqEDob1wupU0vgsE6DREKlSXOV1JaYTeiAiOAWD//fOC+yTmuVpXbh7zzLAmrQKrKx9E
cynG4KbI/CvU7071PX3flGeWxkVAGT7CSBLxCQy/y8+ckJykYwuj7LrNdL6ccMSg7vuP4/1Lrbm2
wYVJI5MSNfCcLUV2voVtqeiQ0BV7xO1/W7WCeb4LSY0VrLs8dTWzABrbZSGqvimwbtuAhtyOj6+Z
HCflYKOAuzOitYdTYrCI6nJxKGXoHiBlgmlh6Bj/E1NuAn0T+mp3UuV7Ola8IxFZkvmodZ79hCaz
GEOkZijMj38JgUx7HvfEOxrU2nCU/lu4qDabsRvLz+xWy6CTCnpo8p1Er22UfseDNkAr/sJuYqIB
vE4lJ0RCUrm1mqW75zVa9UtI9kFxhfw/Ddfju/wrnKpozqm3ptfW4KRR8q5vXbulhWaLvZ7Le+Tj
sIYfVnfGinTH5NTAICAkeO8SnEK88tlo4Hjf8bJMFEeGV59G9Q7qKzNZfu3b0lxH+PbzkA90bMyy
Ck0sioRS9wvjrKMypNJLTykIqwzwwYOfmia0biRhpSdTndBZokfElAQWdnYtIRAVdOKss8x5i0Od
hWggwR5WedSxSVAEXBjfnIjdeD9wFB1X1L9y5j8zJpc/otiaBEl+A1rK3dNfwnMZAC+qXof4vAq8
Frr2Vud+ghGmkFdbnoFtAtdzlJKeuqRYuVPwoiv12qDA0TGeIcjpRR1THoUHnn3TQFG12bnIUQm0
kFfNRQmz6QBFfGW17W+LemODUS6FYrKH2iLc8oFNvOS7ekJOoT82NCYSGEhkPMO/KZuXOJSlN9ei
3tdWZfLR9pcN4l9df87lxSgMKRyvU2XNaZ1LbL54Q2iOYXvgaeGwVzDyi8MZg08P0xzHKbSuKRoo
mCnRAgnXsED43tfxA2dX506eUqGay24m8JB+sOzX9Dy9YPlt9paflxvVyfERs5gndt699rUZFbVA
8JoDG+li5vHtplvEpJr2H/0nYT0QADurGUjXRAd6kIS08mUWrxCXhlGPvKf02SNpEONE81r58E0e
V7hZQaWjb/uSVUN7hqUS9R9OsIoOBlWPZXVLvp0vjCBrJaiBFxijeFo+RTTekRivMMAoXD/W1vKu
NkEyEa90+wcZbuyrSSvRawUw6F7zE+8dvJGajmmuWu8/qySz/LfBYcHDXoa+D6smJmMrEck0BEO0
A3OgonDfunt7C+b+EDzKQZLJo9kGNY/1qS7PBP4xQ5bGTh7jKpTJ+1JkpWuxMHzaBNxWbG8ro2J4
QBuA1mNnTvJhG8bDMah/5ZhW0X/gT4RG8FllHSPK1yKdk7uRvl9o6k8VOZhpRxW/v+5Dg59Bv6RZ
anb2WjFSCF2PJyZ2IEuUwi4UOdnBYr5Y8uSeTJCUdmFbikGWadUOcttjE1jbpdWZeBfMUDpkL2ue
yLHmRq2ztDIWwxfUq7LJNBuzjwE+3oJpARrfMnc8N7k+cuYmFw54KGSxOkiUzXccQFG5SM0KJaz2
n38e5YhlWum+MBvYvBx5gNV9K6iVdQbSHsSSRjG/WYiXMRW1JAd8CfbKaXAASz0FZRym2YRTXFj/
oGNvwn+yzgdWHj60jD814bCqYBdmn6bVtM5ib0pVBAos9MqUNNk+yhHUR1KeB3zsrit5gUha+R6T
1GnJaI1wPbyPgJ/x72TXsG7e/8IDMGmGzmgBTXVjJTwSG5sG1MSgR2bvo+YStVg5+v41Aw7RgZ1Q
rL07ANJrokMRazjPWkdoRHKM3hznxJRiMuHKrLd829vnlVwSmz44zr5CcapP9m8tOT/K2Q9ejXeh
L8edDEtbzzSv4UnZd2J2A6oqFDDKWfkpl56wTHNDMGnhaNVmKsKH/2jTrhKoENY275HcJJ4QQRiv
rXyn9bP042Oj+DtcxC97cKKIDEQHUrborVxIPk1zzxoybrM/X3IFeenK0ShYBaFDkz3OAfMhXcE2
be7H7gbZALo838qp1rynILQZ42vv8Wew+psMGSQIygUrB++Ea7bTHRKbXyAq2KfWl+aalL4GbTPV
birIc/JQ9EGtMuACUj6vNiQAqvNs2psGdHofAmcAldAUW2mDEDkZVG2EhiH3XxCFaCv9tXhw37rS
voJfZShFKOewocUZ8ajkuzJESgcKb+EmqqtNc7YbXNdxh4p0FkEP0q/rXAZasNPuENo7IQuvuFpz
27JvRitx7p0to/RBX0NpEAJccF5hyGh4vTyD7wd8vM0X8f/zfoloIs7vSkN+pYl8E4glel3TqfE8
/U2Wd60vomNAZwqSguE8x8g56w7pzFouT3V2e1p4qTA28ga5EYiaF4q+qIlTtCn3Q0MIVeFTBB8D
T3PZj4a48pEnrgWoGYdSuOlyKjR9f5wWK7tWcvU6aypVl1rQDGwLp7q0HaOBbrxo5jMrjuY++xog
ozx30b/SPi79tFLrjg8bfiS8w9E1RSpRKiwZTZh0xRNctGTABIX1kPM3Z1UO5+aco/ytvspSXhuJ
noMlfdYqaRDPlFZJTWqsMiaNrMYdg1CCBdu/EODHJeVvKuRmj/JHCjuc0XabBzhI6YasN1QmTTGL
zMq1E06vSuzAieOP3p6gpxwqVj9Y9XmjSVwkdcPKYazPub8imvQnUmYhRGccPayy10DdIpzp3cO5
1+iaicpeb3sVMNUVthVqPKnIfTTA0lexerdqbrxS10fD7yBPM0XshnJw03W+SqeiCLb5GDl1nBOa
mmq+qFv1WjFCPbLbyiQfvcorF0Phf0zF0D/aswiV0jYAsaTMxEbFsD5NoMCXI7LVtyKJP2ay5Ipw
R4pPOu4opyMlEE5kOETcnO1yh9Do4yH4cXAHD2OVmprVZBnB29UIOzKk46VW16kLYcDWZC43ocXn
x4TbOzTxdE6X9DTBhSU150PjYRNTNkp04hdATxSzo4oAniJNtX9K2bpZmocvMuGyVfCkd4zVYCiz
zGPewDvYY9rXMi2pWHYHxUvlUL5yQN9+HwLSMpy4Xr391Zbiev6Sax+aOYYZxGYap1mGSsPHGtHi
5G8mOVLpreYV+PNAqqSYO5dUj36eWRDfVsM9gRmWZlkKbg2w/SYnSZ5zTdEN5fMCE0/M8h2dfZZd
fJQE6yNEpOsmZ9HqYBYabQ3qr79GmyvsiJrV68ULI8IoMEe3wWNkV8Qw8qd6Dq06rV38TGFrHc8H
gayEpXu70DVCHFuixha2MZNrZt2XdXb7/KokXqBzoKViNSUUhYJ74iqMyrIHfDgcVTX4JMMO9uaF
c4BDhxU0ZtH1crk8vpaeJFIWVpjQYjbRTIUeD3h7wWnNPH0mq9mxsAFeGOUMXnXfdJcvTcaGIDaE
cQ56eWbdMW21O4bZfte+gW/mr7md+kIUPDXtVzn5sCXbWgsIKBgMCcTqrm5dFxOzNNjmeGgWx6BE
IsBmv40lgnXcFCca65fe0OFx7EKnmOSXg606a+zC5CPlPzrfjg2FR9gYCvK7NtD1B/MgesqWo/gP
lg/GAc4NKka8n56Oy9ywC6I5EPHDCmV48W/4gJw81DUaF2mh7Vb/Ea2ylVAR+nvqfIC9Y5afYI3H
6S7TMBrr8GGjRdVeymW2KR0tXDHS1pWYA+gs4KnCuFfpEiq8NyL1ReRG+O9Yoz1uEeg9JJ8JGkmy
/ZOmzs4NWW0a2Yy09URO4x1AdUMwedhIEVbq/I9RqYvO3UB6uNHz376WhovAUQyfmVs3W1pA2lBu
Ji19kPPNdee05jR4endSQVJuVzDQ/rg7am2IwfqjKrelWdYDvo3VVLKpskVp+GBSGEaldNgg3ON7
3AlljDQi6IbwkMAVYMkyRWUri/MjsA8rG/LasuvkYEUosinpc08+60BXNG6oROhkICCKFy8ToQIJ
NFVCsYo1TtTBpogasIHLHMhyGANd3INbGctglxFhCzPx8ljsKDvqqkbWu4TT0l2AjtOwuJIwNkod
4n47HLCIiQOtC9t+EFGineFDjU8aNR1yChSP5RO8ysNV0VioWJEcBHDNImAJp1eFsiy0L1G19IaK
OrkmyVcPCvGWWStaauJlaXUd/foxesGDIWKnYymX2dyF2FCMEQls39oKSTYlHQwLBcu+ksvZuRp8
r1PeJQg4cbQ2syjIKq55ZKl7YIlRdPRYLY0iqXMZR2+5VdQ1Z0xl3AbvcEe+sGsy133suaLeJJo0
LiZhaPOgGfsAVcLHPI9lCWdHsQTsXhp2LcsvCeQfuwwv8A6S6kryOHF3ItFlD52aEe+9WCabNWIJ
4DlB49WX2hmB8+FYCUPWXzpf76ma64VL2KtENCyP2m4CFFPEJEVqpgOmkv8vT2VPUSBS1dp/U1eB
KmOk2K3ZzrZVVOOYpuRi7QHeKbFy/FSmNUeLmO8umWZoDSb/5cToVz7hED/sb6/opAIkPY3N/vDq
vksY5OR60QlcyQVNbC9GPBG1QGpSJoxRpfE3GzhTZHpNHDomk9yqvg8Lab7+WtZsXi3RBC6cqqIC
9yI+PEEXt4NJdNvrxzlxKW1HSc3un7tmWJzKJMOalMtrL37zRT79AXvvOr93jrModqbMcbAaNZJa
HEtwUu5xneat7ER0/AuKTgT9uNCRpEqRuf4qOoS8X3Sh0accZWGG1C4trsr5ZxudIYKzIPgIdiVj
DuFAwVmfRS3FWRSlwRRPaZH8tstSUW4jgfLCTsc4AAmso9M/okg0+YcaCLtnM8yJiRzekFwz2UIu
WG1mgKPQjU7fdrNTZ8F4/Jh5NxseEGhD3JKEhlDRPP1SSKaVRSywG2hMNBbS/F6+SXXZdNR9ZvYj
hn6WfXaQxYYgC8iFq1izcQbYqYgPB+U0zpP9ObPYEtGUUQlso2HdJmCbyTqf6O/DrdRkuZXMLlYM
2hKGKm34TsNZM6lO5TFmd+jEc2+db/0D/14grLZ70oFnMGrfEGJbh2HBrNaNXMKTwDahrzo5QrPw
mNpy+RE05guS4fD2v4Rq52nTOBr3GUa+szPiE7E9Udfy0oanN1NeMZHzoJg175F7qxPNzSGKc+eW
yweFASa9OGssUKBR8qMXkKR9YCfX0CWW5f3n14QjHPwYx7ppeBuRHow3H2X7S611Rc4JVb2C78nM
mVbdu3ixjNKWX5UGU+h3L1DQSoAqcsNs0g5fBxiOiafmRXpquoMl8C3mganpEtzRk4xKGgErJ4Xk
iiNWvMqfdUDFbqH8vDtEt2BAa6hzmDfCFTICUVShNkZoKSVlB7PRwqILTK829YzB2yMxcCFijxSM
S3TMJNWye49yrPQJSq0q2M9cCBqzK4xcXiepthziOmJ2cDGkrG5u8HpYDTQtrt1KjXTj+L9OPtnN
QIz7KKEVlEkC/KJzg8jP4jga52myHqPBoFg3YDdS/KWFcGSpdr/B6AD3d8404Spw7gJK5uaq205y
LSQf+XAeUIYHU4rM4eNCLBp/g/GAHcvMpnUXaZVpcrGwLuwhBSGr2JO59C3hNrEeG4NIrCjJcvVg
5XBkdqiM9oYju8XKmHGMeSJbDQDqG8Ei8dZ2A5Kjd3I2noYUnJaM9HBwyVDQE2a2hOBI3vhum3mN
8TPwcys3ueaGq4O8UsYodesTR/izLUV7HomBSLzGpDQhLs6yckHuUtA/TRtTzxHrqTFyInIANMWt
GoA/6KhQ67C/DeOj/mJrTyXcIT75gh1uk5TsUx0PFUCFkmO4/fvNDhavCp8JPvMbjD7u5mfiQc29
oX4oC5VlL8FbKNVL0TCx+tw/7lLMrGHmVGGVmHOtjjfE6RL8Xruokzd6dsBIkwYNqeGNN1XWgO6/
HSu6LQzSS9CXUw9HvC3jcNZavp8+iRsUFxDwIHsCWSYrZZiy7UWV1SFmPENCpAT04wAXxFxLyakS
liNjFSWPv3lBd9FHhVbJQfgkVN1qQ2ZVdy0LyG3+af6OC4LNKVdGWL3kSR+Dt6icTmQ5ZGEhdCgL
IQl2ICAnXuVY841zJHtxvtzD3/YO7HaJiJcEHkQojnoXq/k7gH0Qiz+yeDMfgUKopjQhFdpMNeED
84m/2re6MRhQv8etmHRhVOxZMFD8OoB8/zq9J4SI3WFI8jJVcUJfLZNvgHh1z/VJARYaQ2tbelG8
9kmN7zwJzBa9MxmrSTfm7dWkRfSAobisF+nwN7prXi+NhVYzvw9sbn41fTYsuObDsCZxk0thd5Gj
x3gkfQN1dGuNi24BBBo+WiSnZyzALYMaJZpN2aVXlnj9TdYpuOBDEGVi9uhbJCgltYLeAZAdZ/qr
TpwdJOS/0WAfDNvvD7rqEMLSOSUiDUzQTNEeDmGi2LENYI1sJJA0scyCoaXZbnN6tqcNkIxE73P0
kjHIVv+nYkQNke30wWpYzaahow5Zdgh+2TUH81y1QMLHnCandp7S6/i1XxydRHxYAOl7xY5Yi6oa
aJfd3cVBkmI0czZ3QwfgWFUXV9+6oStk/hGte6Wx3ENoab2MqiQqoX04bB8exBDoyHhsNoAjy8Jn
rvjnIzgUKdvyqNRQi1GLcEBizz19mZIzp4eMqFh4DLI5jIGt003jM+h8HFgICVqkNrnDZiT49t2H
TC4NHvnbA2OV0yP8VNj6JOovxlxLfH+ZFOVhPHT4yodjQZG1t+jWSdpTW6B58jLNg554A410t+kv
qglefYwCTna5a9AkeQesUwG8QS/olVau+/GkQyeV8YLwsSoMEz5JI3c2NNhDn1UHXP2L0bJQYYAN
Qn9zwBBg0+sqAEfDlzIvMX1rM1O3dZPOOdCRWDxLvH5wWD984rvF/Tvb9LYsEjcX476BrgrMp+FN
qen9OoV0yR7PB5obObrHMpdcDzxUrMZ5Y6nRlqw68fB1/y1dtY3YyVLgiPVY98rXSYD4mX2kgC/H
0JxhjYlekqonI0LA81EUUmrdDBNJ8SidSnC7OFa3MmIjNr1NZ7regu1efNSK3vhJumUG4+6fOOgK
IcsD2/TGuWUk0VRTIzLToRIwRbR0mDU2CGmd54BkgayCcMkuYuXU5inUZmXeh9RF4SJGhfbT8zkv
XD3ZXVS5H7XtSBRRQjiOHgzvdK6Lw819Ye9JCiiHVE4VCkQbNzKnS2OSSWpmSFK5kCMJ5bfX7L7C
ms6A5NmfnDHVduaac7CepZEzpdRyCexRJre2/7VEEH/b0e9A6EiW7WGDFyBxKGQdomGx/x8q5eec
G83BBpehpMOjcqqbixkBHwuvsgU5wvAao/PtMryIXLOQMKYY7uG9zuyaja/Ix1QQ876QBr4Rme9A
2FqyYcRBi5qbneLWvwv06LF4VjlwOvfX2QJ6PowqKqg8sJGe7BS2dwhfI8MKgJyS4TWnpbrC++i6
qEZMKmzzCoVtSTYLD8FZbZlFtyEppDG+laASdz/Q7E/You/gg1qDZCf1UoAiYmnfPa+AAfWrybme
8L0mnhBSpsZ2OGrJJAPZkCwyEpDNSYarRXE+zuepVo24wh+hAqg/WZ7tkTw1peg1ITW1OrWZKOs5
bxq/1eZO5EM5/11gYAobCc/3YEhSicsNYVocr9gAlVV2mEHTtd6hoqHJqBT+hLwQ7pu9xxto11/s
pZ+pt61TMMYRhhc32agJ59Rl0nl2K748uS6rVzQXEtA6K1m5QqctXMmoFK/j842EgOXr+jSE84MY
XTuQ6WXS4zlXHvP/50qTfSLlod9DQ5kFW2uLANqxRPXfpyutL6cwaIsuFsATYNZ13DHOrVxB4pLp
EeRTnWFLv3/pbBSsrhcRC70IOyC7588HANX5RZ2w58IauvZuPRJoQhee3GZ+ZepspPFWqS5Yls3Q
XGASxWdh13UsWXF28kiSO72oFflM92AAK/c+MTqNDxqoaqO2Gxg+dFGMX1AQkBjXFfKvliH3FrJg
6mzzNHjUoRIKE2XRRLWLk6q4J60EIoC9tCDQA2Lq5XQQa9CMT1nbdoD/xi5yEs9anJbP++koLQ6J
InDtDmGgT0hCkzH4oeNG4FOmScGMX8rXHZKB3rithHVJb+um9GSaHMQ7TvEuJDzvxe27E+zxRZzf
u8BlwpvBvFg/HERCHJALJw9rERPNwOBVXewbz7wBolj+MZzHjnbfCZw+VFPjcHzSVAt8DPEZn2UU
mO8Y8K/29oNymCbkVcCWxyBR/Ow1WMvZNmO0Y+MakAoZC+U7R28aido9+jb4xKVzKoYQl1nWbhdV
ESYAwFA8wbqSqzU/fYUYODyXR0OakUrTdxU8tkfF4z/Chzp7n5sc9XkMO5OxbgDHDnK/0w8PUnXw
yvaH11Zs15NkTGYd09Q9ZtgmQFmfgPsjaJJzl79HweP6Pa5cP65dAJkyx9MMOK7w2iVB0q9EyJds
iE7RnuMOxaX/39N/dFWccqRnIFZ17h+BT0EplGP7s2BUMuDHWTdI0wHFbiAnv2Lxc8ZezwjFb9PO
IAi2xsyzXX+HWmfs5+iqOYL6mviakLtZuhtqo5wxv6CZBldvp2A7WDm8Y1UGA8hlFkE+PgfsP5IJ
nDuGi+WOGkmTYKg10nQnKjeV87HIQAlZeZZpwgZg6Jk0dhlzSPwQ5eNs++jmWDmbb3od9PS68e/h
pQNU4iUP6NA8mnXhJO6NHi9XpkLa4AsicadUqrEVHSVfPeG+LqBWl39O/TEwbKPa+FxZnNgT9gmC
S+T1kZnbZopYYtexh7J9c8+6R/TaBD0JBDJYDmqjhOLtnABULioE8HkCIAU1wR3zFb+xDLQ02mNP
+1ZBScvSmwSqwrowZTeiczv0JmZ4b7zP81Jz8fH6XrzC5MraW2BZfVLvUA4OxSYINuPU4uD33SfH
TB/n2sxq2ajdhV6ToXP63owJa24OovvEFzw64F4xcaiW8SIlaZtEWFyI0n9MMtWxDMBKfSILgYHx
iw1BVhBIXQ0dr3gqduBIuavkjS3sxQLfeynmdXAC626DQx57HOJM8ce7GArJ/J8L50trgjx4j3WL
COFyYQywGafC7NOHl9tt1RBsrGjRz8XlbbV0A5+j3385zRv6B7BjWuGsPzTxXb9WstWAMHUlXjBT
g6493WrPgGoDOUFxPR1XifRbzZ2ixfDBUZYbxBdEEJrNAbum7T4dHwbz4a3PO5H9O1Q6sIaRCUri
Cqd9WXgntd93mWX25DcV9Q03N3wIKmVUJHTh1nBHB3iLIysZ+bd3siH0hYW1ZOIt5/fqHz0USSlW
VyVbvIKKCyG8b1R4sJOl1Lr9N0qroS7ZTXxYNfXMm9Z1aDu2mcQwsX1Oaq1bAtXNDcIKFp640ZRQ
yNk5TMq/x1SPubyFkC9YjKBZQA94Qj0z0afX8laJid993u1NFohuGIF3HrEC1itIuM91rKO/62Z0
CfWnyXI6hI290bCdMrbGYI2kSrs4mXM5B//Q8TQYi9abyij4Y9w4kAQTYxztBAdX/O9p9FkJ3kSe
6T0oiF5Z3/DcuyDh+VuKWM+edntcbMlG2Fb522fh/gzUGYNJVzmeRVpLey0Dt0Y5E64WhQMgbqlq
L84DGKbPyzQz6sf6vIlOskOvOms4Ry+QSnQ8VpvopoJG0Ww8sDVE1hDPQaClPeMPVDhBK6/Fdkdb
iyyLlsIjcgySvKYgfsybiZABeCv+MQ3MuQTqg4H3LgL67naUtwVYDNXYB6DTc3zNo2o5/C7X/x7T
Ps3U176ywrTJRCRfW/AcVORokvMaQ6lVJKoBn7WX7ustqF/i2g7EOh6fAZWBuFOFdPfj75Hdc3US
Rec0ekAzGtDXdBWym39+go3kuIGE1PjiIvSEmyFVIZ38l0tdAKHOAOQmxG5F/LjWponkkkj5H9VC
HqoH5ZJsj0c47PPbmgXQQx3vsGToZNNr8sPxSQYSnDx5Dlh0nr0UNpcT480pE2rG3WGOBLvm9kku
ezBLVm2Sx1bOf4SZbDZsr4yaodaIGe5FteGHRuKh4M/gXVi9aVBEJqp3qMct6qAPzDgyIPCm9SLM
zTGuVTFi7xySoZYSDHgyegTcNUpsUKSsnNw+VsQFj4Fd0VGme5v7c37CEkADFm1BmoCHtALHLP1m
vDAiyBsU0kt2njc5OL2cCjfdat1jxbrcdszftc72lfVDZZfKGZ1cK+Cg0cyx/VROuinfasOKKppa
WHvp8IvGb41ZXVobqrJ6rNRuon7+xSHxRB/RDJbG0PURZO1uwPqTxPjj/ZRwFbk/deYmEE3j/+YJ
HvyvS1nbA/FowQmzczw8vl1aXY0Ev8aXvi17nnVQQJk8IQo90yzArhBRnhkgvuzoYsZD5UyeoSZg
WN73TvxFkrMAqVpZwyc/wchwXWmGawFMHPhaj6B5CCx4rN8X8OnFtDCFoGbcQ/w5JYlC8Dt5ya2R
lULzoQgnjAIguIaRCpL13d6iJoeNm4IY5baTvJYmnTXzbdDB8XzzBdbCLTxixd48rlDrCQLdx+dE
dp6pIPHBx0EwsoVUzhZy7Qarw4vy3L+urEAk3dYU2e6RMVI+5GG+OcdSgg7bxe8i8rNknkXv94hw
Pa399AsgYnLGhlRKF9GDomlasfNUB1nH05gOtNlYk8GUEmEslRUUk0cqxFcSbL+iowtAfFhEKiuo
LEe0hlgblvsOOWEpcFvEN12RR+ZjBYUyI4wlX0775r12zeq6EFSTvhVfRRsUZ8RGXXREagX38sxQ
O1CRDD9Tg1WPyty4SK9+NzemRpKt4V3OMT4LWmrQHZu9gdXBTRtY2HyVBjEMTA4dY7/gVwNNJGiw
AYjU5+qvUvZmNM37MkNUCQbTXIAfaIRJwD9bq3v/wqX6pxFCoUVFO2sZiWSxRbVMnv7Vq4Jf5wOX
JWKQJvNfwYQZS2icmMBzn4D5lv3l5IVRMUruI2pb5e/0iyMqqqkKVC5G2ek7oX/QbhmzKcprq1vM
MWsPUXMwP+vLMInwtk24vDHeUJPLCZ7F1AwAlPOF4izoQ//Y8Y10VpvvXdmtZyl7yxUhnjoe/gPX
XIChIawf8HjZ+aRhGxok6X2CyWiFZqM/gU7h+VmxjlK/t8rBG/8U79hLvBw4RblRSS0LCT+rU4Tz
uj/WV7stIOpoJWnOTzxoxGgIBK8opi0hPjfj6l6p35gIeuH8Cw0JDWuxb027DVvlCafal1Xf7VxR
df5OE0+i5QyZ4fOPqCrXzk950anqdt0XhBUNB5i3uIA9Tgqp03gI0em1kqI7UoH2cBStgDpxAXwa
TeObKK3fTQs9ZN+/zYXZkJR/BGOEe0nr4y9riCHisOYi0o8EErKWZaHY63PEc1nltr719pOycAXT
W1HRW8tceoWoHBMD0liwtVAaMorkc19S0sOUNxGMKh8gQ6Yec/Dvsaep2VD3KNP1fX2/wH1p8bjb
hB4LTWHzxZtV686DUPy2WJbmgqcjg0kdhTRjdZ+CAbOj0JbGk1I29pcoFT3XGwrDkf6DzliQNwG+
VgdGlDCbkf0Q69r/IJRBcNyeQ4wEMegr9TZUsXzPBTeeFE3pDUsb3Z6zsw5scWP4eMdh2PSTWOj7
ot665D4z7fewKT+FfoYTkREGtu7EjdN59CiNmPs8CBQvs0PFiX6lN6fV6t3fGhjKTiUs3qGBHao7
1bT7AD/U+6c6QP2Hhcf9TGRMTZoLL0BNJ5cvwaGV4c9zTnOaXoeDLjarVgkzfRZYhRKEytzit3Bo
iS1UefV7k8xHBcYYFIJb3WMG9yEHInGwwQemr+FmV+2Uc/bLeP2wvGcyG/FtcmYzF+03V3aCg5lh
5JbaDrGuKeDJd+mIlVBj4dubn5riWtB4xBElUNyJPpX6OEEakrrsaRyMEQpspE7C3stc/43gTkCl
Qn5a7PD/gG/Ebe+RKgAsd0EUu0QQvoTjrcb0TSwxg/fwkrPA/n0ayVWz90Kd1m3utK5m2ef+oTz6
Qn9cgv5mExAnFuE9cY9NSIlO1xZUtci9sN02Sy0Y1rgOc0IAFyvaiQUURUHunfqvLUMmCMobLbpw
FMMDmfwYh774hRxk99rYTIy0IzkcEHuoHwBhMIE4O4cNacSEENE0uY76QF+W6XT/GHeUFkt4TzIl
1JPdHwXOyNwJxxG3JRwXRmaNqG0LUHsekV+IlfZmvzFDfMLhi7gy9zLLUw9+N8jElhOV/v2sUo+d
FE6GhlSFHutVe3PcWtKxVNzdyR+VLYCEW7WQSenELhnvGQezeoZzbh77/J5XiP24JFN18KAI0eQB
mN+k2MMyR9WowQtnkmgf5a/Z+zhaPyLrIy0FmdWSdLvu/APo/VlRoMHdW8BJktIpkzBYJUk45DFa
bI/Tp/FBWtQrQlUM6uEJfycEHH6xwDi2IyktOmp+DLU/H5lb1acDLBSedHCFTCgVOCGPB74nQ/dX
ma2/0Yv1rW1NkQWsbiYTLi1LmZfPyfn/NFT0LA4sQMz0GJU6rhtiKY9NgsazstjT4NHVpvvRyq2c
0c6DlELw+iGoOFgcNNiBxl6vKj+9ZHZ+kJa2qyEAv0bCM4H0AJRb+MjpNEuYsEhC0UFBo7tVmWrV
HzryFAOqCwguXrh4Ik7EMfgrhR6IsnIcK23LGHMYtx/UpBmAugjHbeQnFlpbYHG+SGDH7SbwqNiV
5rYtLxVRgZ1dTb2x7JjqCssE6t7v5nHd5tQfm8/CSa3UADGB75jFqtG7gig3yyUfNiuJmDp8jAeR
EvGLlOAoII1Bek5MJvDBQM+Ek8LiZmMvABfrGx+tvOP9JmTU+KidDB/cm1Yxt6qpg+EyP3oxAQzX
jM4sUSGKo2oZpceBUG2B8TlNbio0mCjVWjvDDPaCPOyCHBu2jmue0Ey1A3pCUcuSh8hLv6fBhheZ
rrxE2ijlWmu6IK2MoFfCqggQGu3k1v5o1fgFQAPCbkU+xGnfbhgNgoY13ynzh8IGWslYCwMFwKdB
fwl0490uFBLWabyccxj2TzzpoD3QkgKkZqpw4GPXKy7t5Vy47JyeKOKvML4i2bBmDI6CEmetq0yI
bbgjflLYooC8J6VjwmlZwrtn4B3G7fONY4SWgdIpLxJGAMyLgVKL8EpkOhU+r5KaF/uVbEdC38rs
7rIbzCVez9YxrB3anEGBR2Mla+bQ+VXx2AOafsuvCuR5nZF+OYLcCQJp7l8WrdodjcGHLguApMEz
eH/luTF1Ltl9R/yOh+yLeqkvL9v/jAs3dpB5ch59ffgSl5mOBQKFhWZszUGRPwJFL8aDHRUK5J5k
4YFLwcvYYrpGbi23bfxXRzYiUKfQR5d7Mzu4t4eezJgFsKcuWX8dcr4gnbxfGIY4t1Qi0VlF1BJ6
ekSJvZp3IEXbGpZVp/B1nCbk22gnQYogro/DhOG/+cFLEuSaAs0EGFkwLR5YqM0WRiX5ecMao/Zz
EzCXBk7OMQJW/4/veHtzoQ1qsUQLWDxo6Bf10gCZwmXYnz4yy47Dhe1rKP8DDHQXCB3JsbNJvvMZ
WsRymXqOCAi+AtouMw+ZOoiTtswRRaTi1zDsgxm4XlmWov0dbBlnmo7ee2qXThfTgq42nuMb2AVg
CWxKD+E7OZNSmShGruiTturF70JmlSj7CkNPnnyyQDR6+ibHSAvnS5dU3vOfClcGhUhI2CKNnbpK
KxA2OVvMUneDHcWKxiZbaARyW1Rzhxcm96bCyLtbqPSYVuCqUrMhpEs+Z2L2/vOK2h3HGwLxmqm4
4o7C02fgT9iRCkWcCjllwcYoM8rygMZE7iWNjCshXfp9ZQwDY0dRwFIRYaXj9DzLflnD6rHLr98R
aszQuti5av7w7daLjsYn4S5orv3c4M8DToijwS32iGNszfdoJ5HBMZcHGmJytFRk+DB8bjcxmkCQ
XrDSeFH4iBigixHejfii/K57FUfcMhb3di89Ha2HWmn7M+2mW+GO2pAGg8PG0LgNFxZbewBz4llU
OCzjavreY0LB4t5TOTnCZP74XfA1v2Cl8/YDePMToiDXarspGj2yUso19jVcv8oyr2Q43sggMtrH
ydZkuKF2BALZRpINTOjZH5hjaKDUJRUP5W0XLqDlyT4bG9ImtFpgQWfv8taPOlrK41XUCgP4+bId
7z30bxXs9oQRgC1TH/ashnYLJfVK0AT/a2EuuTQTY92Kfr4Xmi20BHH2nNmzeZXJzsq25hsU+yxc
63H/Ed9VO4L748dmFG6FzSMiHYoLmC6ltc5sLN0Xrd6EOUJpG0jq4b5wJNMkr6iCl54Uudu9qz6e
dr8PJYwVMrnM1Q3T67AdRWgfGvN9JoapTs9TK1AqKE4o8WMWSHPtJFFtBzmRrRDLe1YqsY5y7kSV
6sMtlOOa+r06Dw2+0p2oZwl4Rn2GEx9hva/sr80O+NiU5IF84P/xNoyMFnminzR80MeT+hxtbfdU
ub1wo2YMIlCkLjs3QZdtqVSgzLS4IbXVuPZ0Fu+nN0KIZlxOk6Jix9+I/tIiac5WHSC/Ib6AoDBD
lgxyW4pi243a3myOzsz1y3Wo4+bAYly+wW5Z0ngJvAzR0+nw3i70jUShfODFNHNTdxNz9SHQYVsn
1LTkkrilnBAV2qqxqxBO5FKHqATkQ+HTzy0dAdJ2kBocXqW2Dr/l4A31S5f11/lnL6DOl9gCjby4
LjIDXQSeCQ3e+eyTnKOcz5FApNHCYNiFgnfg/Hq5umzAt3ZWMsIgc6GWIFYUgk3C3mVt0EBDYbup
DSebYWa5hFYjTt6W11kYnY61gGd0/bJhLVgzs4VVWbsBUXz2KzZLZlC6VmjBvIImcZZeBEe4AVBd
W2OxNQQs8daJQo1Wy2OR2kXByPmbBpRYTRY+HpFkaf/6H4jfTvRUV1wTf9Xi0ohuf6/+yW4OdurR
dc0WYQQp6Gz7IH2xQ+5wcAMufcfLQJMs5pZpV04hQNLyWv619Brm51BKIUHC/RP6S0EKhvkeuU9B
4wtOrlPS6UCQRS6ok9nhFvJzksWu+ZQW0HWhTAcHH/JmomKe0xzEgBAG1x9NICn3g3k0hu8TUFlq
GezSCun1gKtTZD8tBb+4/uAWiBuDlQm3axCUexi6D3QKP2dWjSFQs12hSfDvly2f2DU83cULox3J
eEcIvFdQZww80Rj+oZhj5HJxN/sn+GYMAFnTdWh1yrO3fQicvjan+C3oHufaA29wPRXYVADdcpuy
3/B/BFvglJzZ7A4/pW/qOaWhcndGVJcIdvyafeNc9+7CzRO1fG1oKuk6Jt2+zmzreksR+GNXMoiu
daizYauNlu8SnRopgi0TiraPO65xm55rGdnuerIPSHJIXX7LhVVH2QM8jvz/1Xv/uEHYaisq6K+M
Ap44PFUSF+8La+qaAnZTIEaAsHuB1vwdrO+B874hZzEeFwebGfc+7OzJxkPjzipMnvujjC0L5iwD
/nSirAyw4fQ64JUyb8VsMpHHeynPPRY1M56EuDzK7GSKgVVOdrBQ0wxoxH4J/wGxDpjiLAUGffv4
YHw+kazqZyrvenFhxZUAYzeoGSvyeFu3+6FTh2BOoo2UYtl/MM9XB/SBNNaK2vzD+KAgHGH904Ea
WM/HUPYtqL9icYMmr4TNhvaKIagaTqofzRohzIEvT7QE3i+9YdOOBxDgZWxyNYVsxabij3hV/uKA
0Ac2+h1AvKI4V2tlqt2Ec0n2+Ta20soc99NXsemUxlmyQpWUsigt1SgDqVdQNPlfYCvND8IIL0oy
cN6WVrQmIsL95K5koSyPIAaLNaoYj8oR3PYY0tl06K6vVMdFCG4bPZaQdJN7a0DLV9EXurLJIr+L
Oqut0FsVEdIjfBwv/hewTvtXUGx/4jumYZib46fnaUPvFrbv/9Ia8bU7giAV6qzgIaQHg8vOQouM
b/V3IjJqXsykzqO7jPIheFwnd0tAGPMvDEuWVPK8B2x/rM0UF0cJo3krZrBMcJSIVf+TsJFIoa+J
OkhKGNiqan5JYjjNqsnBE2ZrLUMMfYsQAtBcMXesKEZl0cE+dLl09+gCC0ajsHpVDHPPWlmnUP/m
TQe9GHDbbC7iE0MCoTAOG8MIm6fPcESHzouCJ3oJoZoLVsGMV8aSYaEquMFNHEDxAUi/8AmTzBkJ
I5gx8Tgl60YNeuaDEZCuuFcT3rxhTIzC7qcHvwAxdpVK9BoM+4IlvUHTGZ8QW2u9OjDcQQ7oYSuC
GjmvHli/cvpgyu5A6HTEgPYHPY1aAK6YQ8yc1d0XNFxJO6ax4WyegX8XpuY/OyvKbZE+kVHAy0MM
cdhMa6Ik1UC8HuUAbtfiMnv15P8VrJAayt8iI7ukwj3mTZSliP1qOw6FVx/lJPCh8efk7Ik+UU3n
XPpsx5tlBAqtQo9IFRXII52Kp/i9wvZHgIwqJn8lW7y5f3sPViy9oOgmcCEXEiXjIn5I1JjnMlQQ
+JWv9T9XbXI/YXRRSVVtBzvtQs5lNPNbRmWJV3sgmaTilffKtSr8TlCci3cIYmDM9R8M3j1nnbQL
bNyzShwtkeBlvBI4jlK3aAPtywHj2X54G/0U+qmJXvB4nn4tJ1ZWo6U2CiY67F7cIA7al0ohLfTP
YHMymJawTd2t3+d5wEiwtfUC+anA2c8XNy17SNjKPGrzwqv4Uk4v26Ac300ghzg8+hwDOoI1ODGS
fPyjcEYG1Wu4prlhdojYcd5cXnIE0rHYJLUgduDHOAtmdyEDynbCLpeusgTHuUq0+DbLkH09F0+L
JQOXQO33OgOO91UZHUDAlLkwd4EO2oFZLlLiL1PsqbpCriOGggPAOZmkcNPFaqOZeIyCIZyPrBYv
ieamBHHimshyGKs7WpL+6r/HJJprGQwbHzdOXYmxDmf+PmNJ+CgCC+az5HO+srFqauAopVhYYvve
FstPiZ6eqHJWTufkpEOw1kfUkkEeesGNdEPZppToMFTWLcMdE2uxWLEZPBE01t6vJPbWmqMIrg8J
gn2EXBF3CU3ULkdws5aA5w6k/oYWxBsG4oC7pJpBLtgErdyv1XnVXQ6MamYg+qB2H3AQzhd61jzy
rnObecbbZ5+HZu+a9Cbf1iGYTEaiB+opaG9rbCjNroraiUVMmlAm5/zqsnpADZJd8flFRxBuZQjc
qoFqLOLZsuKG3ymjtVrF87i/RyFy21japEcvM2Jt/Js81lYY6FH4YOwN7KI6s5jKCaCGV0NhG7ag
TF5sEopVgIMSwmw8hFAgwgYqUToJEFYRZoxVINq7ar/wSkCpBq5c65QwdCidVFg0TOnLSbSu+r4+
+qvFgaEGktfiL1287UGVHgjgODwi0dUvTlB3qG7PDenUNe2CR8VLKpA7Gp9iFcDNlGrnAF4t7uDL
O0ByqpsvVODTDMFrkBvLlsfXC6zbz3w38tnvJckRmIljrbRGrCRntSTmVJSc5e3257v3Tg3yKrFh
MYDDZLQJ/tTJNgPPxPfoAmFjFil41f4YPGIMiXOABcMR9jE24xNWcCYbXEbDrFlAr0YVEYHv5bnF
hKmNAubGQFlba3G1a2XV+7CxafDx5oZqQveV5t+RXIaiFTi/5T2ZytJORAXvkkMRl2LLT1rg62jA
mRzrJpo51I2f5VTjthdcLtsWMPc37bggWC6JFSIKssok4fJlXj8kJhz75k7mh2vEn4leroPIecv3
idSbW7s5VtvnfABZtZllqFijFG6lGQrDE8frJHGbn9j73I2IR/7Csj7RCcWHiaAN1oIVrU/z9+70
5I6OwwTwtA7hhw0eeuH9ZA04yGSLsfTVvuc5KwiMc9+PPZRSd7/Eu7xK39s+5s1z9whnVrBGwr+x
UzHWfkT5yeSOl5C6SGcOwAWPojbDZuPyMqqM+nollUc0PxBgvmyHYY5/3maYHohXd+Ff2cHx5Pnj
qEdU8RbkmaTqejyi+DFH/hNvJ75krOQd3aYTYaVkjvzTnsHGl1cbVbjXwSZknrXngi/c89qstR70
ultqiAxor4iyctTLBUZWSuqM61ba1aBZWq1C8K17YVzTVVpzXo+Dx/evltAnUzN3IKgvuvf6zCKN
ZsOblsEk1um3EUAVE/yipFpbdcxYKVdTi9hyVdKpMpusSfHtB1IsUt3T/yFkuxWc+5PIIPrhvMO3
C0TQ1zLWRTL5G5ftoO1pDjA5r9QDjDLv/3xXcRcSMp2a9T/xH/LLLD6tLKYXaDMxgWX8H6BS2K8D
rtcPKLCBzjm6qMc+Ky4cNmIk0AJvLd2JYHDw9xJ7AOh+zVBAdpFE3eKgIhLTX40ODuxQJBYXoxyn
gkpFnTvUFDKZeKqA7CXDo6EyYKpI30F6Wi3HFXcexsoJC2oWlIROsHTa70dfVAUogaq8f4Rpotfw
PJey9772bk61L+ZS4/7ejOYqfnq7TN5VCLN5wBsTO0bPW62bUo137Ask1hDghCWIBb947P2uv+p6
2oBu+vRfKlk3kq1KF5B6x2Kax6v7+XsT53sZENd+NkplbrvPP8kOP3Omo/GGLCMXR+kuI3IJVEzH
b2x9/piAHzvat1rSAeNi73kZOd77b9xnysNOREGS5z9K70sgTIc13HKLR6DGfPKEOQBsfXMjsOuc
mavU2KP3hks0Fk7i1TqMsc0SLgk9YpvXAfZ/8roinMbjH8v/3WaG/rAzXyUaGUR0CzwjXWZf4mHI
ueqlRkCE0aWyaP3LOtDf+EpebVYhPnv4Z+lM8zfQcujhBwdm6z5qgBEft85f05buQdznRm9bh/a0
nDAqEvZKAZiW631VPN9czRNp1MHMcAPMMG4vfHYvgZOaijNsC4vWKPSoW4Hp68fyAzo06BCknS6M
3y070NCRcIZV020n+abrE6/06meW6X3UUA48RfwvNuIZ8tvPsXtn4mEWJnxVOi9kdO0EpQqNc0UN
u6Mh6Ug7XDejKFf/BdfC0PJOtjvTVYttWKCn2VrWo+Za27bo1SPXdEzcIOzDaU2AzXRpBqNjkY8Z
Am4TEoVg+V0+CzgVfiiohL+YL4jMTWw0VtYlJ3KkReSQ2K9cy4eAsw+J0yHdfGEwitei5lyEP2gx
Use+cj6Vf8K4HMl5m4wYCXMnVJJWm/hJR5Wp+EZbLoRV91SMbTlT7UCtZqHPWsAqEr8chSXB/vSu
977hAdCnGFWBE3fDTnEKDwT729+/Ubp1c5ljQNEnMF7iyyWJihF5U+B6L7ViirKBecw735Z4c8Z5
yQkfQdtY90Ay4bqEbiosu0Fj7QjMJpmsuRQC/dw3QNQRqCpm2uCyq2xLdxJDDu9pkHBSMpdIiMNC
vbyy2bpAMyB2FzWkiVD0XBklGVG4YkxJr8WAcuL3Yf3Y8OiBmgT2jxgVpO5zbljPDJtP/ShhK87P
NWrGnpiNJf99ky738KUW9dG6ZvcKoB+1EMt2SqX+zAFelQ1fVQwHyqv0IYkqFSqRjXmR0Iuc/RYK
ktAZbYlKUCpDk9RpG0T2CJX8PSziCvKtRA3iM5bXHbK6bKSVVYXJAOkubW2vDSEjCuELwwnZZ5MT
l0V75O7RE3VWJTQYEZJx/MKy66rMuISUOdXVtXpj3QyCLX2EsxcYm7zWbwak3p4n4QBkU+Pc7cY3
S51pVnhSqqRocEjWWBxTNi8eY68tZzAKVWYG+Uve2XZ+PFV1uf8ymd6rTd1IhH3u3n7m+y4VLreo
KFNtbDc5TxU+3OnA7koMPfJjjqLNf18t3hLjDC07YlPcTsPzLtflRqAePWu7OX8ogNr1+mWmPCsN
TE8YtpdQEGtcQdFSQNoPMhCpgLlT6Upfu9+5nRtdXt4zHYNxRUA02bnJWSMDIoKLvbZQ1JiNCUoy
4q4K99GSxy7mvhGO5IkSiODDlJBitOT59uqRldy0FxBGLdPVhyEJy/6ueX3/pAycmLyOQM/EOX3Y
KaG3FU/nwHBmAtnzV+MyV2Mo7nKKQcEgHf52oczg4r5GPVI9Lp0PlO+axTp63uVYbXg+fhXMyVb8
L2ts7T/3wLCx1PIluKzMoJsmDZ114hjFc4m0W/MzlWd9eQF0IAZ3/Wr27BTKGDKr7GDfk1+11e0f
RQlazl0DFrOrnc9GRr/KZPkigIRWAtZaS0EqO5fGVOp5oOH5gHVfQO1UMa18WvyT8RYs3Jkah344
DyBbjsGWVQqc/Hm1x1t4afhoyqfu7afdm8DmTqhZeK6FYqvooDO+Pjz9/esxS6GSe1lU4Z14TfFp
0g7YFmzDJDcL0w0Ts+KBWGyyKovkkFlG/WN7UGd2SF4yc6co3BBGCvrjh0nz8HMF7xBWcvPxvvQW
BsU9bSEPtrnGJL3Z1u07N4QnwWq58BF9RmPDGMMZsXXM0GQ1ZSXTNi8avSkkF49YQ1IVPY8K7QT6
bTc35NMfCxZREx2bXdeRo/Kj1y4RvlbilKFTcjwlNqn9gop5tW1cpljKsolzmlFfjanPjDivzQ9d
LyJFGyadGUcmr+UQNkev6QvQHQY0YjY2jy75xzTns+jfHj8MVK2Kw+LzT8AD1yC9BpRsjn1vKnpU
XqlFa9iO0R0eYVCG3wwb7vLcqBEn2GZLB8AusSOjkq2YgagXJXUbijA/kPWK0NcgsBKvRqit4TXH
sKOXlfrnBYAlqngfQfPjFDFfan+K9dafzsioda6iPhPzYhk8lfcSQaVjRMNGwL5gvSNkvis71lSB
AWX/Dz0v77nHVtpJ58IzpMGz/g3ulqA9JcL8B4ka3YdZi1hiu69e2K5FNwp9gqNMRl87lZ/nVWzF
1W1kTe748Rk9LYpsUVgKkE9bHH1J6tor4chzjUm8UulyxSq/cDgn8KWkj/sUsfn+/X4BaQ2zG8TZ
ZL8ifETpxKTnXah4XDQ3HcnoZUJKUUzlNoyCyNQJ5r9RrNFVswQ6H2rQcTcX9XCZJZ2PvweXbLIo
YQUYamVd+8zCoI6MTm66b+wqJNLiuHp+b7RkF9f7dLp9i/b5zgMnJLoYCqdmI0MNuZtvO4AMGSn+
XueoK7G9Yl666qzf14le7sgQdJi3ewdXWUIojttYecct3eFlaHu9CQ7eRBW9uifWsBcqTVM622Mf
DJLGpgBDZg2RzrAyYBue7KXpJtYmYeKoxyBT4eCh7RzZpS04uWEQlSqBRN9G7SAy3wbnrz7wqL3o
XkaMk4o3/6OE8H9XObwKRTK1IwQkbRoRBd+5/g34j8WUF2pNzznvWM9Lvrd5OKATnf5kTr1Ghk/y
2kCAAcReCyAhLAU6Ry4W1CfiIGSY7t7JFnxQ6TQdSMzaOxzl+ypkGHIJDOpRg5KJRD6QDUbDWpkX
kPnWkSPVmRJazHSZglH6AJ/qYJ4uNwd2Ts1g0NoMogz6VZIql9GXOzyp7TJVHy75VBtqlfRO5d5J
6a9qbByTH8T+Vv+CC4bNT3KAggMvpvbjwLDXLydjbSiGoXpUcWKBAO9rdxqURHeGx25XfRlpLDQk
7iNhJunUQK/85xijCmlFwt6DHuFlRSYgQGqDOSgRk5rJxpQQLaCvGC9LebGlcPCznsXIBKHnjLi6
FoL19XNxRYMDLaPfgj+sUm1W58gnxoUhurJVdx+fHmg8O7GfjBVkMkt3++pEiNzUJlDSoC+ODxSl
hS8PWUOanCUoT/LIwQrE8wIvOFkPfHVfzufnH8FJ20BZX244l85YH7z5RRqetzBiK7WA5WS4zWae
Yo/r/9fLDBFIlOaCSsuO3toJ7ypMWzxmXWJBWU/OWn/QYeonfycgmBkenmnXVuFJjZ+gwUL7Dyy3
NdyvpUKk7dTD/pgD5lZ05pbPPonzOZqm1d+p4/IEOfo7orL7CENkIxucYNYNQ5czvbwE1oWQCQny
rERpb53oukHDTmR6PB5OjPPLgSDgMxDZu1My9kfnVPonXSklffCim9UHtMs6QgN8+fjcSJ2zmNF4
S/qnNt6x1DXM6oJycO3U7ZrF2eqqU/P28A4Bu/k+zhodoOrIEvclCn4zih47J0XVj8Bhl2n0hq/I
bfZ3tdfoGyqu9FGUVfz4xG+KDl4vULdUlCByVh+WsAazyqERk2LoyZ6Dyd26Kju8t1WHswF2wGjG
1lfkRLWDKD+rtE8ATKdU8/PfDiJlTGijeiGgR9h2ZFptfwhmYhToDut9LmVtG4JqiSrhUHnrgSww
vDkY3uw1BwJZ1dwL+o5VNEXshEYqgQOI0pVRD2pfS6OFLVVP++p77TWLZXuWqdWF1jPROKn5Hppq
gRTrBlPOzwRQy4wTfdONnjdaJ4dE7LKM3MfhABSUpwu6TlYPw6+yYjd0CwGaVvCzLxYGwVN2aI6I
bZchvBSgOhP6WYgwkA+yALjAVv22A56NkQB0MUZkPALNJqyVmkfxSLQ9jF9E86GeozDdvr6A0YEE
Vl2MPEgJAJyl1BUZyysxhQc3WJHzkiQcxzBejqzDpxcLn6awTmhzTG8CKpC+3nn1wzKrH2fUHWPG
qDMtVekaV8kGP1vkyOdSF8L/sZ7nxRW84SYRsFEBihOqiKX5iTcNYutofiOyc1NSj7fIYUHCW0M+
ka4ydsyS2+ZLvZ8Q2bqAcMcuPA9rzIuYYMb4+0uxrq/h9WnDzKDGtUlyu60MkFUo1c+M/C+aBi2N
L1FVSUEE1Z2C51Yo/MeIkdOxZgcbF6Vsf3SknJgrzMOIKYDrUdhyMpzsur7w/MRBYDIy4uutIp0L
+kuQR/jGcEQzotZtvu2FFElrCQAOcllBKQv4tFBV5I9cgK6G6Kkf3z0UFZOpfJwmGEmb3ljrITzP
Ox/tz6uA8TkJBZjDmmxm9iDFdF8WQ2uR0HqVVLOv3LKHAoOM+vv/KH+D39G3a4lHTIsLaeYpN4tM
tc8AgK+TdPjgK+RcsXpKEHDWAJilr+WsDriNaOvRONjcwXrDhsC9hG6BzBY+HdgTUojRbdYCmX6o
dwgIVlTJeWmuICcH7bf9CWs9FoZzwWQbTbUZQ0eM19oYBxo3mQEseAgEUtvy7DqQ2IJKbtDP6nji
lt2H2cHeZTCZ7MG5Apv5v/3c8Ow7OH79qyIf5trudZ56iGcc6RpPvi0c2e34/Bub6G+G5KzDomqN
GoNo6xZoLg10sUHdWhmB074K58/Wp90lw+MwqT1NYSpUq0Yx2XSYumb25qVwMtZbOw9zxcTrNn91
kzLv8oOSXVOXP7PMR0UzM5e33MfX3hkt9RMMAVKyU2AZ660mNCfOntAIGqI6G7FlYbbBBANA4xI+
XpOQ68uRmObcLO2ClBt87Agp9KVzf7YCxby0ijjybYuqZb0s1zyD9IaS/wWdfc0aVFtqh45jTfT9
X6hhkrKJb9LHFw6VFA5bDSeHjGem5RiKxCCQQZHC2Tf/bPfBFMY/iYOZzy7vb4eerkB7ZlCIsP4n
X4LELAfsJGfry0cwQZHQCmEKUgLbUQT1ZmoshToQBiewN3i9elxiTfvyzBXYIeVHzv/KevjFYoyI
LmLjKpUZZV6wXS1Tm5pTy51lSY5O43pBT8c0JsSY0SQ48X7uDXfwo1rugCgaS02SJCXjTillqt/5
pw1bM9SEKRfQv9k+6YJNSL+qXwkao1MEmCT/kV803scLlBaKZSIEL/IuJK6/otAS3UZ0SwliUyDk
gAjLmawGtybDQEPxMZDUjaxNeAnxAlZ6V+hDuDsVC+82fuSgZ86gj2mhsqffDkJVRFj8XMWju1bU
QRGSDDuIHZxSYtCBCbsbbebugisoFGjhUYAxCtBrYqm6pfxqrpVf3u5hSbd+UP3jRV6oDDiom1LS
M/Nr/68Tx9Ud2Lv/Zk487mG8Sb4iEXKloXp6sV+OPwBjQLq9WEFfhxSxk7u6waY/2hBGDBIlnc/Y
0XQ9MDyURtCoLXAwL2tBQ/mpj1P/1KIPpHGjW8qNP5ZveBpwPkZO482+zDATR/8NT3+SFgdAT0OB
hUlS25Z7hxDPzg67fzXI5kwftUOKcQg9c8X4hVDSuyZq044Di2yrWpSWWz7Jy99A/JD07LV4lXnA
Z4EajexZ0LlJgjTBZFUcPjzCoN2eUNqe+fR/YxTCgbCZB8r5iOcsyAcF/ZqRXxeX+/HuidTWTd3K
vcsZ0q6kVijGz/8FTHiz8qUvQttt1b003c6rT6dP0EnT0hhLS8/3x1F/4LmlNC7bdQbPXxFf92ly
R4tyfkOssgKlztti/YTNcWhaw1SuqfNucQBZZQVkIQLwPwsU+QvbC+x1rfKu+2W2Mp7W2gM07f2x
P69gc8jMTkg3yCK+82qQR6RcB9/TUfUADQyZYr9eDP9sMex6q1UsAzmfZc7ARY39UBrlXM8XhB4a
BJtQpqFulTXg2NoldqT1MHR93tuSPq2xJEPVCX/gMF7oAB02jYea7HOAuV7ifVLAWbmfBM5HqyZw
+6D/F/+LDwD2ksTJ4ZK6An6PZTr+6LBEeO35kLIlIDw7Fr6T+Kfd42ph7WAy9F0dKeHlCulgiCsa
6QOvIE6hSS0tdomqYjYBoUPcg59h60NKS6evk0aU3qP58duLY5nGOMlb1gtv6OINSBdYhEilR/Q2
LFYzk4G9l0ufvbUD9Yus0yDR1wSEOqI+yZ4perRnrrKd4UGCD4HG7+dFkOCDrk4xpmWO+7R3TxJH
RBIDPuPCK3PQAs1WLoiFNF4yHpEUvW9HFTrvndkbV0slxAXO6cVgg2xrJaOGZQQ1SH8f4pzp+ftH
guCJ0iTHjpX1tSpeglg/LhWUlqCv9Q8UoLyUdb44WSAoA7JnlBj21go949nAiflHrJF4vnDYjQ6u
eTKrWWvfPlqeut6gb9AXOzfMi2ku+twASBaRHoCUebWZbvCTSkIML8SVlYU14w+tIc1T32nsodKp
noDwsfW8z90bBBYeOMp8uxvmbPlJm1uXXj1wlBQFmrhjWy5ypG/IDlf9L/DUSLXfEA0Ewmt/PMp/
NyuNh5eZ7EdvTU8n15LclnoF9SX0DCsGwmKC963WARrJL0e66JJnxr2NXV3ZYQMkKuBMix+2xtGy
d7ef7Ue7diVAHIUt4L3F1gCG25Hoz0grPhzh14csGqhinCymTMeJg+Yr3aHodaQHRXS1PeZfLrzQ
8vniDzhW2lSH0cTLsDwEiZO7mj6xKi9MUMg6h9sEkPb1aUzv29lg3Z0mU94uaViTInixZCUi9AaD
Lp4Dnoh2MF4XgjfPSb9qxph15ZJpEvWjMzxuSLw5Z6c/Z2AdzKT/0Vh/xw0sOA/M3ROT8tOjLKQC
BwrwykawP0730lt3n9ggRANrB4v6lxNljImFQICbO23Av9jHLfyaMrMKBCDwy8Eopk5zR2a/DO1T
q53JoHmIQMaXYKc2QgSGsGYfbxyXWs+QKWwbObbql8SLokQvgMzxgCTQuRHC4FrBPicPz4oUsb38
GN0KpUU5GqgBgK7BMAk07lvcsJXGJ/erjIZ5IWOgogKAG20UK+h/YX92UqSFlGCMMSJc2Y0197Re
eIQpDCN99CO6rfrdoaNtJf4uXTiBbslQkI2U3C+7SFBqig0xD/DfK2PWIKNviGEk0qEi9dfNvSLW
sUKmDxrYKuFWvtLp90ZjBH43wLHXWoQkZjxBKxJ4bK976hUlCY4Tvfb7mdoh1tAh6dU/ouPO1HfJ
dOzaKpnT4shxBs0rwt/wk5/VFY28JKmza6b4IUbH99dPRnazP/27+f0e7KxQINkeKGLY2ITZncuI
CfrLl7K8iNzCa6VMNBw1y7S+ioeTicRhRDY/8uDFrAhJb0gtAkm3uMB+gCFjDrkZaVW9woeN0wZS
A3OSyR86JIGdMz8DHZcawtkxSOf+rrTpsrnymeYbcb+apXjgdPLBAB9KqkNORA5IfQv2ig6cThD9
585soEneZhPRiST+7FXoPB8zfNkqT9MyvmZv0CDUkrD0aUCPol5yNo10tjoAD8dbOFkmHqSTOiJo
8f0O69uOfrnqXvMwxOd84lm5L3dLgWfv+bkkaWMKL2k7wZ0Q1cSj1+BK/WyrLRfN0y41MVSjJDvU
M5W3d2qltKZ5Meos6GChvYm8UbxQqLWMi2jWktGT6EfZDDzvnPgCIBkHMnpK7ZOsLztGT97tDn00
Of5PEo66OZ/J1BvK6PVOf5iusYiK0vABNMd64QiGxYbR6WiQ46S9kPrAudR4ALdbgO4nfoo8jdTH
eyum5ie8Sr4/2LzWGBslR8qXQZ2TCY95SAUw5eFX3U4py9OrMGfqq3ODFgIqs2263mw+889SolWn
6hOneaEgo0XhggxItWobK9cx7DXv4ctZAN9T5pSmNFFHLgE0HPa6DhX48NTNhuRYVEZ6HpoIeKU4
1WFhJgy9W6HygGycgkLdzk0eVPwMJPYu2lgr0P13hMIe9iDCxZHL1I41b3x1LXIB5Ov5N4KzxaS5
jEjxfd9qLw0NyyF4vYdsedrka0N+3kvatVdbZRHu2rpJgp02yKn/hoWBEjMUn8MYy7dZOXAxaLle
ksvtJhQgNbLCFxfve/y50m5Iw3mpXvX0aolTpyn5qqPfTmOfUAbPmzdD2JoWu0+B4m+mTWDOSAcZ
MXDxyi9iqIhSGV0+DwAhS6fMdqZKYsxX26olpG0gl0zwJshwLLWhigSdAxYcuJippnbzl+MpjLnD
YxJbSkbBRydidTsrQTo0UA/GMUK8HAKYns8EzFc1dD8WBHGIWPFo0E+p/DRtD4TC/wWxewKEtwzV
ZLezh6PPOKfzJXZWB0za/mGse+Dm5ZdonnEuEWh7RlyEHfydcY0QL7ACJe5rwh3T7MO1WCjgW5tb
EFDX8IUU3iuadMp7svhmibU2Fokq7Y/kyaZpPsJqkw01uUwuTghpfo73T9P+W/JAXzMkvVsMxUX0
YA37F3FAeZCf53KKpUzFsvjANP+hR7VGXhRO69dFyK3lQLnC8Ch+9td0GbjpvG4/x8UoUMWM1CVS
DXTR0a2imuuJ7u3QtF5NcBpoSP2hoNNgqiigpIa4lpoylzK7p//d9A2y4lp4gyuCHyIyf8j0Gp3k
g6MpljjBVfI6BPBh5nl2UTaAj/7NvN6DbBMrgTrLqQ21G6q9A4TvwCn5RCKT/PBna75pYwPQJKRB
0CfmpMonA+lxRd1m47XTQc1Qt6ub1x0sDM0c7CpVTASbRGHrtwy7b+nQx/lU7w89ODO4QMk5j3nV
P+tWFNUEuF9sC8/xFivwvxBK1sUOdwVOmL8hY3nyw3Vd4Ei39Cma0unZACvQ4dzfm1fvxlsFGXZe
G2XZxCxzQSZPu7KQz+Zo9i3uM9Lw0hsup3RokbJvpPBgdsBMJrB0+dpMi+Jn/1qvVu84uQLZo1OL
KyTNhyJ2VxDsvUjcHzJ0vUMk7yXXS3Myof8jBDA1UtuWB9EsLsKTJfejg9cYpylGpP7SlZ0fYk3T
As/mWHrPs6ZRD4+7FMQu5HuW7mKuNiHmzsoIV53SGil16zoccIA2CvmADgffkmFnmkk97jM29WoB
TNPx31XWT/yw4iz6X1I683ziuhyo9tZKZhuvd3uP+t65sDeDlAJUjIjYDe+waelfr7RjOjnJVM/a
petK0ZP71OLkg6yxBnatpa9YIT+LykMLfEXMmNlG9eNPgjl0QpbB6moG0bKxq5wIJh++kv0m9Ilo
e3YeJdvSP1Eh9aiJd5AInfOcHHf2Hfug1X1z0SvDXAWc3jaznZ/4k4gqExp9601P7xrGUWQ9tf/j
LzlNafOyc9RXNT5usVa76rn26gbHRKLHdu/ir+UHhgX8kG/wFoiJ4/b7c6N1djDngDeTCVy3XPAR
He3nIJc0dlXJF6A3PNLaToXDPCsHiKsz0W0uhy95Wu7DZZoiMRhBS462HGApJz0eUfuZtlJ9/lL2
au6eFTQibZEAnXcFrtoM3LQNV5RFDNJg8weBq9smBbZE8QTwlArY+advqGOjSzljQQBGhAMkN6j+
kCG51K5eE4nrVmPJngjYz8jhb15nFM7FVc2upyiWsp3gu1lax286eMoOUuIeu2abYSOFkQmOQqS0
x7zy1cX3RON8PLra7HgmGMfhqXSTGPm2IMGoTrZLcSdRA4aVz+90icO+HIqXZMPmGHPqTphyJ4zb
t++geaIOWfyKI4S6E0EvewkEEi36DcvMiZ25opFwHWoyFjlWolnZt4F5fPZH9V2xll54HMcrMYvp
O3LbClJTyUkfPZ+zS2xrF+WLKTdlkQKBcf8WlAMXimHadZZEcLEqK+qRhLwqR1usRWLDXyq4dfVD
yTjNG8isnQH53XMObmOwgxzW7hufS/RLbjQeYBwJxbxJZBtXt77Fslk9aaE3HBLuFheDzJ0OrSXQ
ho7CCk/CwlI+P7Xh4GUQonuQuCLrqZtZCzJ+Qhw7CpV48PE4XMud/nT4+wHd54nh9q4GrQ+R8wUa
1yW4kVRa9Y+tRTmgR/6MkNo60Klv/4ISnTvjGhUKf7a/dSRe7A1OjLvNk29GWVWuE1ylrZ6eZqd/
k+2DtSjhgNsKDTIGSySHBVCFP0o5WlR2iwlGKTvSmUSRPsBgPe5l+ElL3XJfXSFG4OCmLdP/Jl/R
YiCJ1hOj2HoiQyT0TGwev+vuA2pDOPHLOpxpVgl3rlgM47ZsqugrQFQOgWhUKGdVbxVyxv11nzLn
ViJDY1TentrfU8JNJQaI2AQtP3xdK+PfgOkNKhAOiY4z1IoiPC5FQrG84t+9IkxSNQt9Ot8YXDBt
GvC5XybTzekmAS5QqQYD+m6rIqNKIV7mSZ4a3xyRN+zclCefx3xrTseHDOVfXPqcQV3FaS9wpPvA
hR38mja+677ZmB5yalwMVkqgQUyAC4otPLu/PmHwgo1usAdeGhHoKUFhmFgplDp36y0D9CHr0FLQ
N2eMRLLE4oz8cObxWj/spMGtEN+lTPMNgkzuLSLFX3Lt4NgO6r+UkLMrOZmdtSzllZEk3U5QswSX
44AA/ZBlu/VYWQBUQMgzCFRAeOIDtZudeEHpYExR4Z/DfS/gVkUNJi79630u1+iVRbL5Tl88+CgX
yPYlii/u2kSWOc3bxyST30tqIMxxxUwtJDFb8Pgs65OV8aLpEUSSDLi9udkma2HWau6VgMt0JXWC
NhCDvoCWLHBJq9dEMm3hT4HqtNmCvE6BbUShkMHPxM+HsDqeQ+yKAjEVtlVA0focHBY0JItZMnG7
yrdTP3ZfudckSTYXGUKQitfHTMPCJJmccgUMebYTMcFyrLDWtMskPy3hoSTPT+lI1bVN2ojrG+H2
i/jJbZq3W4r2KfXjQsNi1uW89i4BTO0t/QVwN4CvX5VNKaltwry3f8OiNjP8Fr3Dqlh2SCTzzWp2
OjQwynvB1EryQqPsBvMvi6LesjP5mYAPGdQdai27KCgiuiMUW/o+0e10fB2WYIaLxSsnaCf+l5Bf
8mGJe3WeRM2+kcjBWIpvXGHwazghOZQbNzOlfLzVgKmOcTNjO2LjGEQedWaGpYSGoa+TW0ShNrbO
5xFkgs8w44lx3CCwNvERa5QyEuuJfcRCHvf7VQhLjVMQfjbF8+SPP5F/tT7PJaKJAMdxIblhfHPb
re6+sSCljrmDOzaSqWdDaKkgx+dSOwKOQigvoHFJ/WA6xOK+FxkNTQctpSxI6lQbTsalxTZT4prK
VM3f4HEq0um0dq+25BASnUM1E5rqk3c5lPTIEbkrwOLLxkiVzL4T3i3xCDwy0cQ4h1FOKCGU8RdV
j7nMGUg0aXpOwy6H4Dfw5v7KHBjVU41raE1m9a4CWzg9Ht+dRiZsZBEVWrrX0gX1rmIV/PAmcU7j
nS49mroDFqBM7bKXARZiNCNS48eYjOFVzAJ/8UXHb2WZOdCI5nbb2Aghaov3Nncjwt5w9eOnvO7n
9+D0CT0Y1/J4looaeWzFI0o49BL+GFOOS8AIen7kKYnyKm/jywtCU6l2Dr83Xu7wClTgyRebxiZr
cbxcBQ4YIAjvSvkVNw5WRGjDxDAelRNgauw9rxwqgjJd3jpeZcPMNhymoKuC3kwht2B6jZw0zZAR
RcIc3z13Z0dIbLM1vnDR1VKPN2CVXOs01Oe4VmnSx7cYk9a1QScycuZBuagH74CyGMWQxfPnim7M
k1frHuJjRJpwdXog+u6vbAR1J66aFviG8jJscOqJvKV/a7r718HT9ZcWX6OT+4QWMd4xo4mCTH2H
GK5QmYXZXPnh6YsG2dNdquDiSBYZfIXSnKhpP3FxsCW2kOpwUzjio1ydm8hw0COxdieY2BpkG3Fp
bW1LDOwGo3zTOUfmzcIgvfA/+1R+SOrqp6cBmzK0DBkVVCqGfl77UFlf5Mm3QyuoghabtdA1SO/Q
IrtwDLnwgx2rOT0TXYq2++RmJR8tPUR8nJQoecR4z859ZiLABc+KSp7Xk54S53cknS/C4hFNAg7T
Sv6FtCIsjedApWG5j6INSOWeZaSZWbOaNXaqMD7EkBh7RALlVIxwQD7pS0vqFUtqJc+27JCZPnkC
jsmRzUs+3BPAGmz3UIOSABZyIpyUmU3V/oYUN6cRgu5zkqDLUWvd51P/+oKTtG3uuG5JgsD29GQi
Ld8sBTta8K6Absmlso5hx0xiKX1GdMxBJ5uMW8TyAUfRp8L4K/KuhDuvrcCaONPoTBrFc6aULXDa
ZV8Te2s0JdbLYvxKxFuDg6TUb2XvdgrF8ElvDRVshnbJ1SdnJpqztASrmQijF3jlgT2Emk9L8nB7
SnJwkB/+pxDf+9fOLTeAFEBfMH+JspkLL2BZoy1TXwvhs+9QldpLJNaQ1FJld1ipIrjDTQuwBNzV
A/AXDN6ZmwzRv5yQHcMKZI7YwTz9zYwCDyRY9IH9rjhUY7tXJ+YVb0qjuKjxwW9DbkigqGXw9Yye
1POPWHCRISKqgDWGwKAOS4FV7C13/9UxCGbUfw1E3rywQn5++iUvNEAPpO/abTHW0NYnPLx/yEni
YJXv+9IWGkJhmQjYBAgKMsO9OvDIaG3ipScXJ7h0k1cURjJ+5XOFr6dbN8IFRH3/a9/7qq/ZsTXg
T/sqzERYW+7bF+8BBjTR9E4ZsUb0Zx3L28Le79yNzkmaGhikRbfzgF2tDo/YOXwq/6YvKAclDDcR
Q0cPKowImeK1o5tTyYLdTAwIgpuHlCkrKSlaVWs9Qi7UYH2Yr7ihRPrE9K0o1PJ0suZQT7B/+nJV
BlnIbENCKAkocoLZ6N9ai6G4ey6ltEkP4BhnEt0iPg75FZIg5Bg87TCiHiupjy1l0kZuz65XPLjQ
C//G4DTaCe6TyCF3rR+OO1O2fo+fwHfPFCj6f2Y0P0Kemrs0oV3RXQZp2rHVgyfXeEok5XzCnkRq
tfKvc+jrziWar51V6Ds31qwGjau6Mmf63rHTbJS364eo3V7WDzwK4iIOpvj+2bRKwc4ybSHJxzDg
br8LUg3yrbnuUWO7f/56lJxkXN3RXhWfcUiVhWXLsgmyMfmP86SER1efAPcEdTU27J8kvaYcfPE7
RtgGpdscTHjysg39e4ybvjDG4iCVj0fvJVVrgfdIE+Ho+EAhY6adveDUlDWcXXdojE6IdaZko/Jc
/8sBQlth7JikRnN3PTfTb9X/1DaHgbzmBGesgFM1GsEhfLvbaAXOv0PiSrVPPjwZf2oSS4MkZtJY
sk1KHbqcQWBIyL6YDMQCreXWB+EFaH795g1dGoUPP4yHnGsiiqsA9xijev+roYlJKbjxDpnz+WhF
wGIUajyVV0ylg0CNYK+NQOVQjqZIWQh2/xz/QufmmYXTt0El8xAog7pvPo4v6or5OfbIcacaQild
KuRVblfQ8OWjYGo37AOeuVnGJoZaHAAtkzn+auROBX/qFJoDc+JKkLLMPnNvuMGQ/si/Dar7nxx9
UkXFucc5xXG2N2O7zboXYHaayy2IUt7ruWNMu3yv8ywisPj5pYxPNMUv8kM0+G6IH0bKEWShlCfz
ZSjf9UtY+Nxf1cXdNpA3C0NJeALtU7lGOzIECHv2Z/MCIajJeIoL8Hj/rzI+ZHhveS5M5ulAaZeX
yIKgu5fQ1kl3UWKepOoHgWL9o4IGMY8oZwEGMcZkNpvxsstKGpiAPoFiPHNanrO2+6SWtDCgTwc+
JG5j1/hO4+QBFaEokwrFQdgWjIWpPsQ3VG2dpSr0NFxskl8DY7wOR5nAlZ29H3O0htcDxTseYeDP
MH4CV41bGsUcTNQPwflb912ngvajxM5ounRFWW2apHL335/OI+PbkzCTGa2lMKGvys7MJVsRAqnh
/p5DbUycFJIFFijHLLjHkRQ2+v2Cv5hUN/pbdHrfTGqR4PR7PC6Qwy7e7nyPkZ2r7JGAQfvpNoDa
T1wLjKEkefMNAH0Wzh9gpcmzupa+qUK1mpGMaeWpQ3pErpS1HSq5Xjd0BjJZXbDjxqYE4bFXHwov
vbd+HQsS8aQqZD6vFACoCOXSUOWsBXbB+98TNXtAxtluRKRgujg1lXrDT4Bn+08f6jBciNKhJFTF
dsiTe4euVLE8ZphDpwlCSStC1lO2hPjxrFq1YEzd5wvrI5HmyeFFPb5IR+LPb2FB6XpY4Lq+OKQW
NoKadbRDxz3IiyFSlO9SuohFR/QrGCyqwidVEy/26cCg4TmJD32n5tL8OxcrysHlZ7rIlf+tgvUg
pZjw1bLLqyw9DdvkiEeWIn63h6Z2JCi0o4W9MfMkliJgSh05iCqxgvEJgITTzbb12UIReSAXXx+k
HhBw5tJ0y+U+lxBRmB5ZQUMxa5UxdHIomQ0XwsaceYv1VYcp7Jw16SycPOJHOpWLuuXMmWJz0B8t
Dp7xnf/mDhuqYHOE2DFbgMktyvSN8d5iQ99unXkK+SKEKRrVcCeOV0Vpkp/UUcznPW6fCoj4GFFu
npyxuPsP1YXrtlAUQDjVRvPEARMC94U7CbdkSq6LRNTrZl8UvuHQRpbeHNKi5czOqgW0UZ1ITRrr
Wtf03z/TGBzRci+Q0EQFzWxOI+YA53Td38Hu+ZUFONKdHtvk+c3fUqtxYWkmoWSP83FBiHq7JACc
Mrz+mP4eV+bOc+VV7rTXqsjODic3s04dXlUtTr6FfD+oiioqt6f6REIwbNePF7buHHviHMRxv3Wf
mv5RjpB/rPnTSpihesKpcbZc35hH1wLHjolnXMpW8syNL0A0bbSqRw4O5uoCOmKbGTd9Htfnh/Kt
VgZ7u7K1WtCiZFx7ObQon3MRHULHltz1Y6mjYjpftSA2eNpOnuDAFRHgrBoAtLFaEIo9VxlpvWnv
zW4CRMlYH2prQPHWdIEXRdvmsq7ubTJKA4yxvAcb1psYCL+paBBO94jmuxM/4blFsnpYXhJc4+6H
NQ68jJoHqqvnqN1CTsJCczqyxScqyZ4/h5NhUxpBwIsBVTJ/AFpgBNv6ehqGZuNR/JlSgG+7nyXZ
u7+NxXABJ4zk8vpHxE7yGoWKCLfKQQCIYFGK5iv0rTnWQ0TEOmC9SopXPHyVenWr0J6oznAkuSfJ
ne6r+gY9fzumn6DnhzFPPhp+vgJR+vfUsId15HK4Z4YQFT2lVkezqE/r+ZSbsKSDgcQw+jasLlyQ
14g4wZSRKGWGyL08q38veG1cGGcKy9YiFuXccunEnqgwe7qStakDkGckf7tEctyHg5K04UCxdZ5W
rO4wyU1LuoN9CLuj0SidhE5eUGPRYuyAZJUsyiH2wnGpsxfBStQMraA/jMF/W8+57qkuBV/Ur73i
W1gYzZ5aNMADXFLxbqRoUVd0Mnk1t/CP51tPXenIRsWcJtrfaALrQvNN74qLGWbUzRtH1HpHdXKh
YgkkZdxrwPZSpmxdx9/habScG6hTses4pRGMYEycbseZ0YO06uvtWVc1b+pW656kqruly+V7vD6y
lg1R2Rqr+apTWjB2Urnrd3+Cz236CrqvnHfJsbJlmNiL/O0KcGdUuZGzJctyhz66FvHG+akgPujJ
haGy6VeVJ0Q1BzBJv/1MO+sNxf0OidhcHDtGpFcygL3MxJBA4uLu/m7it18jgYBPsWnJSlZQqCdv
Je7PVMH+q5gJFDSZMADl5K/692Gkwzp3b2xAFbzuaDGQC2G0bc9u/nP7AWAfdjYWOLET+PhVfPNP
f9gV281ozYeRaI5UiGQYsFCB/d91815v3O2qD7AtbpOgrDbxPhK7cuifKni9iH7rttkTewT/2vEy
YBl0D0BaJ33nDZMFec2CjbfRV/CpX2NCArUfdQ4B1UdUK5oSmjsGsIW3OXrNBPjW7c6RjLr5SiJa
+AtzrkgmPiMtrNbuVU4UPgyuTa1vBNqgOx2aSi/HiWI9NzD4/OMXiFonLYtuc425KNu4EYcrRLmu
otjHxO0Yy9mGhYD7ww0I56P0cjVrncln8EwApxZJBcNwLnRT1VfbsdIMJLPdVAVnOIVqg1zm+KIa
yUEkOexQdc/eBrM2FxundCrQ/FCMcEzOVV4x/71sxX6g8Pwt053Gxk4ytz58uNeR1/XLIZUbV9jI
g1oSehJOhSZDGk8I4UoZ2rB41yiLwuf9fYX1lNteqyLjH5VKCuG+oEvudJjf09CbrWKIVserNHpy
KgvCMwtNi3HasKpFUiWqtYvbW+9igaKPOdxcwwyfV9ZP6L/a/x7hsXNLub0bE3JRdFitaKVvgviS
LYJFQ07DpGzHkbEUSNlE6kMx/wjT0e2nLSRwpZn6gRB8+GWeiDhaMtG85dUz2NI8pM0nRP+1UbWf
nog99wGQ8z3udcLKO1fTy5pagfHtO4tRQw1ufopjwMe/Z5/3idHS8q5CIvkvJGtq5jfxkbuh/j71
pPT+dQYfVGVHJoBjw/azl6xEmi0m0gfmPCqKqkZvnV5Jo3cknXH2vNeUUPR/pQMvdB8wnSoQzVh5
BJfTworT5uRPOOlJeSa4IH4+e6ysVuNZgvbJH263uK0md9wQbaruwEWs0JyyXGm+pyvtD3jozIly
LRn3gbnAXWUh319HD16Tqe83ZsjhJOI0+s0+F+/L+xc3gnOT+8vSTGSHdP/d5RAbU5uRFYeYRbK4
y9WdSFy6GMniWfWCTiHbfvLX0dFNNt1++a4BJ2DY/Hvrhf83ry3Ed9EnQ/mVopEhhj/RFjxlEW9r
0JuTGerUrP2iuGllA6foJquOMqPDq5c+KY6Fwn9ED6B3dL75XwKO/d8f/tkTofb/HkDr3LjeF5WP
XLXTVpHCb0dx9SlGqlUPGPuXRLuDzDNHnjDXFj9tPyJU6PE9RAyChDsy8y1JIo3gQjOKYXO+i+je
itSHsFhhy7Gxsz3NJqSQyhtZAdyEodZq1lh+P9aRMAfvKllcPvWgBucQgfIra/JIdBP887fZU4qX
sl5Xm0blxcvONZEQ0PHJ3pNkhQ+o8tZcGnQfJLXbVajl2UtCghWAfEYdKdC26R3BDgVxTpxsD7Ao
3vFzaSjjPVd7qEqczQa46mzg0TSp07AQCeisYc390uw+lfiyP9nkuasl1AT4H5q2ZC+Hswa25pt6
cJ9eU05UgeGDBoOx1qquTLVAIPH8M+SKgtVVWi4JDkg0tDLp5aNR0tCr2jmGR+RQLzUrynOLzUVN
zaDLjCTN/GUDGi5KWfL0hjC61xYTcFW/wyLZTwFaKVV1oSMLs7t14M+OsumTK88fQ7fAolojZjGq
fd6NHAo5U/Nefikh54FJeQrvm7sq8ZTCbBonokyt5Z29kuM31kHxB4MNRPrFwQFeQ+hXaZfYUlXS
un7QAwQrO4aMBuO7LAMX2EO/IyI+xPzBO71RX61CE4n6hs0Pjx61yZ3OGKQZUweHh7un8J9e9vBe
l8FvgwyNa+H6qIspeOGzAhMLF2OOO3eBMWTuqcGa52xOmjW+P58rmzYKkwS7sQUo/8ejAcamm9ZA
mVxIsdhjjpftMCaWvpKr+50m8l9hjO0AWCJKCCmrVhp9OAgq0/S9NDLKXl7AvFc6I5GDSD7K3ADl
F7h6n6fq/6jhwWzDz7wmPplodFuq/EIPKEmNo1u/m/aG+ED/q6iRvpvg3a8LgtUTOLgGjOkVmZkM
VMclZ2dg6uMCXEtGu+kGkLqGlcvCgbYf+X99wNz+NY5aLxdQ7DVddQkOGitugzYmii9ofx4iUqH2
60NXhBiRk4bK3zA2iwHPEu2dtXE3+56bKO8HB6R4E6hWe6Ju6sfhOSMkwhZvHoEQ4MWnjD5twWbO
pekrgqss9GGvvgc+hGVxT6ol/kbuaYLnDEaFp0ZHDIpclWCZnAxmK2f4nrXemg03Pm7ibTHQzorp
JbYPNrXhWgLF4lTcWIP+y+3Cd5u9tGIT0r+Bpy+OUsM8WvXxmNO9cThcq9wOMx41Oz1Av5e8Os1n
WhOll6M6LzQjOCkQ4hLM0P58CMhALsQlad+cATIZrPrpb3x3VTC0WmsPr/FIDarFLkLpGQIsnCUD
HxWypN0AJsdzFqLfPCjOj38pnsEGSQhmy0R+PIURtjrw7fS6Fd79cNhmorHTweEnSjJCTaXvmCEO
v1O0wqqMknXgn8JkDJYad8/5lbxxks0j2JSKPhbuIfsW4CUfoqbvRFe9YaTx/V8GioPRZhxS7LVy
vMDKR/02jxwa82F6n6cuOW6kv/O8iRSdMAylFtR4RrP6EtLbLyHYR/pLSdzIa50Tq90uPqmMcgZJ
O5fbNwvXzDf3fHPKSWt1sZ66exDuq1jJYUkgBbixxV9oJeiw8I6kLa/HwLSMoTJC/jD1VcUTyo18
8hOxsBkfZSUwpPhVLuJ/HevyM6b+IKksV441/+bs504ZCu+KnfnVk58qFXK3wokZh9p0REOoXzAe
jIEEHsuhcO2ImjnzgSi9dJCn/ZBMbpzWyTp/c+gJujv/sdSrJq19kd3HkMITshq/4FOYjo0s9eER
MfK+Mf9UwhbaWqkYwJZ2McTy9qyFOYsILmKYgDWaBC/OVXxQ6g+FilvNg1WSnY7qNSa13SYGBiwZ
ebT41ld5q1yMgUdDMNZxA6M3PkxisGKN4YdvbCnpvm6K/P5ONJWqpOH9q83PU9MkmQ7VAilh4sV+
9S0nPRVXs1yDeJLG1ymwRHhGlAgGC+VvV8qPQZvjBu8XxYA3BmCqGS66nIuBB6Ba2DaTsMDC2wmQ
QUvBK/rkcoS61Q+zO5teaNMzMHPjNyLZqPjda8vNlmOLk/vSe5EjG9xCdG/ksFAnRHhRwsvPjIS1
Kw3ZLKLVrvWbIi2uP9J1pLRpZoJpWBv6hVOcnH4iuObkhairbAuYackFB+of/BxJVM68biqdE62R
pHzoIzUQ1ApCA2+BHPGPTaNKu8KB7lqqfQg8OoE2K8ZkT359OOajNjJ6V4VxuXq53apTmho6jRwC
HETAcnjMJzhBIQ3Bs/jcR7b9UUJnhcvQBCzvBQiC0VwYJhU7tshrEWudA7bPl21S9rmBVbqkY0+T
xGYhUHVmOUJswCLF/M9lw50+CUa5B+D/DH2ltWlN41TuqYvx8fs24vLSUwu1aCTmewAIc648l3Or
kEnjvZz/0HZ/V/54wXU8hYKTqTyd96KESEWONsNWkWV7pqzDwnJUco0mYXcQ9YAad67sCYRDtb+r
McKvs1HjFYZOexaw7EXgzqpvD5ToENP9jnfYXjGz2mFWauuLGE3rtMHmlJHR4Ov9QEhs1zwWkaQ5
0HrQAs51ueObSIS1gLADGGuy5HfUp9Paj2Q0CKS/ScqSSr8TfUsKkvnbhzIO/ClscDyrbF2m0gIL
9EjkUgU+kY5Plp1dNfCoQpvitn8lBEkiZoWao8pA97XXxyYO3gqTamhy
`protect end_protected
