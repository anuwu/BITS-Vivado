`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NzvuEx0G5HwsRW6LabE9tv6D7miYm2zk5H6PW0m/i/QjtjDng/QoHKP9dRkjbY33CGdh9buWzj/T
iTEwIfiPpg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uegFRRymlgiluqMREKLn3cmKVsrP+ARyKVAzvWBCZjZFdPGfyfY1J+5BT3DHkkLkddk6wXmHAzrX
ex9/7rPxn+a96Sl0KbXb2fdynfQE4js4WZ4s30akpkF8OkkOgqy23iNrGN18OvdCrTBqFOvQDaql
PF+LonzhjBYxOrtUwws=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gjd1vqFRZ8aTV+TyahY2j1KhfJ593tIUNpKdAVhQ+EIPRnR2KOwC5rRL8piYbMs3haRMFDq/M3IT
/aem+fv27HwFPFJmLaqjvtVRcHzMFp+FoyAcJ2mxiZH9qUywwXzjLPC2Ts3AYHsuVmpURpaacNOm
cFmCLiN+R+wVCW+cs7dE/4hICriINqxB5Kl0o4ROo7XXB8/xYi7xz/etzt2PGPKbrFy/qH2lBU2d
WiZg1a7PxxaMbHGX9OoSkm/vIR1ccWUUzgxhyxc2V5sGkjZMGjZa9ul1SfswjtT572WnNbWtQe+S
lN3rKrYdh6Gwx92X062U5Gybd3T/HBAdBci5XA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
geKqy+6ber8+msEscNCFadd6Y4er7BUAQDjrZkOBYXPalMttTjCT0+XMYDc8PJKznvwRMh6ooDsj
LZdawq+bmAdqcoz5v/4rkkmAhy0/ncLLCypSXP5X9tWWlUoEnvVbtlwfC6NwKkePEGsy7Fmll9Ad
2sL7f410b6I9rE2IjhJIwoRdTu4EOu/DBmpRZqmekQ8pCo7+WwNVxtdxvTIXxS6muy7qQay/fcbh
di2a+gCDWGkGZihCVDg6775vyIidmBIUs4RCZKuDaNMpUYm9/mvn4/V9TEHX+dBB/h/2zp+C9tX9
ynvTIfmzZkBKJ6f9vk6mvrM5IXwnG2qcHTKIdw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dsuUaPzLcdY39SvSBqgPXClrpHS+X1tsCzGy0CVXwJqaWmB43BH2+kL42HsyYbHdRL1d1h2W9PvB
NeliTjJoWFWFvteYzOezxoQPAKCK6SgqxafIETsM3orD5vr18SGtTi/27/T4Y70CI97FZK29oxAA
JItt0oJqYNVIthIcBKWVAEvAm5ETp6YZ8bqYkDu7w9Rc5BGjflKjMZdaIFkCkrvcZZ8pEKx7wlFE
NnHlPu3SR6Kg0jKzfjb8z1TU9bx7LxEY3kORUSjwx8tq2Ba59wVbVpMd2sUfVwCKuzW35pdVhJx/
EJXk4dh40/eC/1Hc+4WQopogb3oGihfV+iXAug==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L+I9JABBUZjbd/CC5epF3i0eyHgklkuFl+d5sHWFIHZaeNgsI+CYpI7zMU0TujxRxfXut/dDvlCU
znUHjYaZoSIxQOknBNW29IlmLFK3vxW1IzTKUT0DFvuI66bCtIhVRMdhW2j7hIggeulPevB2fnaI
YkWXP3KoSbtPRhHzRDk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IBPd62E3V1LjxCYxudvor1B0/8+0308rs3QbnuE1+UsNAPZqssy8vAjEL4xFi8qCeZoOXq9+LlbN
yU9VHjZDJBurvxM4T0rHxh0E5u5mGThlHMCOeTi6+syqAtm721hpkbPDe4TDjU/6M4uKwh0fRCm/
1rV3ZeaSGS9/RoSU7wzUf0kFz/BvgZ0L669JkBQVFeiM/p7ngOhhlXZvPksUVkNTFmoa5U/dV7P1
QmboeZWjz0j6lpYt92ON9/ofUBtpJf6+WuHFpNxXsPjScFxhnbYRXM0w7GUtVfZ2VTDP0EbXwOAk
TlVDgbAqmCGp2OZBUn7nvg3nMIcXVY0axMVNOg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YDu4ql3XCT9RyldgwN4GvJ+W4jcRfHKJgosq8hibl1HWZYq8WL8TKFYqj4JqsEg7atYHTR0Mp3R5
YyCfO/2C9da2AK9U+XFlUv/W/ba2Swm0HZTdSn2DYsfeFh6F7zgHhgjwHpr1DnRqd3bIXcRMVxPm
T7bptSqCjMDJGTaEJhy9JZO1/RuXxA8CbNkrfR9zG2Uysg0p8sg9BRV0Dxc8R5wPj1KHbYs/bCxy
YDjiii9PoM9ERF42RFALedlZy6GwuiTb1zy845keOhwWyzkdC5w2ZuJlgvkTMgB3KU+H+6kvnyxt
B1qfyGwWxzQtacrl1R6XexCXBW+tjYwvdEeDbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71392)
`protect data_block
XaiUK/idXQRSskPNNXxE+6Fx9eqECiI2yJ7CpdyooLZy3qmeycs9anvzb07og8Kze7c5zCZGgeSg
7qXsavC6dbqFfPRRymwQ01Zbncb6KFV3ZUG53jgT4hWhYVdU9UGj/KWtvvNZnz+GC0dk94/xKxjm
zq8v6YqFFvmWWYeJRC9GJkt8UyQSMEI2KO2bek3sXiEPIfZWaKqm5e1r4LkW4EaeMjbrOUa7HbT0
W7tkuwRG/3G2tAGmY+qB6jSpFDFSMlszExTdF/eKypUgUbLABw2mQ+sFccEsJtt72igD7c1UTrpu
jr20VkGOEG43d8CamMSN5fmJbTdv3yvoYklrFn1ZOituUKxK4dhGdQtDssXbwH99fKrXC390dKRa
rm7kYkI3Y2U6juhNZ1nPTag1LUGMdorB8EIFpiMSPTiUei2yfopHU3ZYb1Urng8rsdXVXs4b9srT
GBl+PyuV7/XVKwBVuaF8G0bHeJey0q2kQhLYrU04SzNxchrzXKCEw7lueSXf7g4dkI3vlFgUzE+e
Zb0hvARR8WrywgYOrQ24/jmcHWPpB+jd/4V03b9QWmi+o0B2kmqpNsTp947w9+0fMYbaG5Xov4+j
mqUoAtMELvmkj3SPjSk0p+sEgQWw9xLgI+rUKfDr3XRDBXZ4GioMLZ3r6k8ak4cxn+WMzpdxBD4C
HFnLnWm+RZM86XjjtmyXg92mt6cAtscoCdXknkrhs41qavz+YYcP1OfZX+OiPYefIElN0KfGTHaW
DckpjGTs/44/fMd1rvHc2WU0mcYwnXFhhktXJe/tO/wFwRdxq/hMhmjAvKB0hxb2c7e2TtpmyStC
FZJsBV/j2hG0Kmpl3HvgKufg2ymmdVrSocEQEgDc1jqupqOKyiUYH+87JI5GfFsxiPlzaJiT1l1/
5dy5tfHiJyUn8/v11iGzPYiLv8RIKjTyIWT9WIGk5LaKRa4h6wsaC2iaVd1Qhef+XlaHR4icM7Xr
FJqt+NZZMDfo2S3BbpBBwsg4cPUNAhiYAGiLXOAMMHPdVgIrjrZecXMYBaEg/gbgL0lLY96xcrvI
yqOkvmHpHIJBCYxhu1cOov39k5HtqFmh6MQwH+7uKbIXhQIgnUlneSfkOf2y5bl6QjqYjXEReMkI
vKVgCQaGQyr1p3yiWdJtlp7492cbdSXA5JExJVtEERxHbLVLA72m1QPlBDYLxVgqJJ2cRTwhwEee
lkZL2wzsg670Ua6+NzdsphpE7841nUeN0n31csfuBB/jsHBdtW9POTO+GwwWaugYnfcQV8hNH9yb
WKoG8qTTrdlfO1lwfkmQWksDarPKWqmj3n8uvFBgyTytQwlJolCktBuySTknrXMfRPFF2+WYJD02
alCWr3X7/5AJp0JeI1gS9niPXTgl0HeGsOncgj0UK2RRgzUsdf95id+75RuRqQut5gCksz5j1Z24
LgSJVzP/G8RXKZ2/j/REC3J3JmeHS7IMhlpNGhKSeRUBIIbx1XVbarUOvRNCu+sFxD9D7/lW8RTz
mxG53fwO+Q6EGKb8/MkNgdNIx+LKT2KeYc9enhD6FpfiTyLPKIp6jjTNImRJgHuByrFy2e7FRobg
Rl0QgPoinbBXaKRKJolug+0Z/fT2Y2M6ElSRDkaKTY5/YSDyaPwSYPSvnPw46xvqdhOWrMYfWJsD
cQIct+4k2gdpgECSSMz2jvNosptA2iRD2K1ZPpbooi9RN74JnzBl/Iwf8Rq/juKLdXyVUGX+c9iG
PApZ3H5Wqa+owBjPfhElSmRhwgJx/xmrrMpsIm99e5xcfEVI3/2mD084usSOiY31mzZ/WnU6eL2y
ivlMuTWxAW4DC6YS0Aqba++kCpxZFNd0ubNHFOnT/l3cSQx9XdR907Ts3L1xz2ODhaDVnqC13FXc
Hp1J71sFZBQFgnPo3liXOnm7Ka3laJxbWE/djRxk7EeAzrn5TGhOprAKBShNQJ5vWqNwTHyoGETm
D8vp59bezYl76e6poMrTE5M7bxK7XHyJGNKnBT9Z7g8xcp4HGE2+Q2HecyU7eYemfw5zQw/Cn8Zo
XcjwER+AoTuFf5RhQf40wji0bghoeQcfsUkw0RdFMCKI4mtfe83/LauXsPZvAsBoTKVQmvP36GcM
dVYmNgAWsq+Khb6gcE89O0/1ZQwCIjHvsm33hMX+oRUzJjiTZt0Hv2oakdTor+bwPpepNmI7Incu
A/NIojChByZFl1TEaCTz2LjZ+wyihnGyQOwBm9JIXaVgU07QcE6D6Ubn+tEkxSc7lO5dnSzmQ+0A
r1MkXySTht6xVuHQVuzD1gHXJnXFgMvBIVWja+ygsUb1iLN+m5IAyYUxruSx1boz4k7M332T3QQM
ZPQgyzjxaTZVxMqzCnuuYz9IGYzpanlGE6fq0xYN8IrwMU+oTQKbzj1n73PG+DK9Jvo8L5sTZzWr
MTt1z8NKZSgAbmXXXArbJ8Exk+hOrMKGX9Ti3Jlmt9pXe+lq5um6tzXQ+/VPeX31hgKLBZKK5KMX
DAz4y+6/jbvK2fRxTTiR9uWAsdW5LQ12MwB0qu4yCDCs627GBYPaS2Nd1+knIfUi8ROpNw68OtEU
GvbleuZA08KWQckPjTaY4jnzRH1Z5juK8RtVCRsvI3xZZJ3N/0yUF2/gZN/ro1NJGASylaoA1d6F
kBIlzLGu17arPN7vEDY21dEznlbGvqblvh6GSPguMgoXDd2tRYD0b2jOk7i4ovYs9NJRDv3DjkQ3
3Z+B0yS0adkaoIKHbrSiD+I5idLDYc4NSYtx75WQEOd6Xyc2UyoK9ZY3wzf7gLj5wTxw/YsfLdQM
lyyfo9btNX2vEbyM4aRmqgkyA5Rw1/UC8I9io+iDTKeyV+joJpMBycBk6XfXv0KwO8aGIw7sIgbh
5AT9YNm/KfIGzJiItnAv0gpr9RscBJLPXC2HDsSHN9G8qsUNLy2mb+Xr+jovS2ky7+yz13eFsWHm
Xp6wYDfiTMxizrFi2VZi4siU+ib5qEI6VHFCkeWMf9BaM9H/kftLAb7t3ruwTFi49flhLObgDkak
TjMqmnC5n+RGA3yDNmWpxxm3kijVgLanEvw+axoA0Aw2e+2VRymmPSfxNRS+TxQRp8NQA2Ck0hVz
E9PJ3xZC3cjFJLr4ZvnVBDsIqSjQxhCbbzkbWHzl6zUlv90c6WRVjPgB5mXTUQpIgy2iasmTMeHy
4u+9XOtRoM1JGclhSJnKGPV/GWSky0S1Mi6YYC0ZVtgLrjlXEb8W3IxI/T8hHIg3SG6OBZYpek9l
R0c/3szeDeET5QJFUP0X+QC78Kqg1oB9TVFvyRH2PA/CFA0jIZC1v4X+a+CkdU7ANFZzAd434tjF
N2O/N8J3vd7sA5GhqFgng0N7+fxNdfT0U/F5GsI6Uk+nfEZ1CwRKfP+AbpC3Y+F0R6BKQOHo2Cn3
o/+PNtl5ntaugQV+kv77943KF5Fvxj/RwQZt24FNeCW7YQRkGpNJlDlIhz01AuVWvSVNpLFMgc7r
2KIlsBAqyB2cU4P1MC42vIfwQMuVDMfgJ45tzR8FenMUZ3Yq41J+K+Q5p6a6cjJehCNscoiKv1m3
3HtuAGi3WQBy7QjQmOHv2+e3DqyCu40a7L3hJRPMVvUw5/pBVQoZX+0YEYdstF5iEbKDqLKpWh5K
uuGbn6WPlXDPaVL1drpBWX/J7hJFAmO2dEf1W3QZQyi/fzWXScgEeifqDlIolBBQyq88PEl+Q7LX
y6SNbVneBvU7vQHoszHblT6yVel+V3MhcJ/GDXbwQgVx6hwenqJ7mwKVgaa6BauijXzC0h2Fbb4p
LuIpCUIljBOzASOUrabKzS9aWXFHWvWCBw5JqyVjt96PD+DlQdoGPvdkgcDKy2saM6E5Tu4PY3y2
lttsDV5sovx9WsAcA2bupNhq3Gc6MjAvkJgYQnERNvx8w0kHdoWphlrffx4x719FdNeIJi4k7IAN
eCjbUxndCJyeXrrewe+eKWR8xuyZMQU2KX7AngGHMLUjSIUdByo4LsdB/t37vrlk1QOfo8XOexeh
PBv5+ILGH3vY1kkNOnWkIqYF1a915fk9aSazuRyOZUeDl/0OaOy3DpZ99BCMtIxa0qAWT4YR5+gp
tx9adDgkrRBMJcfKPm1L3rLw/lJRnAP4bkWv+IOYXpIb5TpnwXjBlxtpzDT3vPPsS7EehAwSW+xu
3nUThhfdD/4u0L4GnYhWj42sVRSFNflyGTJJFTIyUgmKCDElb15EkOPQZbQyOwitHF7k3ntPyV3u
XJURxocJtIouJ1KODJKVvkXdC8b2s8/BPr5cUUF4El5i7jctYUKn87+ouhcSsWwouWgM/BrqC7DT
judzC+Voc0SuTyDomY4OP+sOp4SEpe7vcT1XxtFVylWup+AUm2bV9pzphzS8YGdaElYAoIHoujoz
Pmjqf2VycCwoBI3cWOk8AUgJF9vTUIvBxYaFJD6zvNet2om7sFSAdatMYhfIjsnWeW0EryxOrnRE
urETZO7Rpj9ROOOkxLEV/7O20jHoAUhDfhP5Lse2Talz/7WNf4ccqBvzwuEqTG9Z4ttqJtw+11XQ
H8tv19YJ2yGOz3DdQI8q5MotzpLJYilPDHHcv81hR2mN571pkFW8wq0cWlTYkc3h6mUXotpB+wda
RoX2FllLr63kyhgXwgDI4PGUk2uJZ/i4QmnnKXzOXQV7b+S163UiMFgjL/nk9K/AExPk1Dg3qy8v
gGAKIyYYSoYwgDmhD9A3XiyHU1gDWu7KWz83pxbHcsZZUk8A92gUg0Pevp+DtsBhrxu1QL+GmNwp
3+SnZhQ9no8ezjX+9jL2Ve9pys5Z2L4Pa7RZpCjs7Oj5RcRE9WLcWVtWfcoI/kANjKA85YqyMQ9T
gduTPH3wtxGZWS13iVSexyQJxqt4NsN48GtXMX/Z0kFwB4JVJLVgYUj9qTYEwQwvBCBZtjZzQK7i
PFwmfgz6L+oIWYIosvnO0qlsY+Wk049MYed1ZLhqD8Ng0gQT1pyHVeDQpGR3vyWSQCZsLGcMwErW
H2Jz0/Y2sMALaJPFT4DOxoytQk+uuuAxQipj31+ffE4YE2f447t0cfmtOJTXNPaC9LiAMAbq65dg
+b01mumT1y4oS6Zvot3ZHxjUPbPZzdYRNyvCoCSint5VayqJmyFoNi2AwzO6lwIcIJdWriDjzmMz
hs2FkINlke6FJCYi86DktXrsCb5F4ElxBmm+jvGygZG5RSAzIB5SnCC8+4YKtzhDAWGvzEEeluqw
phubSGwCwAucwJ05qNqkPfUPkwlEblvuLnzJX6a+xfLhUuQnHONIdEsabcf9FtB/gu0+2Unpcg1k
jUxytvIqeXoGtKCS8D0i8bGVzc6YLwwagQOsbCGWCOg2pqxb2KqZMiS2hZFObRto5X1OwpzSzwoa
al0cR4Bg1zTjnf3e08lo/ixqSTswFV1fZ4WSSuVHgwsozzGk0cIX/GEJE6iZDaN2kfKElhT4qtPe
lkBY92wS5utX7eVe0OMxlnoPOtL1IVFHTwPBNWovZibv1kCGxhWD6qttlLUlpBEJ0bVZvKAV8ySd
lj3W7KTWa5Y9QxT+jXABgcnUMEP48FEUvNVbN2F8xj2PfXUcKaknespQW12EpCk/oNrkL/PEz6mF
j/CXgAEEOHc/0RK7yOobZx4cEixibP+QED0FMMmOKKjFRhGvs1jrEgKQxTZDA5XUtR5a045y9Kok
ufgkvduPKPhOdpmOJwi85aEOUe7fi6XXaKPLHquY8bXYlaCo+OWdD/6SvchZOJzO/e6OIomiMMp9
Y0kgkRMPKBpfcIY03A1ppkKhLo/DNmB7MCb759RR0qoICdORPSPNIw1YGnWhU4gu59Xhi+v2Gpzt
kWKRQR6M0krLqUZIFmKaPyC0CrjJAimlg9Xd5iFCXfDCKn0f2qCmkLo1jzE0Snpff/Dx5zfskcwt
smYi6GNYecw2330vl4f9dBIgyx5yHa6okfz+Oo8Mz8CrJP11NxoCLNLf0ak9BwC4EEJZGVBt5x2t
7ALnE3ILSUzOtqi4XJx9QLsozRaDqWkOSlW8nXVWWOV3DJYQXicCPol7DLwNYPmsX2D3PS/JEfrI
0QoNE9ph3oeMySDn/sz0laCIvdqBOWBR7rqD+08Crntn33bEVjNNYRCXpW1uaV3J/xBnqtPdzDQH
H0OoJr6Ihw+XvHmM/1K69NDNFESK0OCSawOyzgeypyvpqAnbA+PUa0lSrLaiwiWZo9R4fRWLnvkt
tUeWYu+vf4b/3JGe6CcIzMliauiuyiAkup0mCiiuePSRgOaat1epvSa95MP83qP41pCBgaplxIUN
+ISqwnShRk56HD7Nl3ti9bEM+TxdBwalf2dCiJwrQV+S0siHxwBDkx7zVbWG8WckoHyCDEScsMKS
xjyzgj9NHdqqbAoEvW01xjlr6HA8AqxQRlHlttfTenU8lOl1JzcKA9zhRyGVzChfDRNrGeEIQ1B0
jHc0sZNNOmORxbqGD7EByGWlmGdpi30deh79SqgEwJyq7uQ0y/TRRNCciivWEty6cyS2T7VjfDT/
idN/4SoaXNk4eXB7anE+riWGwjJiRE4ZUWTb5YVM/o3wLP9r3Oic9KRIS3WhqhGe7mapLqWNzk6z
5vXgx9MlLjx61YQxz6Ke8v8Sricmd4k/au0vhIVKkNj1KfaGh0j0ER2YjwBVJ/eIVACdoFLSrYod
61jPAlobG2biZWEkGvp+B2UNfhLyqFFIOttwWTU1cG/dsF0zjXimJGlvNKzv3dLr8BsDCQNREYLg
AcvJ35hF6O6RTLv16aC3DhNM334AJdvL+8WTVDrEm/mEvRPM3Dl/gFp4oOJa46eoLVFTxe/iPJms
YRT/BOnyK8zHiUPUqYsLJ4c4hagK4Q6hX6/OA994Cts4Q5HreptKRevyr/KzDvg5GvhaK98KMeuj
kDT1t79EQYXZQY1U4hQXQl3eWV2vwKGfKlmXOEETVR3EwOM9z+m0SpObC2r4eq5qtjj5vsPyMXRr
74JpghiLuSZ+CJoJ/apiMCumXd8DgKzH/047lid5LvJbCFf9zWnQ6bN5sXaBZB5h6acX/sWj/kl5
vjmxfSgVP5ydkiLzUDP4JOPZyaIlJvmtu+y9SM/OwI1K8iH82AS602dvWo7OdSau+6HRrxOIK4X+
mvKnUwkyui3zL6UPfdcyzwCiAU6px3JmsQgbLlW6u7b1vB35SQdzu6Bfyye8u5nPSWh/RklqABEW
MeE9BOPPhmPLqlADYDAIyYg7D1FkfeEXlPJXv6D3XeirNJ3MTFY2HOodrGfecJaH9VXVAGhZkzd8
MIW2QiZfbHLktwHaoY5mtDRU1YqduEobMIrFSnCvlnrnTXb6M2xSwv3g8NZPH9HH9N9p0RTCcUH9
vtndcwzUAyQbwLZ6dsPbQvX0FadVLX/kOH+QgXrJhAbfq4arm7MO144KWsOlgKn2DHLzs7K7/c+N
gH3a9+K67i1uQAgUtarak8LSENxnTXsqBiFwRjGotOpkPE6naqOIo0N7n3Twu6ZPxpSpGYFMJK64
mmRc+RQVn/UqTjI7UIeAhTU2S2X+jk4omn5+wb/NPpiNQih+LXdlSDLbrHFMimWgcGpcU9tokV6f
PR960KSJHmNfSwLYln78bX9ldln4eQEKW+UsSZz2uMhuKLU8YOTZ983B7VrcF9E9bZCgwv0U8kCW
ggo+POIjlysgCDCxRV2LQupyc+HxBQ+eXx/NI6ylWxqDcxtT+Ai4M35PXfc/xvL2vtBIV1opBDwE
DSWrytCoLeFGv/0un4xMvE9dI38D8XASmx0MZQmZldRxp+u/GL2Fc+E3XOA3LjwSbzk/db3T+40Q
o8Zh0nlenVJYYwTleYIXmVE0jbdf3Cx+yFybclpbMOmlpifICf63x4qmz+p89o0cCerS5u/8ql39
hkAJobldDn0SifvTBk5fkdJeOv/PPnRUXb8Xa50EPzkh9ITJ7bSaHQc/LPr5sZxmviXJ6FtLbk8k
bvoR7igVajk6xydOdM13nMnvhF/jqcAfxbnnKi7qB2DyJLOonrPuR10b16eMsBXPH/vmJEF8WWXA
zzODxMBbGBOQWuVK9tNQ4NHTnOJECsCbXU/PcndW9N/yMBeQdoicem409aG/RJGsVFzai4PckAzh
FwCsCZ4nkzuixh4bxIaqg4mz7cR0nx4E2ajqtyycqsFv0G9RIJwdUzE/Gb6zyLcuZhepoo+FH1EL
B93UDKnOjpiV7cetWu5c5frj8u6kk92q3jSNQhDz1RzKiSu+G1uAMnSiupIQYr5FpunLBJmHFv1j
IQXyxEikmgrL4N5UiabXzGrMguz0jYDcWXbp9dN8ZGJM627gyOtn74Cj9bD8NMIyWdAUSS6uR5Cc
PJEwkxDjkCHLWuA1r1kLyUMAq9yLwf0ldFkyQeJTcY1WCu8fqt4Ih7cFM3JHlOIY8p5aM2DAUdWo
vpPc7ZenZf8k6DPNtyuxKE20MUw8ANmNeSViwB5ljTa2j8rh0Q61yRjSdg71Ii0e85r+kbzyNJFW
+MJH5p+BCbCT/7Z+6Z6ruuo66D2ZAtgeAXlQLKJL7dSmJ21MgnFnRXLOKcD1VBLjP4cQKbNz/vMv
AZZ4oWKHvAJfE1A3ROL6BpwiTUkLUNzk5Hq5eMPBnD0gyTJWCWwCXcvPJQrvLXgb6yKexYzllxsy
tVB7vfIXCItb4BGBS1+3D7/0c07aOvWzDKV+MM8qgIajN6VR822ihLfPT2AD0lerhzEw6i/wsF65
iOG+ZLJwfF27efIFE00imQ75+CQ8kRqVjbnAl55JbIPPirYP8ImL4qC6ySz4UMGD3xWomiyMF4aC
bmefZBGS/nfe3vdLbejsEG0z/UlwHS+65V/OcKdBu4Il4GymObw/WqNeabJ9zpWo6AktCOjztaOH
nDGQAjmY+d9kJJZ/QndNPfUpXdTF4rDs1Y5Tsxt64g25UFK0mY8jF4ORcvjAIdu3zXJEUwiRQPut
Ysixbz0lVm/OyUt5jwfyoslcduUYS7TndrFv6kaAJvMIotDuYl3U/y1Qonttc22j+Rkgh3oI3Qfk
I6AyEieiPxqiUlpf7mbQrMDWtoPZua45NBztpeV0+XsgWztNgYPxgdhRfyLb/O/ZqBuoID7fs66C
eXYwbdNkoCGuCbcJOlqes7LnWGIJc+Gd+8Vvr5iZxVSYGaAfBqazFZu21B890Nj8yDQqhflUUGpE
pbEXk/G0d3pMN7ufuBzy/jEXM1oNuUGKyrxQKEVAMFMMQZMNLhJL+J8KEvVRySNS27MUonT8kX1f
5/57kitXQ9a/12rp6mBxrgi0NkG9+WyhVyGVrLfzxeiUMdAtsUSnvHgcInQMsfrZQSmIh2bqprP1
tAdC/sPYCZS6BrQyY8u52uiu3b8yU3BXsRgDgv5bNhBJayVnwELnsFxBgc+eqyqKSIdjxHwG2mE1
uqrJYbvY2LcTRLiAw+sRGN/qiRujSNNExnCQeTfbSt7KuDHUyt747FgFN63TUQmKhG5C+oRgjRTs
ab0tHmUxIMZ3NppLbtLruAg6Nn/k4L4i1sWk74J70XE0dVYvfmbwFRhRCef3Tz3Knkt/H4VqAzje
euX2ELBP9jVHtDqf4PlchpJ/zzUggnmF0qf3CdMD8NLelP79/KAvZoCqvLpZO7wSgHGav3j/dtGa
V8xGBqN27vPhkH8tD5bRCwyECk2ZGjEAse/KXgvFy78NywuJk2uPAc1RtvtkR2Uxd9qsA9ileZgI
OHXJ3vYqTV0fPgorIHV7sJ3Wz3OxkGwYskV4+mCDmsau/e1nNjxQ9Dj6v21rCiZp4CiNz6UPAN0B
4nCyIdNlzO1Da7RcDABhTyeb4Xw5uP/wWfwrvdb+Eiovj1gdtEDPuo30t0OLVnG+qL19pW0Q5BeC
lih3vsGxMMrv/CL3GHmwU3qU3jgWyGOdfIM7Ple5SV2klJNoXovhDjpSCnJ5s8RAdqpWDj4ElpMO
s6hTn1nxcLemx3BKAd2mxzEeVO9Zf3ah8OVMJREiUxyVeknLHhQ26HVvD9HDM5aMcRjzQSJ0evMr
e6C/cWsQGS7ufwY8pxQ+rzNXWolQiAWH4DCy8Oa/VuvFJkCEuTFjOyy+qlwa3dcmUu0636X4RNYu
sRArXDcjSQyFTo33yPSgtpVBQASumr1qh7X3A06Kx+VyAR9Z9bhvf4KJLWTKvZgXZtClPH1Ms7Qn
ngRwJ068BQHPG6v94sgg7p/uQzJVvowXPSgzLCwgHMxo/BhaiUnl7ky7CDxxL2jjCiqOAWHaSXUL
PTpNA/L+wrsXVyizaT84o+Tn/M/gdqlikN+eifCkb0s2ADDP0ai4Ke9MK5kDUG17WbvLgPW74bQ+
ivKhJv+9X2NW2cPHKo9xCLg/jndBtHtR3S6L6A3CQtPLRlBkG5Te3lLk7AJfUzFiyWgMDmgVF6JG
niBZT4PbsYRLFYmvM/rpj4a4ZNKNccgUwTMJO99CBLS/NB8z1vXR6kchakpvWcVJQF95+eOOlMVI
GY4FodQvSlssdnreGrURnzXOUX/2Tc4a5TASGJU+r9oTJtD3NMl7/LWqmEsHjJOxTByIFpV6VbCj
aU5eDqOstwCXSt73Gz4ZJR53qwsa59PCKhu2p0QE37hE2x3YrSDbaVUJbJvaqArTUR5YX9uhxENB
4QFyvNlOeAByzq5ZaWyr2rmN5jM2gzNKxRmDi9VPx2/dXFxsjFZMvyrJNI0p1Wgkb5B6wZ4pjzKo
lEz/6QmbgWZlr5KM7dyaNpNiPuIlLkT5ffTgbXRdRsOyodcnc2IqsemTF5oP4wx6g5RiNSXEQCYx
6L/8HnvWWVYuKrTbqOMNm8B4+0ss9lV/Y8KVGk4hxwSlsIynlhl5NRsk2V3acLTVI/9e8WioqlAQ
Nf/Pu2wYndNe6/TuiI8/Z/NW/fSMDCBxVYWy8DYtf+NhK5eiZ1c+mRAgdc8EUKBUaNslS9fk1TTm
dALFAH2SKugNEPDUfDqfmRHxGcmVvRoBc68DGFLNu7q2xnrZKLR+gvJ8GASvW4TTxf9o9/0r/s0s
aWKuniBbsi93Q3Zy8Ls69ErP9qo2wloheeLXndPU4NKz8a6Y8opUEPuUCxIuCL3h4h6lJEKlCB8O
3drruZjKAEWIZHS08Z5z1c+LfkdtlDGggUTdqiGsaT//pexrQ6wwS2+1wxZ6vygeBdvF6PYir0NS
1rOqWfrhh6BmJi2D3UwIpiWCVEnkBufRwwdCpvx5fdJy0uZay4ilPsgkhzOsmjYtg6EJTCReFBfx
GLWANBpQHcu94xbmB0ufdTvb7oX6iwa6hLKvJhXxVPHOTfbhRG1l/9DWe8lPIjQ7cMvzSUIuTs3V
5EQMOKHfUkq/XZBOgwbIdvxB9HmS3PLqaUt9zZrEjgrFb9NdwunJmk+egLyU61nV5OFaUDOauoTm
4GcmeHdOgiedixfmZkuaWtlrQ+IbAo+s0qXEgNMCqUBA7wLe+qO5f1OvJKWLU3GAO4xhwwmHO5AP
47D+qlFigYHRRAJXvFSm6pNsvEyD/p0MnCjar6isczyCUrT2U7TxgsHRHFoN/r1gwxQ3XqzDIBqX
ZpuH/bSkgG8blmOqpEqablhUx3cIKxlBs7ZNT0cKnZb9thYgWOsdjvB+8KrdfU307Q9mZ5qSiY2g
hOKgpfBHTFADJLWojbYZdWTr+FsQBbjYmhz+gjaX3o9+sYV2/GtKN+tedDdcuf9l+LCyYaS2Byyu
BaS2Y8C7cQcTnQTezB0CR7a2IfrObSI17cQUospkkMO0GWm5x/p/nvWCkqOkCNZYH8xxVW2HeW7e
BZG5MAQUxT+Ni2weV+8M6kQi7I1RZq/wQMceqkyBPBS0efZB3/Nr+w2nH8xne4nzpLLFjVVHEzLa
E+GLmXpY/g+YdjAFRu7+rNdsgI12uItcgWurU973MlIM+/uZvfC8QIIinHJOWzRyjRL94fpS7olQ
EqWY6Ln2EuuO114UeWa/q57eIK6Lry2tAJo1VMxwACeySRRclhOrkTZs/mKM42LjEohltdZk5cLm
jYMqWv/7310T294/x92QMtf9kk8AoHDEKTuJezKS7k0EG6DzK/PWdV0Gtk2l9PMmqmSpCmoibC3T
NJowRxjYNNDnJA+BTGuphdWxVdKTMyhnbLpq2urBYb2GhetpU4ejZUsQFPg0vv1+O8rJieKwaO11
kUnl7M7geApBSKHWn9dKnL91AjPYCrgNC30nfbjpARS7i/WCjvU0bw+H7H9pnPvu91A5Xp9SRgpp
dHLpShDfTHQwihf/oI1nrzUZZItBZi05vKHSUnUxZ3Ef4pfgpjdke3nubaJqG5K8xB7hNhzy1fwm
+PPeXtrHE+Q3RzzcCFoqffg03KbYF/YZsnYc8echE7flTmtuCIMcThBUNN6d0F5AYcz2veEA2lGt
QIXrg0QZnuXkrg5Aw90FLZQ2/BYgbOkj3Kz1KNQG735lA4IMAZ8x15ssElLPOlg/Ax9zXILwoCW7
XN6uKorE1JuoslLbBNtoyrAiY8MFZPJj6NwGxutrFU/POtQv3kef/eomVdnxt7XklU9RheuPtO/W
+WLqPd+TqmE6hA+iEoDrq/L35sOKNuib2XqAWQfJbwidWfgKhacLU84sVdQc40YOTUQgv/fqHJ1x
Dzml0oUUGzZ8n+gGnoXNTwuDZM/uwzzWehak/B27c+vWlZhUiXld2Dm24ct0g+NpVNJE7PKN0nry
V2zGXtWOjeDW6dl71K0QOwHVXT5GPOLejCJzVhV61ZT38pBToeiKBmzex2UJtORcW4+gPGMtM4Fn
CwHkSvpo/+cD6RYVrpCuVrQOWGanW/EWA3akxqEQYtDJopPmFnFC/6ZIFSqRFIZ4uFgLWEZKz8k3
WIbJFo0tktWMqgftrLeUvSIYn79Foz6DSUpxLzZcLcjpeBeJWkYqPZ9RP9Cci/lRBhW3JQ+/bKhe
rq00hpmz6zgLEIK8MoZI2bwFzYEBM/TlfDudml8rrn5IM2nS1psc23dTbdmxVUw1dT6G0VZ4kXrU
DkNdcw9zgBTFdvAM16AT3T5iA871DdJITZWslxWr1yoUxPfb9TgAyuvd/WgdjnG/YdDw1fs/fCsZ
UkQi/nGwlHaIYzlBO3/FE1pUapwLTAiD4BfNwaDsAmrgeJuK76MTCFoUtTK7+MitFZL+S6Yf/CzE
EEX+ftY1MlDEGI9fL+gFhWETF9LqMArP9owina4SY2uF8+Mabnv698gC4pRRcArrYeBGoGqDTzgR
4lqyliXH/geZ5vVowGoVwfAJZFrhgDU6kj3XyNLmK8ktZ5VFaEkfiA9//nhajqntzi/Koo6+pIKd
pVizgvwJCakyupK2avQTXnimADdR1mhvgDSaX0mQ+HbIwc324GhVUMy2jEY7vH2iTdaALTOH0vIx
1cRRhUvBgZzOjqqUJojlwlJx3pd0LE9M1yunckea0V3DViPlJnds14glxpThV3UTRbNSAoYQdZbC
Xha7L94nw8v+HSUzC8JlcmUgv2qTd5fZ/n1tEUtOIKzWaBt/lW9qQmygpBQ+f/z3nG0VfXDI3MuY
o8sbqTJF2FVHEHkEcae2imgYxfpyXL5kBw13neUz9RpRO5VjDUpgHJEo9kKPH9yK16dgosQsLgam
op1KZKMXDu6dAp8dMDMSdLzpzBNc1IkIdQBO50nRDARkQFZbOCia7y+uE439du/VbCuHdy4LW84Z
iiD0gKK3dKe9Trux/pkQQXTU0qYtTsLBoR7jzQDuVyYXWkKPLqzUKugGuuAoEsqQlOBvG99i7Fm3
HOBFwgxlgGs+kmf4SXV8wacVzPeNUNuzt+jr6phgs3bTbQvb2P59OBCDahJ7rrIxIu6oj3cJC6GB
11wLENKpXOsYNa5Y81AF3LLLWdnOJ2ilTYPfRQCr5qlAFY09lYU46kHcLsUGziB5Q2IMqVclhtlm
4Q/AVVcwRqlNlKrrlszeasWgvZH5j1bO/hv+63jLvCt1ZqBneGW4S/xgTHsDKrnLoTmn9TZItlOc
dlrovkyKm50/WvRdXOxlO0jEe7Vi7JQd3mbOhH+f32E8RpQ6oj5dO1/oh7vXXAaB7lUu2zQr1sSl
uQ0ODRykykGg/8zjFnM/NTYv18yjPZY9meJQTj44fsnd5XBpdsm/rvu52bQieUsGnupEQHS2WZXO
L5VxDKq1J8/wLNc26ig6kac17H/AClo8COIEMoPVOCyuIrk8w37ngmPQAuuD+AiYHGh4t97KF2xm
IhaWHrE0Io9lZKh/ywK/FnPYIiNLRHXwFh5NLMvbF+Jls/uzdcRe3Xsbo6Mt0uVAz3y+ssdFgfv2
nUc3qhENPAjW2uteoY/0MgLXBwPj7u31sif9L5IHuqudeiFTBw/8mHwX4tF+pDLGLVo/Le084n3n
REj/tRTG2NFAndEjHsc7ZIWAktu9XtYFWuM+82kTW7QKgmcbvtCJA5kmF83En5tVa3W+TeWEeN5H
8x2ZJZsnINcOVIvgitZOdJm6AFhFKlgOxRO/bkdbf5MS70/2zaNLEYLhHU9OhZxjVXFDJUiwZrHn
TChUlR0nMjDFdsr4QNwhjSW9K5dzaYQvtB1l48kAVluJOIsRX0kv2+gqZKj9bsCTSlWqrJhopXnC
Rj4VpqXiKn9ohHIo7F3yodLsyLeJBSOQemBZ5axPufRgicOCDi4pUZgMy+28EOoRQvtJMGhY3ADR
hl2BJ1Hd4CTAiqkhlvs0Ql1TMBce5VgPYyhM0UQB43JOQlneUb80dJjALxoYG66lz9NHYA0BgXjs
/gU5eSIci3k7uB+nzsdE6iWs7XrQh14/geqfppCRm6aLQ8LQzGA11tCh9L+oU/7+sk4vUb3hhEr0
XkX4t9hlCHSIB6JoPDbqZY8TcI8nHLAVa5MIvKX0CphrHPbHTO1HVB2lbYvD2pZVjYH08A5IbeWM
Uocqb5+WlzmoVPiCsTdxvvZ1BifJeuFZfyemPqdWJcoOd13Lrz2+0Fk6+T2RgSeyfzJYkQk/KUfh
immYZ4XBZ65lsS+yi31bMWkX/H17WHV8N6si+wfmYRlEOoruTfqHhvFTM5qlXaq/YNnxweLe00Jk
gRNyFEh0OXONR3fl5fiodqgYOFQSStSTmaMURcF0vv0nRBefCnFabYKusw3qwJTbt0VO2H+KB/z7
j/RPb5Cx7dMOed2K7HT9nQBM4SL2uq/fV7JceqSdnTCmUf+k9vUkI0eLPYldfMqm3gPS4xr/6WZ6
jv9oeg3UiIbAMEHCCVyIKtIP6vAzJzJnZpLoJkiGPioJs0E0UX7Ls53d5ZYnk/HG500+ofNxBOeB
gBT3U7ho5syqDsHYMrNIs11jMIPzfSfZQkcx6gIlRsU85jVoPdDTddZo5mTaaVgK/LuIYzCWt68k
m6TJfVq3JPgeSRREiTH5f9GS/d11IMT+azl0JGQnJZPcho0PfeqO6YJbvxU8IiGPLPN/HmfS7ixo
bLeFl9uij2k0lMWxZujaYbq/ARP9OjC6gxxcFI0U8fOFDK4kjeikrnp6Ch/Bwz3Sc9LJ04rKdKd4
m2o1KLctsJwPPByDEtt/9e2uBzeXeWZPhiAXhvNcBbPhvMZsXbXOk2IdN2Ux5cosndDtFXY64vQe
j4/jB1J9s6GcwHHbaTFFiMyWSYFpZ5FZO92AHMMTuv752CwKaEKrz9moTVgqOGl1t/ZtVxHUikeN
RIyRAiRWBTZqRqNy2ygxewhqfFeSKeDcJLoZa5cOaxn5DCfCiIw+KXrS1N426bFERieODR4y3XJ4
6bdN0OppodVgOpSSc1BwOBpNx+Us3fPTOrpMxm2MqzWB1oCs+J4+2PYh6IvDdsJ5HNV6583SQ6x4
TO4+Fd6FW+ty2Uoc6jYZk5FlFkAwaaTzdoLyjSmHf5Oz1ORdHOmejiJ2REwC6FvnG109/1sLjpAQ
W+DLp5fGl5WHLbHzRTvd80JTLTurXbrgBYlBxwF9EIOb4eK+9UAagmDHz/4GOcg0Uydi3bgg/Pnw
yG381nsoNHXMmSLSw6JpmjvLrCuykzDvKem6pPDTuJ50NfVAi3U3lUTG88/qXJu34V/MHnlvus4d
h7ZoMYOUAPQO/9fTDaWP1mtBKKuQ8+s1AC2iPh1PtgE0Ca9nCS048QvmNrmmvEGyD4JwbOnJ1Qhs
JxkX9t7raYXCKZto1wmIYwlRyu6I7yNXwj0wVrgFMwtsIT+Ng+5zZ7QyTmTNxxd4staj+kfpAMGz
LWi2UBFw/J22qZErh+R4Uv7LZJk4hWkHkiyKF0TJYyL0JY1aEBv7Lhp+nRARI3mlkiCNthrnq8/E
tzI8Y4NDUqIfLY9hCgjuk8hCzgsfN/rIYBHUcLnjY/A0O8TCJEXAEvpqs/fixRP1OK0bcpHGjH/n
+uGRNsVFcrFzKYcAESGDjppsz/5n7aJz8OXKCCedPo2SnD6KIb2yi7bVIxNexk6LCbfsTziwbYCa
1LENn/28wnEpbGkHmesp4eiTKlrCk/avEbnKqOCgADmxvirWhJWuXd8o7O2XUoR3X8EKZoWlScPe
135bHFqagsZobusuiE6n/ztrjQrSxrd0mopMTJdo3StUlZeIIjr4hRHTWbL/HgECkaPuLsXrvHPh
UviikW4LOHpcLNw7lRXvuWg86R/DGouMebSqrfUKENsChhbWoz1g/YipDLAFmdDipCian8VQWFmk
+Kn5gw4PO6BashRCDutt2d5d96B1H7Og/U6Pw3BAv4drE/KJJtpbPpNj5R3x1RmYTFfmMsTU+sKu
uZ+iXwcTHB+Phy4DVuc2XD0wuqgjfckZBnPRRdjVU9kr+VfhhRaSUGOYwkQObrI/j4u353dvw+vf
hSEVskcEKhnNv9yzzg3pX8vhM0HLM3rYyg7fB06V/DyHSraQqhfuRNKBChUnQ157KhJvDM7Q9B11
Sxvfza722cCApiRxa1eUjmF4NFYLgSLq4xj9lhZAU3hwr7Vbpxrw/zpOWxICNfibE4vnb5H19ZLJ
DH9JIkp63ERILBLYcbyJTVcA+8eDK+b9j/XRFxQz/A8n9MPoCPo4tK/V4lZKF88kmKcke1WueuR8
msT81SjEvfEfgbEzbFxovU6LWaek61trYnnv1yOpb+PI0T83zGZms89xuLwnUOsJ+PBGuxLUYVM3
i47ZG+ROaoef66FCwRfwiZIDkayKNrxITISWwlH7EWaaJYJGIFCD9o6JdRmOQ712JOHJtgwgM28d
voIOd7isMpQKWvHQlz/39cU2VMJK3KQJcec21Ga7XpnqllMBb3xoadBcgQzTi+sV9aJRo5MKkxFe
r69NEONKvBkmwhMwbFa2t15dncadLv8XDC2Mk9W+qr5pAWdd9EVbkKcyNZP1letH9MRIwtoDy+zF
EIsQ95YrlQwfbnX8TEOMYSgp2BfgQe89ER7mLlte05cEFghB8jjCH++i20q2VP3Q/lJujuPetOJc
5zh/4NFziGQM5n1e/vpaA2FITNRlsWKxHePiiqruNYYnha+pHjoF7K81DucXJ5qFS21+jDCrmrPH
JFmcFGc98OSUAZ6tUC1WtQ2knpXr39JiBb4BHEcVGKBvWsp00rie7LqFRck73nPC/n9L9TcicTPz
qtXXIb2KBEpHDhRR1svNIGvbhwnevPspU91mqxHFNuMHizuRkspnh0f3rhdumk0FYuOQADxE2pP6
pVkQABqk/bJDmJER000Oi74HhoArqri4Q3CN2Y5T9x1mzclOR936zA8VrWT+09etKsJKpH57L6NP
EKVpFdMY81+5NXxVF50kJtNDE/BwFicFD9g+sv6Ckr65JW5gA4pNXlppAizA52NHQwe2MHvsAuB0
sKQ89I6gh7D3iJ5iwXKuzXxVRFMb+5q2oUS9wi23PgNM8ZVWHCSt8qafF6F6ojB/j9nT+4FyRtyg
CHh7PVn3wLQNZ+IgwvfEorGBTWO+72H54hmLTFfdgTpc6hpmRbmdXG0PEW4dl5yoLmfYze59Xylx
WXMXM/VHP45U1jv688PGp3W7pr9EMyyjMy3C2N3xpwH5zotKBxAqQ4n+2VVVfVe95cdmHgZ4ejmk
amAnOJsAg6UQpaSrdKqDHFYYHy7wR/Srh1WG91F2OiwC0vdFAVG/bsbJi8dnnY2xQBv1QHGY2jVB
6F7LveF+9pBgRnW/dOCP8VH/1e+bGJ7oFodGQPWOyyS5lRYOnRtrteeftLtkMO8yhmU7JngsSOh0
U8HAU+olCYPIR18WzwQI/JE7xGibpmLouviD0VkLutYbQv0isda0WnqQnlaSnVEVStNDtlJ0bpzg
VbdBuodaf9jM7SFD/5nDQX01ceCx5kzL9y5Almp2sXz7ZCw1r3umc18csC8mUZ7EwZWKDXtVMX/X
MB+Vde5GO38X7CGQT+6ZQkeERKsp3T8IOn9DCzvQaf9osmoT52UEQTWIuUgwe0DwnWroQQ5OvNk5
O14LzToZw4CT/8XMaX7eJknQTiTw/GtGRxxcJCEuMDSiFvE2ww7ZjkL72/7BYjnKf/t5q4OAP6M8
ERcHDpgEU0egCNa/XBCTnQpc3n5ZBlbarQpc1IXDyX/9dZou96/7QolEDvRDM+Nk4XYn0MpxqBA/
PMSs0WPofe7bXMLnCDMke95ZVOq01y3MgXMxziw3FIQMMA9i7i7GRKTaHuN2TzxqysKHLnb2Nl03
k5F096rw4UkVom0tpeqpvzccSNbtURPqjuGFwTqJ8HDnJfUn73QND7wnaL80pyf4vCYLj92w7x/3
OC0igxxuD65e6kkNh9jPjjdh2cWXjGyN2f3Q3wN6KpAtXKTUxy2wjNGXoc8uuzYsVFeczcWTFWyX
4B5O46rlFwPeGA/Dz8mqHcGVF1hjPGKw29TWFu9msiuV1GJIfFGvosLTVYXBt+GLX53kTKg5mVDT
FkxlV/e5RZHf7THN8wKrxOp4agoprFDcCK8zUzzLnVId3Rz2qmGgV9eo6u9iVvErOCzdWcEufuO3
/XS+x9F2McRl6f/uW1zDVdTYqDjC4+icgmKg/Q6I5C//fpTrXkIiTlTyofQyLZGESsj8vd6aPIZq
k41u5eUYcrMmogXIYq2WQbhdhxP2b88mLKk3wqJA1Wz1+kCexYXUHYOj43W4DooKZVK3cw/tuLeb
R2uxk5apAfFI8D2ihRYheStwePRnEwM+d6vcCjx70tRB8ZgOnqGETSZYDZ+c9bvbkPEdIW+DM5ml
+AHNa0SCTlsnyd2gwis2MB0hB3KHDJdHmarpKDJh6CZO93G83sYxrB643ep37XBPbhq34HYYSvXS
TJEqMWB5LsXJjObf9dFOdSygX98FYSvmfA5SbskQx8g6hUEtOUgS8eNNhMDbHaw2jstoRd8MM0T+
WiCv8WA0wOMmCgYJtokx8WIk+cqDYSME9SmVh2SwCqDrhCNv58Kaf+6qaeEyNO1AqLN7+EjMZHlK
FL+w5tgA5NQRhok1vBucXTw0r+3EWpkPZGPqmdweVVRcjzmRJcNhAdg2kvEUrv0ls9ngvnx3h7+0
7P/Mc1uNQSN3kHHxXIw7fHvyin4/C01eYeLPcXWmTJ/6RtLzY3r78BWAPRWRyTIWNhM/U7TMEWpI
5qq3ThAgBFraIghHD6oxmxnRIvf/jNhl254UGiprIwmEDDoO3i1Y4tBVzhC0zOrYUlX4cWO1NdaP
ZY/TnoBgRCzjJKhkVlJdvOg5pho5kVwdX43kL0tGZNSgXwGmXZ47bisoh8nvSIeWPhrExzEH431K
eOhbwCHBTMPaER7rCUSuDm2B4K6a8rCJQWxuwla/SRYdrZJB1OZpJGtXxGaAZ/YnB27wucUZVjIS
P6dEtkdxWzMKj5g91OWXNW7QGborZ4eV9LuvHPKjCmutkQPENiZ3/B7WWUGzaVNz+xh3MM2wsjLs
elHga8XVm3SpIn6gFL3rd75dG9tAwItao+yn9bl1Qk2DCWVptPpO0GBHe8+yYa3uB3EURplC9hAl
uTtA9Wz0wVVCVxMQCLF2pcfBHSr35gmFMfmPOAgE5gwny6xFE0yAk9IurCKPfUiiCNOrGDItDLKV
x6Z03LgQqH1SPFCeRJQWFkUXrx1m/NPttuvOXSJvsPq7fzcYjzvxsGamO5xXZnrkX48T+ttH/wNl
93X+qnQBlIv1Kbadfnre5gA94r6ouVQA5nzBUH688Ub7B6BFnyKFUGLLwWQSdL9mNnGS9E3jTaIT
MBrViH0dA9OnxxgWQPoU1ojJuTRAupyyqMRvh+WuPlwRaJXnxhcsbjmydD/G7YMlfJJIezQhKpNo
cM7VluuCpxv4feh9Sm3xz/MnmzWRYt2CCcTwDac8LReTO8L/xV6qeLXxbsMi7HPy8sktxnStnIaq
UR67FNu8UoGomg6MEneLfKyWVcdZSjJFamwxi/GCSZD+bks61wE9w1Hd+p5+sIi5DnxXEQbM0urS
6QJIVD9I3XVV+XpgOj61VGJn45SzGE6k4tnf5J25opGmPevSi09Y5q49Sdvb49Wfa5GE2kgSjJdP
Gff7iFYPsckMiZHDa6U5zLzAtiZqxx8o1DxOo8CGmpT1FslTfN/eRPW78ezBFuSuMz8H1ML1r54L
VJl44wEVWzjzh+Vtpqjr821krSg4uEDH9u96MF7z0kY+7fRoCMJKW5jZRvt9+Hb8QC4XiLKT5Ky+
pMiOSi9B5pHqRi4VhR5p3ofvLwze0YvIVj+uYLA75eSRWvm6jFVgIfB6RkBkbakn4VVCqvT+n+qh
Uzn0Kn+u8aZaTK2dlb6jqF532inTfAx9mlfhQh3THSrBHvvfl0zBb9O0QlUsQsQrqzEf5z2fMkMP
VND813iGs8ry3QwZP2oRKTZ0RzjxuOnf387ZJZkK+jPR5UwyAXNnRkUHRCvKYFVeQxx8r6fHej5u
x5oafY/k54u1952uxIZaJThkK0cPEWF35z7aRAVB1g723bzHhb671DbkkxWlyGcXcotfU7nrpsTG
cNYylX73woYmdtDK0OsUr+Os3PwnA5+yS2UkigZLbLs70JIjLE7+ZIPEmm2CnpzN1TsX/nJLiiEc
aAE70op8LGVgEupNLkBj2S42KHZBA2GRVfZvScjmdLFG+Hl+T4VZLBGey5CzjhLbORjDLle/iW8m
MhUyYi3he/hJoRQa4mFAo3Ovz5uCtu5GYQvX6cdbF7zwnvhx4vdXUKAizX9QwnsQiRH19FAH5pbh
zgmeY+j+6kVA+JXJEsI1yRk0h2j2TSpqOKnuDN3eeba+agDN0AdLcqmHb1fWXYC3Nho9hyO8c06D
swa33MY6Zt9bNGJo0JYS1cqCDU1yT1w1U5MhBDBNdjDDPneZMY25FXb56wjhqDWxavPVlbWLGxFf
ssUhFQbSHJSsxtyiKWk0rIULjD02mjxDm9yx3sqP2EDTA5Yar2n1p/EUZPhOCXZkCnc82brDiSzU
2poTfPM+2EGX98CzaQA6njpQFCUGk/HLmvEQU1uEsmh6t4GuDC3+W0h3MKDrBMO6iQnuxw2Rg6en
MWgymXkEYjpgbzcL4D595JuPyk8+8DMP+2bqiwiq1sCd9aR2Bmzt5w4+QPM110Dcqg/qq6lkl2fL
iHXKHOS/IWKQTC6S3Eea9SGuGFYm1rZZdmJ9fBLjNHcnS6kTE0vDIum/xyjVPgKCKrOhqOr/NHgE
NaiMFMWn6O6bDyGgJoUvBtcw5A23BZnNVX0eps12AAqQO/P8UyaDbbZX/eCXbZR5xLqJO1nIZfIq
5Bn91HbX0LKHdZ3qxpL6SRpauAqSeygJqbxVTCr7EGA8IkyHgYOrlDzRBxvuQdNdtTKlpFo0Xbto
yjM/5VlPru/O2YPwyOYUo0GDI9HE1tAfJvlafpqr0TxlLvxxWbj2e4StLigaGVnGo7wA1V7ItodA
SBCptyzj0SsGrVjBiR6ZL9GJZmcomJzsuLp3IXKeOz1mIHtU1wJbfgmUJbOBzHXBcdYbc2ttAv8q
bVkYt53Jr61saGSoiuKyef9mT2iinqxaAKNhLHECzn/yFc9uMmCDasfAGt9KG5D+8XL9Je59eL54
gdwgvM7NGtRzxY1dwQfoK+KV7nE4NHgF+BH0GXBUc4kc4DFAHUT28IrVYvzVyDQ/VndpGhJ+vvGr
KT4vlpHzk6VkbS2J0/34cG6ieAcVdK5O/7W3kU0lDK/SL/E/UQbjl+KpQQFbVO5CoT8r1xRmWNOs
owQJ+WkBLhVdWvcaaCrqt+7lwyMyI31gc3+ZCQ0d9o0d5owDyN+7CjFujhn8UisKk+xJ+iWAX62H
Rxehr85z7gZc5EE45SzVHwydMRpEZewpXEIOBh83qMFKA6eF6xwH/8SO2pC8yBeBkjrnyCr4BErX
+ML7MviM/SUY3L6+8VqMRK5/yvFiivRSP/EDXRTuo3KWYnliJ7cfyRnTk8pQG90GFJgWrHQwIhwE
1W0wO+Qfeb/ZmGwvUUrh+eqHIZoes3G1e/udz8SC276vm7scWzg4zMco1N+4DC5K4e6V+8TrJQST
H1rnjR0U8cvAhkNtvVRJRiTRmCySbH1jkvQXTWuYyqPIWD/BZTOHNaxIs1DmgCb7+UO/N15mgb0G
R+JAIVqC4usgcyTSzRF2oQdnKUrYQDVxO60z6snc0vbwnclpsMeL8QUq/Kz1bJJzbPyAKmC7Mm9y
hl7zsym92FHHzNLcdYKRVNf3gXgY1iNu9sBMZsZC3rtUusU7/C0PFhKZdr5lDZytr1H2Zccucy9V
KfOf/2TGk7sn91b3dC9My/mgHLWXOoLhERwdT7lnhMFJlB3J7lt/h3zN7gu1mzk7aLiB6XbZBkRn
K5+azoHC2Ke7fO46K4WNvs35F97oToqGDq+51h/B2JI+9cav5oX4D4iFbTOQwTWc2m5+EkeZIkzd
A7whshif/4WbOMxYED5FUugLZsCJO40hQlEicwnowKKbXlBlFW/gIPmXk909Ah+hzYJf8YZmJhdb
XO33A0ZwkmptGFsjnV9ehRaPK8bomfoEn94f7rEo1OhajdZgd1cwVc/xMzYNPjgDTcLrMrtRX2Hl
/ZRiXJjFj/CCjMIXynS2CecMF9qTQsPXE8CrK3gQqebtUpLmDa9uSyM0CesenbjFlMmCjr5R+BOw
gmMhZRU8btt24026BYic4O96bESjCK/Bi1wjOaQV+hCaxToW5hVnSIxLpUZxCmrAFgSP2dvAD2+n
c1UtLqxGbefKrxCtfnJuPn6PKt0LeIqloEJ8sBC8qej73mb+E2A390PXvYsE0nvnHHXkWBYlt4hl
QqYxhkP148vk5IQNB7Z7/ZfouhVty+qmlhrsDf1mFXTbNkpdrCteLN/NeagrLEKSD6Lbpy5Ig918
HWCy9cW64PfDljWs7B/P6iyTJrVP3PCFxasnrn6ivhF+8c2LD0obIIl7QcQaSw+Twmixv4JtQXiy
eR8stieF8iu4rKu/OyhHKBuwLMrumHKsYsDVIaYa/bvwCkTBJ87cPX5CYcfU525v4GKbUw4FjzLT
dQoVVn8zBxekEuT+lpS6iH0Z0GPZWJERYWVIkMQGt76WtAuZ26uzTKg4nsD3ugBFAQQ8JWOMPo8+
yuD7+cd9CI4QsWrY1QEbyBLgwSu8MemxhsqYTE3AuOCmrWWxuV3ZxYF8oW87Z/gMeIzmDVdcCYgn
UWNlqjRZqLx74r1aYFN4GP/DZj3aFeNDp6xJ4zOo5N33Axk7RcCKxJntpOCoXeLDjiQhuJfGkXET
JgMUi/XlJ+XEWxnN4k1zhBWgSLRmZ/rkMpnsprUfm7LGUyMT8ZrziixbNtwPd0jU5mh+B3Hyp/Se
WbxsM8YeNaPKP2H7Lk+b3hE2IMLjqLx+NZZGKBZsY9cJf0Q0CspB8LFPMRhPoJ5J2+9IzMB+DO6/
bwZvW3/4JmpNMl9T5JcCgrqluKCZwIyphn+rfKn7gT4yheDl6RqVkOSmul6gDcQuZ797bwLj1WJh
IYRqEr9wr1aaaHug1dY/O8q4cZ5PS+D2REWhLsBdcTM/Z9ls8Wxe1uOX25U9Uu1lJsSeoJznGGEC
sn57ecNPqS7nwNnM7FlmTJp+SNkULhg8zuMcZZP8Kb7WxpG2UQ+eno794gNdjIArXVyLO+U2kyO2
DHopQ/Z9NVbJ4gTKZwjQIzgFeqYQWCjwsVsyxCSkbughYBc2hjg2DP1I30W/KR9LOT+QAD+hrUGl
Up1Zk19hKxn/V4FnwW+RI4O2vBzqrHt5Ld+q4ZwFdUwQwfUVP6nr/mLMp6yOZsIydwCLHGOnY2AW
d6Ewib5OgHEKz6tSjzks0fQIej4gcn1evYtyH7b6dP0mo5XkhHVXhohjOFKLDuQmH+wz/bZ/b079
ZkM49PJjrHx3YdsIiTIx/Fy5poLJ4R4hSuARlAtn5jZ+Bnuh3uU1zfA5Ii1nXz8eKNkOw0cl3ugm
s0KWTSznbEbSYTnfAoHJ5qzl3WmGS2KNJ2NGCNj7gSdohY8GTXjS4pTJ27ZJFEbc36ZUmk07JC47
RcznK4Bo/gxlaw2Pb39RBwaef2HjzVA+w2VKABnZD91OlkmMLJdcY17992qpel0HBFn8x++Dwpq0
duJRTU5HMtVU7rb62nOtQFJy3/yjxcJNuG29evLWFb2rqoVOQfq1jl0pz3weXZl/RZmsxTOD6OvU
mxaMJv7vvVsCmQ+AIAMkfxnXTqydCKU+lm+5CiE/4wgKc0FQZR4QC3zP3NpSmB8iH96NAQtB8Gw6
v2bjxaPgXMEYarLvh6e8ytBgiR1mmwnxaI0zXzQaBwREsOa8WBWs4dXzKSJPoeLk8qZNwRbblXc4
BTjCCOiJ5LqrKrEFgIlRWgm82h5e7+FNN0naZnD+Qel5Z6+y/wIiGtmzCAIGHhNN+dzVqxEAhWnm
L6PMa8aOWS4sRsMhHAMoZ06xo/DVjlhRq4scT/pLpuzcFtnElv3D+Q+dBaF5jGmifVBq1cO7/4Am
kSNSYDNqldMeeMh6rwWVAArlDqRl9TtbTt2boN3VYbvtb8LkNHvrpilY0iEj8+tQVmo4E7xksmCe
sNeGjRLlfuK1K1FL2e0JDornFBtpDCeHnzkjwqYPcXZJjjGD1AMVqJXYrAhxWsZiJ6iDftZCJU3S
tAEftEuFe8HD9UY+Xw0aYNO4LCS7IQjnZIDHgcOsTmWTqA65+l012jFIuBsJAHkkRJqNNKbRVsGl
1xGvzYRXjT9eBVh90ooYvKz7Ig57N2PSSNTIEvJRt2HvBTZ/M9u3FTvL0vTGUgxyIkf0j9ipHpBB
WcOSdqQK7yZVzn2JE60A5lKwliUoWVcrCembvtkNhjl7MbaNox8RuRAvcKk8372EPNsXIRCAijQ4
Kz7b4uEsGcga29co+qka5+BLHa0xa+n59SY4D5/I5xJJqkik9fZmLaF6sh2aUN0UAvnYtRr87RpZ
9hlURB72UKtC7ai/vyE1XZ00BWMTlughuPJ8vuOxLK+5rF4pnyShsUSgKXsoIohwck+MCAz156Vc
ZfKa/V5pnH+tq/Hu8TyGLV7k3ayGPbcMlrfUx8Wn9bMJa+bbhX/Ode5L0QvMeMaydol2QpCNaINU
uQKfLVU+k0dkgurgCOznEooOpIX9m4U6VNMhOWuoy3yhRKEYwovfPk64iz5vhzgKIwypITeByaoU
tSJO7mjNZlYYyUzJ3Ve6fXiohHjWTwce2TearuiQ9Mkx594dN/0bxn09HXJJa5sY48l7/f2zSQ1k
JkKuw/d3QwurKYaVUu7+k8V5DBs0TVnlBg97Mks6DzdmZs6wyRkbuD18gNYYS2/QurerWHJLDEe8
U9YTzx4nEEwSbf6mabwal7yimrc3V8UpHVVCmPUA9F0h0FkX7VViRRtVScVVdmyPPFbH4Uh3g0Gx
igjdheO1fVj7b42me/LvUbSJNeHWUDHZespIFzZlBbVf7z9H9o35yeWgnaMVG/bbeknAU3YW6oxp
PGS1WKGFBN7Se+OGlg8k8dzRV5o92Zl2D+OWpETZYsQXN+PKC85BCHdGqC0sFMlfICZB3Ur2Ialp
tEWippbrgSfjpve3p0Pv9pV2Z3zpZzqy+K54gLWKaKjsFbDMMoPBiqc3573OJY5I8zGQEuUqtWIA
dLNINxugpkYe2Bnb36+wkks4aHQST4bHekrenrkAgKJWgtcOo0QdgAztRxCqypyQAwQbU3MzMAvN
+mzhig7St6pUVxPiVYLy5h1yrARYdViKMcaSEgubufpRkPVEwyWPy+Sa64zoutVJDFd6+TlNIRpV
v01hn6zJ1q2ppPKAu7Lcq7bjM0pY9VrBrn6o6HwqtnDgoJ0uVrTeUU67VxenV5cSMV5nuXHuK9pb
m3Zn3AcjghFMG8CZA29QhKMntHbil1DC+yMqnMBlRqlh6LiBmXlzl8g/R0ilWGLKzdCEHXbRfGvG
kFjnNz6u2+fRLb9m2MD/HaaydXeXF4sFu8I14Si0XfaHYClXQ4VgRaxwbpUltU1I2VrcYu52KroT
OQ6atY0vh3v4yhnovU59HvZcnXnQvIir6Fnd79tUsAgMkpYzits6h7CwwmdiZdhy3+SdzB6/hbbZ
XWUpKh5suZKjBHAiceMwWbuScjLulp6vBQUsHuWcvl0YYAUGRoU7T8/nnBBDEdHOVwMYTuy0ViZe
JKNfG1i3Bi/QuD+Nr3qrbcJ/9FM7miv6FxgWYP6ouHxKr6VAhK1NML//8me9vV3ujKXvTpszy5ny
B0pub3rCIVDOxOTzGx423szMLKCrlhiKWv/ngMVCJHwKd3fpsy71aCBf6rb/2kqQbUHtWyEzRR0I
5OVXpBKSocauTpn80hVhzpIrxsYV7zdq7phQYmp3d/jfd9do4v9ftWyZWoAvzNo6vvVpJjVE2SsO
6IqCj3h0TeGelzbtJUD7RTZFkvgz2nN6aVA/vwGePZjhBWattTrjHmibSUrYHb6/5qBohTtQf/I6
Tn9AgIayWAVxAvvTUigjtzdoLYxizrGIGsqVs52RUyRxrWv69RDAL031s4RV9Dt7cJGxHV61ITG0
y8H4toMyjG3Kri8iahjxwTJYba2aBC4OHKA8PiH2qIblPkm7N2wyzYO9q9PwPnjVuUV9wYDa3qEK
v2tRzkAt70BtaN/p0a564//iI+qm/4Lp1ed031N+p4+ZgD7zpbUXzYYaLd+H29LXzppFsdUmF1xm
Wm4F256IGEwd73DzltTdAFDofZvEkJd3qDbkINOWOkPaxluphadODRFc9W3xb4hCQzuWtfigIsFN
XMryx1dxlrDpc9BeBJAJaJ0I1zJq90SUCTNHBjaRQEjulLaLIA8Tfpx9uiqTCpa7PoX746zQ5ZWi
dX+vAgM7/FBYwQ9dhi7M9ays9fGYlLWEdTiFrZwZugywHJjAmsQIEfAORHnT0rx0CP4hGRFBEBKx
iEWpmZahXHjkUobKVRw21Hqc1nvj8E0W5JWM0+G6GGgIfxejdcKvdStNigWTrwojSHxmUAlHa90B
cfLeGgCnOLWhXAcbgiIjjJpib/JGhPlre7O/AMzWOctPLi22STXut0ocFT0AVythiwRy11YC+ai7
nXEh6Qu6BrtrUGw5Uh/G/9unjeag/nbQpjwFcP/+og8HKgNsoFtXMMDL/xx1vCmIGVY1Cp9oRxxQ
8DplCgpMFAdpwKat0VbSpeKx+8ktXXloyglYnx2ps9y4luwi6y0pWNTv4FYsLVNdAlHmQdFPxpzk
yJHPEuCqN3mHzrSTiP8ZWwNEv5b/dEeaKn2HAvceZWZK5NClFPznnGCMVHfusTC2gOeAbTJ2ZQ7W
5cYAId9F1RSGVQV2xDCLlOcaUG/vx8/pR2brQcwGh8yRrfl7N8rWouOUdXMQdMJPDOXSLE+iypRV
vkpNqCQaq54sVaQ6/eNPFhGZybOOQPTvrwEn2LdeCwrWUVR+IPXImHlify2ELbBJg+BGP1wu9Ngy
YLG5ViYiGJWRDYcBeBCZ0TL1oQVUuA9fq6BYXPmR/2vMbwkMrlp+MpyPQ1FNGzAIE2nPTWCRQiP1
+m5HGyes1ca7HP8vwIr90LSBJszLLUxr7pkpNn1teCTg4REjX7HuZ5iHQg0mgXo/WFmUoxB9/3BF
4KkKw9f5Zk4AT+oM5jEeukMcplclh7mRpp2A5GOKHAlM18hX0Mpw14Ksk8BBrfVQgXo3fpkIDRtC
R68SBRD3ezTqUC6pj7rNhWRiU1x8SXOieIVRIzalSj5uFWOSha97SxUesAbfkGpUkO0AJ4HKX+P4
QH1ENlt5OEjg5XjNB+mYIBv4HubnQTfk7f11mQXdumsMWzG1xwmMuL1Vbm5LeKlxtdaCxI5wofRC
WtF5yWlwdcteptTQSqP1LjGeDsuSEiYTc91AerzsDUxZEJNhGBBgmVHPa2SMCGtDAyqsqCZ7UPWx
9ZNG7Mqcv7Vq6Twx6PLvBE1rg06lGTTpDPGZ3vjhK+HUJvpEv3kk/P/FtHyJPZdaO+0MLD2ld3BA
lp9IIRrJhLAmJsZkQDlV8lGiasb4AYfqPhrglsPfj/BNluHWACAsJy+p+zu/KYDLXSEHq0Zk2tPB
Yd2/JuSJRsT5fN/23YeEx12Fui3mqvG6g2vUECNocVFEZedF+2vQ1Z0eSfPFRsLq7fTe9jj/Z5hq
rniEhOSHmcSidMQrpOYGJlJCC5hDE4IYWqwvBIc5y6hqdRrVBY8xxJmdktnOb8wtJlW/HgvDZtaZ
b8dNTQiAT8omglCe+DpLLYLJxp8pddwMztL2hHjUoNwugowrGxetpE6Ooe+F6pKLeIGZzg0kYYRa
3ceOr8pyNXI5tvwwWVU/Xz53/dVgAFt15dipAGEq/KcYYDxmkG/l3p3/8goLpZP4gDQrTY7XBIKq
AeVE1pRGM/Dl1yC7kSKpOP6XgIuVg9o6FeUDypGsYvk5FH0noNLYYHoRXd/DRXOG2zmgN+nZ/SGR
5/4Wiy3ZLOajfnqwbv8bE3lVvcArws4cHdmqpHzWy94wIXFX/AtIHCxQR9JNGJqh/gznEtNIsTsp
reNyJ/xPNSg/f0UenOhXv6N0ZJtsRZhtxGvJa34IDcthLeAtZ8YmmkLg88OL2cuSRDaEkL1DMXlp
TTgpCk0JBl5099+2ajMz5ztOdx2rg5JlJitr8Z0INkDs1IASxaOeJ1TKjvur2hSBTAGYxTVQL91V
o5jZWqZ5L2VleFnzQGbruNOj38dJcX9mkllBHN8iMkrzJXWK1V/Wvx/3Wsu14unjqyONmBO2NL8b
4YXB82GZFwAzpPbYTrux8pnf1cK3bKn3EYljVDty2eexqLzPNXtrYj64L2ibVqI5zC/9kPjnUc1+
E56h9aSOsCT2cLeuE4M9HpfU2v5AFZuNHgU/OcIPXaiz/QTC9snTd9vmZl4gdw472Qshg38n9mWT
DoaXjxWdH2QbywgaT0mh2w0Hy1WaQcQCZHF2TFtOCTrM7e1OrFy+EDnLma6KwALUwqhKzkoXqONb
wWFFwq4sEMq+xLieQ5yoAho/3QZbH3PjLkL6YeY5/mNDcmeunNDqci7T6LKQzsxmaw6T5W4hL26L
jSXOpwJbkURo9d0McczBqjDKSxahZGDO1f53y0DeM7GjN+ZVwQ0bgpnYWBtn/NbRe+DTLIXUOgMh
vZHoZx8NeJdaD9xELZAcS4iYmeGEhmEw3X04UyF6QU30ihmd9FulJq9YpSQUy1kJOa4JP25Ctt7n
NaV3iDmMImij5B51JLjR0wpE9lvMj1R7s8muNpgye27aKdAv5AiCemooGMUOKafmt2CK/FMw6C4P
h7UBzcmgMsSpbdtmFEPa5bCpJoIWF3UXLknhM4FzKvcG8B0XoL/Gt0QWJ9mGqcC9P33IONDKdJAp
LdKubH75fgwstTCrB1pBPAXd5jucHNKDnSdGkoMqap2E9xC37gqexweex2MxzwKeJdysq3wpeOTH
crUQxCN9tjLti2icbGYduYGKcMepTOsExnHcQktDiCi+7S7qzUmTdWuteWrz0x1Bwa3Ins7vZX9v
yhnJGGTsGHKT4sse3moetZ2YJ2Y/Ru9gBbli9GPlT3Cmb2BqozPHzrSwQKSa0In3P2F1DjpngeLB
W1Xe9TN2xdLubI6dwdltWnJ7xWbzyBd6zzWuunQsBiXpSDfEdFhLhVgVz9cKccBVZAWpIryPaSu1
wUYQCAcGdtNbmz8+byjijDsnTiIJjjjnZYKdyfQjQTA21tKAuKROHDwrUfoKsOgZVJwDZc+E6Fgz
vdZtgoqtZXvF0m1ghrNqGEAICBKh/0X6IPDJUjqk2SO0viQKqbUJGT7cs3C2ci4GXNlg7tNcw5IU
x4HGyud5nWS0fzlv8KVpscuC1Npc7A1Koed32ZVHzKVKjkg6+U05hKoRWJWzxOBI2rHJ8g4OmLKg
tiMHAqcZuaQAMddyWfzNZsudL+fUa7NhPTx+8BRNZeDFN6UoVTfDwYp9J9TVz9OsWQTFtNtwjBHF
TeNiGAYKt6rXQLsb92KBV5j1cqZm3qjm0/1n5OpXJjSWgJN8UHCTuWgEvBd4R/VZf4+X5R2qANzf
JCjuGruS4e+ZNw1nSgT+JaNruNdfpOOhTQX7bYYP+T2WSHkawojnRNWPZRCvNQ3PDgnhRmNVKvFn
xj0SEyvlxjp0plP5U1oCJ6Sen9cqkleWjG5qxEn5FVlXu2h+FflwFaqPmByCRzqS8OTKHTqkNoBA
r/9L6j+VHzVVHd/hm9YhFON5dJ97NV3tPGfio8LkHlMr+c/ojTX0ymItp3ANRxdZqDLeNqPC1YGT
Nwr+vYEzrG7Tinlr7Lbsd3tLCvsvfiqnCSpIeEvq1x27UX6Q80+I04TvAxi3+a3sDai0HZzxX+1D
RF2FPrB+umDj9NJygb2mDzpML37Hn9vH8CXWmwuXdQ/Pedxwgtg2AUp95AXvAaifDFMTCTvzPTRy
vfLhAJkVXObKIkMzCZWVd1HQvDB2ESKyWnhN9laWnMAGFDXo55Ps2u7m3QSc7cw6okHa79xevvUy
/2InwkQ2WzftJ8ezuLeFHM4aOOS5yYGbTyUbvKjgeMtGhalvYVPBureNFp9UahvbWVDSqteWON86
KnZmnAJhV3B2c0LM590Cb/Lq7AQhFMxQbdTuXRJ71TKaWVbGF1Yw4skRynQl5wucg0lJOZ3RoGsn
IShshiN/o72wBTOE7NzwzWFz1T9glNeaVw+2Urdrr0cWBZLz/ZkHfbPUiVkVg91Azh408mzF57yb
7PK0NRB7XkavFUPnyn7JJhJIWoFFN/aiQ4/lML7ZzTEjB387ZyNPPh2kggPenI3vBoj1tlH0IeYg
l40Gsv4GMf/UhhELVHW8CmlMlk+ZN7DHOz76opEkfeKV969O1NYzczjQ0qSi9WmrCLFvOmD/vbtG
FSARpUx5/34RBb7s0IKckLCXPfMkRPfiqCjeNBuaLT7sYzKJNEGi0QmO6vz64oHlA3ckmvNVGsHZ
ACJvfUsEdkqOTRyng4qsRBtlnBPzpVTjUCI74UvJyK4A84rpgZFKivSUnFuOG4fIrMVZm/eGDUTa
KJ2lS0ZLg1CMnMq6bVuZTelsOmi26UPEEcmpMCsoDuhkBWGtgrwpVYfpYfYD3hITjtInAPSyqF0s
uGUJSSGqhAllgMQvj7OSSE9yFXCEpoaeNBWR9C5wQzKFYp+OqLcY4cMvdAeiCOFWMJFHyZMlZbSF
b/q6DsuTy5LczMB5MARRTXThFOh58AhU6QQjYC9Xx1OuMvFYwVV43sFO/p+B+RQVD9OYlOgiwSQT
VPIPpwQdJrBVQxxsqLDlMkEHqdGGnUcZGFRttwZvqu3EEjllPs046I+J9k3w7wSuHysdK1MkqE67
xwUijMqrNbmkdOBmxlKWJieVq0NJYaY8GWZLuJPy3ME3ndwlPYZD6mSoKKQPY5wyErTylYW2zf1t
We06rrL3FVRViDYoQUW7BX4QpFv33+iMK8bwc/kH8OUQqAf2DoVVu1XdNhVhRomH2E7uR8plv9F6
tTvT4avz45nWt3EUBMsgHqgKM1KtSCNENOSedEwh6cZLbt0CLaKCR/9CqAaNrr49EjJk/YD4NFtN
SxjGAkkQO5jUDTFSrgWfB1cI1H5uuWMT22ndEKpb9pI0ljAPGhLjT/8aOfpg+rcKlX0jCwqxEA47
FnjLoUeVUKeOSwj14Dh0JaFJ1gINryKIPiH7/tNkEldewn54LHMqO6B/vjgh4HnBX7TpijTQMJh3
DPaDUUd1my/UpxoMUW/4Xtmaus3mWp0+O1AC5RolyXCVE6xOnFK2fzp1s2rYkj17EKROX1gbv885
VNMCauhM30CItMrH+k2wo/xvqH3pa0853VU+NcV7RyXFMR+p3xzd9PgymyN6CegMrNNqXbSC33Y7
+1PYQJdvFGqrnGhNGC9WLxKZppJJGEyllzzezQfohT9LnxqFhKXeUov04cCwYreSLOayNt8ryUNs
87iI5VKiC4vXMFwqQLdqn3YGWK6YRDJMSCiaaepB0SalM8MKx4kq4consuDbwdHzHaTdbRCd/vQA
94RThPpuyvAAhhT1CddUH0QX6lBBLrnvCSrapEyZ08u9Vv9OQcDr1qdoNl1VCYB/a4n7eYbPzpFo
Dkq5Fbj+cPpqmi16QbMXFN8jCo9eqF0Ze2iTfpUa4sL1S4c7CmnjLfaGOpaWX+Tna6zj5XvZtCTc
hHJxj/3LUN8mRUjfY242U8IwqUp+Mq1dzLQwxjKK88OQhPX1IOUrYB6M6k0X52w9YDt8TiqLESpA
OW3SCn8rG0cBBLt0ixZndvq06dNWz4EZ11I5gZXS4ZmTZ65UcnbwgFAdJTHnps2/nUqZGA6jZmv9
SRN+HgITfG4JKbFDrmxi9Rqv09QLo4B/c8DJZ81S6Q/H7iE2MXf/zTxP8OZC/ESmNWnWoveYcp/U
1KnECjlXjVbKSWgudMU5g7qKZblcTAKA/awZJqax7u7OiSNuk35ZCpBEclkde10K8x7pp0GF5uxe
mo6OENSDg2rpetvMqDzIjKecP1J+bfmvW02bxdcp5RlK/Y1hqaDdcUFWg7Weqxaxp9a0Kwps/ffu
lvZjyS6nj91AVeUpxs6M1tAeejO2st//osAK1FeXKwtaDIan1Zvxqrhh7dAcqMZUTNKtd7Mim38m
JKFo5/jYXPVqOJYwo5ftcPSEI3BlnGFJ6/V+cDm84+3D3margpRtxZ4sbju8vF58oFdgI67v7BfT
itI7iUxZ8IlxRb61K7UM955gS52Po61OPQ3JBW6Wro4DluRbURlMB4CkdyIBX+Ww6TuQXvqGyOX5
SkuIB+bk7pffyuRQizDAYlDoz5oIpXFbw/8Szg/CY9QnCAtAqEQ66/USusRmxdcx4U7wtUfxRSBG
exsYZTwRe4I7KK+Do4ze9G2oedBLPGFuHPhujSFr7qoe/8d2goqQEL1soAAT6FBPKoesmWp1EWEk
HqX0krPmgxg2+TP4uJDeSx7Y8Qq+9746hvmO4SGuTFmHdqZofkvqwMir/SEStdABxqbWndGr9TJp
bdd5zC3xdWRn6YAN8Pstucw4R+bko9sOYQ4Toss1elAU5NH70FgK0OwuX32qyZDNaUFbI3RtYwo5
PBCJAVbB4Sn9IP8vuvSzCNrzN0ueYgf1MjvGp9VHP2VigAl732ESS+cR9KugX9tvae/CHa/V6QI2
pou6OM+D2E2NL3gisoGwZIYegIZNz9XJiSVHHkwnDMaLtsZ5fUkmR2L9LSc7Y7PeM6mRL/mI0n8j
YQVI25e5t4dXAlDFty7FzFdxR00BzwGtxJLAyw2N5q3PrtBi02e6ZIcVxwW4Nz1VEozjzbfd7WGQ
JxMewH7/sBikjU+TwQf7BfxH3eo5vijn8mYWZPPDpyK3ZgXyS2oQonr3Mp5teeqiU7yDEm8LK4F0
lonZOjViZ8i7ygOckrt+D/6DwWqfGmz87gmHeopSAW1L28/asyZtd8/OrKmL5lcLqpmb7T0nWeaP
R+uThuCS3G6U+uXR/RmXbkwYWv2nDTrI34RD4dhogjL7uW2ItcXJ+OhzOeUaC4yvagQxjtLUvhgu
B96MmzkegJaYB+5s7gaxY5Oe++LAK/Y3A7XFQ9RqbN84irfp1V6R6Vm0m7rOBKLnSH/TtqrU5+dT
TMBKkHayHDPH4lm7L2xMJ/ycuqRH9IgxUNAjj2kRGyf3+MaIzMF5sAqvTjrwGsrJQ88HvJPho+E1
PNz7Gxhpk7xeVgSyiqKvOYhGkacf105/9z9ttcBMiyxyRE2E4Ykhmw4E/Jqf40dbYBuI+i3JlQQE
xblqVH+W95gLNm1R1xLfckkBGG14nU4G5+11zSXhxGOYjBL99QZAXGPk6u6OpHTVbu2w+DSfPTFo
kK7S4SdygFk3rMy1LRNoVwBTWhHNrKnmz6FdClt5m8dsblgCL2It4tELZbrlvsfwSWTGP8sugyim
lJo7TnS7Zk8fPmQA3iS+FzCMQb45YTXm+otTDoXq7IbXkpo4PvSyPsyDNS0gDkQZyFZr/LAI0Qwz
SLKkMpFrSd0cqneETnbxIge6IJPCCrvisUpvNoNVyHYzBT2aDFkfkVE4MT6PXN33LF3HBbqrhYk8
r3/30iR5vqliyXG2TdktQhxo3CnaXdZmnPpItoje9JbeX/sx8DwzDyjGVaxgWutrid2O8fwzrpU/
RDUJFNfpRco0kABxlCtrIWSPJvS8rFTJDo+j8mjM2ox9XGFuMIwfAI0jBhrInBgNAZKs+YY951zq
M6uHLIAEAZZ1jBz4zWTZ+ZvbGplHU2qwNln9eK1gXpET1NADrmEErUZSaajJe4GMLtT4Y9kRnrVa
eJxYxO+tW6S4R1J2S0PaDFfPmf4mqyeFdNHrKS9em4wZNyHesolBZLb84PqvC+jplxAbh/OGfQ61
CyqeOWSnedPRZV1FkO/DsmrePQXXZzYa/YSCkOvKyljYjXQxrg0dqeKxzmYdpC3DjOQt9CeEnLqh
NN2dYgc0aXC9SjwJKUuWkvrXYFHciFug3LpMRJU3vEhXiSbBnKQAZstYXAEwGlYK3mZY1lWnJDcJ
C6z6lfIKsdF3MUcXgziC244ba7h9TPPm2DdieXuErMYDR1Zqhk8/tDanWdmEigJnRWzrNbd5AO6r
N9cnwa53FZNA42hK3pWM0rj2rRh2KY4q0MATb2O74vwhDNvIWUKCjO2/5AbakJbEJcpqi5e2GFl+
ufcj4W+SoWjQ8r7CHb9MW4nekREtJmHpi9TkTO3aUZjaBOm6nhO5UtFWPUUw5Jr21Xcx3zTbnqjO
8SR8stkClk9YBf7+Y/VRiTjCii/o+9ZQ3Unw/2KLkjrJFeMtc80yI58ai78mK3CypIUBfHNjRSOv
PA4GjyOPYFL0a2hMPy5PcYstkE+sV/AbBj4rsqqW+qNxffMfySn/WCEfPKHUzEtPUuSZeYMy7u3U
o3UijWV1x4VT4bkPHIRzLNIF3E+UHymZP/u601rWr8c3egKQp4lbFjHK4cCsRA5YRQHuL4z7Uss+
HV0t5XX6ssvEOc6gQG9+EwPSiYjC9221104ex4b/87Ep+m0ZIszOLQphYRggm4R4q7eOWPOovh/Z
JH0CJ6X+9tc06H9HeVYSPE6X8zRwD6Mn4qNiU6xd5WMC0hiS0xax4vv8nADXgqyKyopOvuxp8yC2
x3hde0TYoFAj/6J1rAzXMaydWUEiEmxVH1N7uw7uU7qThvA+UmLDfUlj7izkQrB6pELoYxrnIJ2k
AemREZ2wzzMhDbW/e+WZXRHzUb64+z2xUR7F47iuXIlg+NNad0J3ExfsZWDS9MkQ8bCKGLCxVfU4
CQmnE5gV+NzOLJmmxM+EFVPoFxW6aOgDrPkhsuiTMMglm+jBKVISM4v1HBdapvGp6l/nbCgsWsYY
tFnqsqtKgCXIoYX3xB8WJAivEguPSoWqrQ25enOliAJICwQb8AhgBUWecfypnLuWsqx05dos91Ol
yERWKFJ/8kj3+RjznJI6WI1QZsST6PaR4XOcLGIfTRsbQXBVpIa/6z1q8BESjAm5LtOSxpY1xI0i
9adxXHRdEIzwm5OXtNMNWHmIojsfnUhhKsPHpE0x6YkGHuNz+VE5lRiEe660WsXtFvqDQ6JlLQuw
4irNvFLSch2qe4gvNG7HD35X2bgS7yUVx3zdmb3RcAbYdjlVi7SsSJBK1gx30vJmT+BjgJ4yxsGe
i4rS4LAVdoRfsYyUBGzWq2R1Yefavxq+jXQyofflZVNUEcc4sxB7E4XN+kqpjcfGXmZ5S9mhniWu
EvjE1DjAYjR7dOQkESzLEcs+fpq3jh7GW3r3NInohEMYoqyGm9oG5RIvGV+ArGN9Xilc7vnpA+Sh
GRXN731MeaWqwxMxv2F83PHOVw5Q7SKM4MTjZAoBrbOGIDj41tGgDS2n/BooQ1jpl5mpPAgfIz9v
0cKB7Ozak/JC+PpJuVTY6vK6Xmte5zilFpC2tUAisGlb0l7fk1Dh++J6fhXuYQeV3sWNFSZFnThC
aN1fnD2txnqgaWauJAXnmxSpMNvuEnNlpS70IGg06XuX7fE27Dh3whJ7Ml8LqhZmHOBQjyBS5h/G
xmSixLIgZE7JLNAk3sPdpDdnOcMvY/CjJj8041NZCgbspmuZDxyCpJlaHgVBrHy+RxPbKdKFmiRR
ubxdecHK6Q6KxM1XfeNFTHV/F2pyODxp98BNW+f7CZJzHDLQ0IxKGGdsu3SmIVKa1LTmwrfQvL3b
rRtUP5wU1toRcc2Yr/MqcoOrFfe/GtwK12WMHMue4gIj/vqsJaW0Vci+HvNck3UMajAa9IDoBcuM
PzB05EieJRlxilX/AMhK4K5Gi3379Cs3dlMmM0q5xSaUdIDzeufzF9P+0YAoYg/rcb5ykwKpxATi
SMtH2zNb4FXCKzc3CfRTJkGR433cOoyHcZwrJDS9TnMk4sshHrWlUVMnhDgPSv7gDVv15v3AvNhc
Ge07NELDTLyGvqYhX+Ddo/Cin9bMhG9N/30Jb8zG+YsCnEYPNYDgJcrctlSe091CIyuX/u3T+zi5
unYuD406k9oR2liFBxjFrf+a3C/7t++9pFtPO1tDfIYJBOq+/6efFC1sOrYcIP2lpI0ogQcR7X6o
KjeA9QVqpp3pJ1pqDy4m5MzBTt1RweqcTIgeGfce+dSXJRx/Mf+DqQ/eZLcGW/y5CDu+tWQSlW1W
mAYlTrmb5Zir5+QqOJiqLxHqH0OvVq6B+BUeRe3UH/96KicB+E0oumwjzNN93V6EyTsO8Fp5RrZI
z8ywGXzZK+Tf7lNpTM6N4bY2aUjmk0ASL2mXgoVdOhXazyKz3y3vut1dNAGdzW4dsymq7jr9AhKv
j6aRIfBNzdPvLBlZOnsW7m6DQJAVApeWy1ZkBxx1frhlzTZSf9DO1UO3fKsl2UX9enLuPx2DaK8i
SKEj+DW6DCEnmInyikx/wjThrcJ5CaH33TfkUNMbpSXeWv25hUwtOIK627I6hbAxoX576QHgYu/6
h/h2uilWL+J+6UPswKJAfClT91BKSuviuV0faHYY87Nvt1TezhwSgbZZNS3det+9BhlqkI+g6kIw
zgRmh5KDY6NZYAlf2hwnI0lzkitJIZDCYExCDaILuCBEXSuKkcyckEbtGKfDNft6OPgGW8s0W8Nc
wlVjLyHbh0fvPoPOKu+ruMk/gjV4/eJlZAgpftqCtlu1+cun9n/Wv36/xiSE44G557AtK4wMvOoy
r3kX8gmvDatTB2nSOyTAQlsBRnniTHDYk+AWr63WXHkJ+z4J0DciBuIHEZIY5m0Bd8o+t5Gxrdax
Yw3r5ForU5XKcqzLOhbI987tohupMKC+n8tQfrJiIPJpGbukGiOEgu0rwY59EGprURShSSYv/ill
zHlLVRsuLw7DWlc0lpBpdXD7vbZX7AZ6ttSbpz5kOe620K9zTmbxZegOTn2gzm257JnsYSzpatI9
9yQiXiw19Z3BW3jYKnhuaUkpGSp0veGe3/zYNa0ey9e/MLiFbzdvWXI2IruOdOXkyuJlLeI9qKS1
2uyaSL3G8IWAeUhlpx/4OcM9efpt/SHrXKm6beKyCbm5xaHCC3nmHwRPUJ0TIKa/86NKewgbJWhe
sMqqTjxehhjAIR9hR7ad9fgT5POxqOvkrOWS/sM69ZALzaTkHEr3rZt3tdJyCocHr5ogtuSdl6yr
+v8yU0/OpjcmfapKHGZNH8NnZui9Tl0vHQQdsuVsNrRMUQnNDTDM0wNgw03BSXqVkwd9iTsxQW+m
f6FpRnSma6CXKcKHXsudvZGvpg9o+ysGJ74QRm+AZhnhD1a+x0Hcj6O0cvjH7Q+Y/wBzspdiAoNG
aKytvh2qsvcUElhIm4Vfe4e9Wae3TRg4BCHXuT9/Hl2DVTHMgEfOVCQ3/btrzhYgqWG/Ec/BbqVj
MGt7wzyQjEkgOAIxEc4dZ6Jbm9Q7tqMk9w2P2XLe/OH9p0UayyhWnCjf6H8VcSo1Y/19QkfIF48H
eAi4aPCEQ6HuNkKcRAnbQ/yh1P7YtJk/0E3dxWbSQX8J8/1rYP/b5sxOrA3SwLsVdwSH2rwAgpj6
S3qANAKod3TlTpiiZA8gKBiVkFSl0/I0iwgZuR26H0ZoL0IvLdmB1hU1GGoGVPBPFeP6KV8RqKLk
e6J9LzB4lVxsa179Cx6q+WxOOy1uNBP+qAJ00Ag5JWU4GE8oj5/FmCQsYzcwMfu+ld69861LCOo2
Hf3ibR156/sEROaXZ5ZP0byDBU9D2gvAJX8/TJIWXi1PYGLNSOh20sk41D6jMIUUPl7tr/lgE4oc
Sw+2ExIP/peLRu6FWZ+7rD9AuhPPtRAN2y4Myf5owSEl89sjVnQabdNW4PuOWEYfNU3ZNsjNOT2J
2TSuNfLBz9fC/xSk9N7f1DkUZkbitpJVap4Fzj9KFZUsn4Z8eBvV2PHISZU8hjNIwdHB37JO48jZ
cjsV3TaRi96VpXEH9TSU1oetYMs1dKRB2ctbYQ0bN1RjUFJXoUbCakaHslqnhkxT3XnMadbGIr38
drGEyFdIG7mX+k2DMbYL3ZkSnRv5LefUf6PMW7ZLY/0C35gQ5gSE0AT7uznJ3ZDK2zb40IPecXu0
NbRA7LSNHPnaUd+OIgTxuJhKbWRtWwn01Syn7tQ30ghyiJnIoATwUncwXSM9bBn7ctvvJdOSPK5s
JVwAuwWhYNd6UqCB8kc7EuT+DUWKovNAQ91gaCmVQXogmTn5Rucetih1v/OI/XDRAElHtG2oQ0Rq
B41sRKN0POvoesskb8DiYpbXL79HKUnq4UUMArvNz/WKnCI72sZshXQvd8j6wyWmIEQzPwBu3+67
Y6AaNmy0CFA5S+JkEPK1tazFOyAVA2kHroAuAYFkXhkJOwd4rIxo3NjlcaNDF4tcsYliUEpP/xI2
idQHEjB9wDtdjrbFOAjVtWGLvoLZHw/K6zdVmufUwzW2S2WoUqsh8IFkAYVHzS8suA67uxn6APRF
1u7zXLRbd+PdS4XOEsRReNd63+F1dyJj7zUpa1CsUXMQm0f3GSPFEK6+pNZEVY36BXs4GsHpZysz
DXpErlR1csa4p4P2Kxwv6riGhnVm3MGnWftlNwnglo3xeEa/cPnIEPZ0uj7O9mm9ImhGldQVqniE
g7JSluHr2RD9S3CDoWZZMXte1UI5p99G5oYuQ/UrBJly2+SuuGG7oCyLIPJyluLHx47mwPG83ytx
O2oG1LfOdW76cP+kEJBpYm4Q8yyWKfZPdL3am9SW4FmttXv7ro7gdydT3WH33rG3SP4jeyG5TB1c
MXzyYYPX1NpkFAvrOb6AU5iGUZgwY7W4n85zPAaOjEWazQX/kfDRtqwP1Eb209eqc8iqISnFQX66
GSxq+mmrZBh60h3HsMjd/pB/LvgPT2PjrL2tWZhxjfoFHWiIrvvaNrKJ8Wee/GNWh6CrPKxlvNdH
3C4vmUS8vO+ylVTo5GWU2DdJFz5SLJuBHeBl3oORakghDBViHBdy7bpFO4QniktwpK0tgsVjbBmx
c9CP8rN11DOy0KJlTCfct/PBNRATTXmgkB2a3T6IfFxpAyYAZfT/WcPWiCKjAfRtzj/J+sQp1Ui3
mJMVzYNro7IRNjXHjW0QToUmKwEiZrka9M3eNiSIdad25dwN6Ln/kl6baKCiHFAUW0qL8CJri21V
2vvMmNU6+PEpRy4haHk54bESBA5d7uqLskTJz90z1Te6+0VgVfLbTcSOVHRxiXPS12+Fq4aCj0tV
EHnMSPhrf9z1cCbwsX9QXBU6ofpbHyYXxbSnatbzlbHPYGLVUdJbGNo6O9L1zhDzh5IC0hMLWtcV
bhGCmZJ6nTnZW+MdnrEKABEXt8zyLn60Ir0DD5FpQ+sNgHalr0Gcrl0UiIG+D0HvJXPbAcmm3NrX
PMQvwRxJDERbLqa1BN5imMfzL95T4fdX5m+5IdZlBmEX6volLDKwGl5iNAt2CSyzuKAcIe+Gjh6g
zsymaoxpmUR6SXZulkXUdLOjl6qgwYkMDez9wWSpGDm7BVABplhBCSCaH1XxniBZcI0Jz5BMmmJQ
v+Yb8Uk5UhFOdFwb5TRErtP+3iuugTrGtMhb1vLwzC2hgaUta9aHzMgGhDvn/beq1JzlSZG3aXnf
xY2GzbqHO1wEQ5i6iPSNnDbc23EBGpEfzEhz+6Xr1l53UVa3EmVvRd2qSBUrvAHHV2rVv5mysPUQ
KVfpaZo2X8BoKCRzGwSgsDx7JR8qNbhboRuBeX7bNS+EtyOzIveJswxDFnoyjs4ez4AV3GPs4sUd
9dku82lkTSUDmO4vNbCYKjYLlNrcO+WPioVy/sAZB1/RAUxcGcorp97DL+hsa+8LqNt1Uf1OXCHh
wB8dewv++vD3MtizklqmahKyPeOhxIOjSMxBRORag3yhcObjeZdmPk3aYXUqOtOOz7k1JcPnnrXN
M7vBNxQ+CbLEDKmxXK07FIBdWnW4I84N9uWZgp6+Grsx4jMvb8pffUklk+4s+3W28hL/Td+8j1Jv
h5LEPkpKjtbm7/sukZTvjzgERnKyFOs0uk6RzR/5tYPfBPlCVUj3/eE2aag5TwxlNRXqjraoGkQ6
eXxrsI29XoNfTurZ53Gb6dEhRVhyAYnSIR1NpUbySBNl6393SQJLyLuyJrZSLdWN0gEHt5prurKO
4FIWrkDy557IEP3WSwH0I1vEKDgw64ahtr5CcXAJL1eQlY5L3BItiq2ffCWqnjK/DFr7tGJNdir5
ZXzAUlv+D8WdYeQQf5bJ2xNIAS6b8mgZGy4yYInDReT3QxF/nUn0c1uCswE2pQ/1IHL0pXny75LI
faLYuAD7/X3t6qy0VeqePpI/ULQFdz2YlH79ueGgCNrWEcM39BAR2+TtyZMFLAWJ+nsCY2S/Lskg
tFrfpc2rGk0rWKjENS9ohc4tS9Qc2Ur6C6RJVFIw0nrOCOVmzXCSPw+t/G5SOEGU2kc1YAXUd2zo
344FNFc3ITuTADvNCMAhwVin84L0vWC5NjmzRdfwtHN+8g/lJ42gZD+xTLwUMRNzNemyE5aIZycb
uTXHWrUT/OdKya3uxfs0hLK33Bbuu0E2cvjWegPxLOxIv3+JUUMTiI3BfyG3GgpbJmRIcFibvZlD
M7+a1vKWOvzaLm5CFL3LGee8IAbZnmHz9pWjyHTQprP128CP/Vk7iRG9vakaBwsR4bKkiTd9hc0Q
tCN3IYyNIDLSBdtIza7Co7N23PHdk+bOIl5jgUSGMlZVrGQs/mZGQx5TIe/4sxCRUvKWE5sCc3E0
AtuX8hC9o9oOBBigvdtYhvjtUZPga6nq3EYTuZks2yS1RpWPNj6jcrRhy39rokHqh29yCput8JQy
ohtrs86odhO8oQmngdwa06uKYYmpOiKjchZqbAp494ESOVPIFld3fmvz5kQt1j3rIynhGPEMpAaY
8TVqIsZ5O0u+QjiIno0MXW+ebzeBNNNUESln7CH2j3iUE+k17j+256OgdiVjzIVCrqA0gmieTmdY
5yrSwngqu+FpxK4ptwrff/ZBv0U/exCH9x+ZF66FWEPxAufrbW+4lq2HfGcIQcg2YmII8SMoil61
f6OjsynyILJM0tJbEZ8j0lf/VVfSIlDAKKRDU8aC+mqzuemWNDTb7W54ttOjODCv0tsU4m9xWxv5
RDm5UvLhUNBOVRyCjb25Y90IRv+WDLz7/uIUPU+zd1jGKoVwJZLpy1HfzjxGUkJBpwk7UOBHJjeZ
MadKV3OH+8CiWPBRY1H5LyY04kf6Lapgz1nbl7H1LCOZR5Q/T5dNn2aCCvmRN1w5XJJzwqr41KI+
0PbBLEn6oi3BJZJW2XucoiGc04uPc2oh1GJ/FIaKNQnrFf8ry4/QhAfKqmqsl7uT8h1/W/tnDxsw
nWkapwCEZoi1TL2Bs1nYYV5F2Bp3ZhZdV4gOUIoiGHpLatlcjCNNZ40cpKdwhhM4yDuZaKRPR1en
ETeODZq1SJP6ucWNuka/rNsMSDW07OoUtsfzUKQT2LaXl1CTy/5ORbARdOKDuQjsl2vIdq8Vstgr
fN5V5vGX8bk9n09tCpuXjs5Lhs5rJHOefyXnCZrXOMq76piGjzH+MJal1Cg0mobHHwp8q3rszVuM
seMuLPR3EUSLpcGIAyNN/5p2KSghFKYOry2oqXJ3JNaUstpmHQve+o+KffT32UEdtMC8O5+MEsjF
OVP0Wf1sEEummtUXek7pc0e1RKAdjhAEj1fuW0ACLluCuoqJBMnCoF+RwC5e2EcRfytY4MS5mYGx
fVZoSrcN30CAxk4kEYQgbNYDo2fBtUQn07OEhaiMT+P3D55lzVg28CkqS5gDgA+SMEBZo3LIgyq9
nfRPcWCchFCZInndzzoSCYp3PUOsiOXlqKFx6RoczoSOlLBPGhAjljLg6XAmGKZgXBeEYZq495Nn
vsbnnWacJiBFVcGTe5JjsyK//dkljP5PbrntYTQoGCN/b/4WPopqRWuLrXxk9ds1cxilptiYe6zd
vF9Sa/nZZsc3gf8+gJvp7a9gELgJe3TN9liiwuKLVqOCvwdO7KTcACtwKOfuOxUI6/4+MUXd4qFW
qoy2bNB8BK3EkIqoapVZZkA6Wy+Xz9w1wQgVllZsgR3dB22vrha4cLFoftl9zuTN8Yqf/pIwfOgi
c0DTQvTBEoDxutopd1JyDrzOKT5Ks0voPqFA1q2Hm0TLTfB61IKUOiZ8/5mpfGTkuwOaRrHFtMjR
ClAMvPmFGfcwVfApNMJUvUIHlYQf+LFn4lVO+WhYobeOpEr8TMBZ3mUZPeeT3jjo6b94rdSPhbvi
I1SEQmYULrqvNt1G+/zJGvtDP9mFNw3M7CQTz2YIPSIqUzuIvD+TirkGBDEuEkhmy5Yp/rUNoGjp
H59/r+GVwtXGPANIkxWptF5YW3lOZgavXlJIz3TtTT31OOsl3JgAp/pTwIW562mw9XPUuNLJ2yRa
bqCrYbpmePs9vwjCBVi+iHGrjjHr30a7Oy2261XDwqQGf5zvfpX664hA5OaJxfMME8eiJvJgmNsn
jnnPuPPT+rMOAKu84+qks5YZzSPEUS5s6BYlM0Q87T9oOjqvMgeqKCQcSKLYRne4/kB+mBSAo9YB
nfaazuXJPeuq7NO+VJbp6xEyIKKme0p/EpoavzNoM9ofOet+8UBE1xP6Qyid4gKhwXg3ykiq4BLX
b+GKMzYLNGvlSq0pyUg+ZF4C6L2FYO9RHPiPQeqnioGo+/nShqx/cgFeTaU8YvsZD+6X6TPbGFhM
Ffdu5jMSO4de+Cae+puWfKzmzUjvqBmMqnu1jC48owcYzczTX9NLaPdebQz4QFinLz9yf9RmFCPg
pTMyRrpyZBIRQ54dZZ2+0wx/wMEawlHyWy9HQkOfXzXgB1lWvaHclJKdu0oIiud+ZtccnAvZ8D4x
jCB0GLW3ZUKrASH8A/jZXxYK//OG0arpzmiGczBSB9+odL1yYfDginv0N9qyM4Iz+W2jLR+REtNR
vSKBV+xkYhbXvEh4Hi7G3I/+9NKjG9TPCsXLw6qXCM4STSSuAv5WCKGKfUa08sdS/YDhEn6v92qi
J6M0EJc75Y8xukP9kJNCrODi++6vChsjk+1ktDA9mDSt3GRdiYZt/gw7fSLHWw42AqCrCSMDoT/d
bk7dHT5Qx/1N/eOfQJD3LDgXCdZUanOTFkTOXLzjOtMlI1FTlRs72pt9iGeDPH1uchq1veKTj0FQ
NEZ6dzM1YAvT5RS0fhV7NbBlxMOruarpP4rqCOASRn/UztqbzqoEaV+oDYdNrK6b+JSBm+qWC0Cr
sVa/ydlLiazZw7cz8s2ZdljocuWNX1wykb56AILEcSaK4D6E/5E0ySkSdYoNkQi4qbBVdd6FMaDS
uCsM8EgHP9K+SiXvmwXX6pyEybRKq5hKuLaP4ABPiILKtrhbNQxiBNW6Cs+4qG6K+zdzg/MGQVU/
kwvy8z6WRuHpQj3Q+PBCWx7+fif+PmGi2IU7j/KfIcyNhG5gjewyVS7cEQAT701vTX4hu0iR7rnO
WbzVPR87tkcBYhX4NmJYqwpDN85Glpdlz64tYLL9JFWIouf1SYZ+WxQL+Zyo1aGxMj3xwrsAPOMR
KChPFb0b6r3Xh2uz/BckvSMWl44RVQZWDQ3T7hZKEiH7DRAYFXQNnZ5/fCwWibPijohBi3v+W6Qc
4CZHx1ZXyqcWgMOCTSetcUSYvp8kdjDp06mIO83YQU6HNdsvg75mPp44oLTtmChloDjuRQa7t0vd
cjdSXbNUxLLQNhC5RsHyL+Gs15vl336C5aVwV3fqWiLAJCkjR2sjLZPTnWtrgNUGxgjXjGrSiGY/
cgURvSZUzcIamIwEqYQpEJuuX4S5wH3eNh9g3ktvDD/IEyH7Qsk1GizlXKL8ytmrL8W5tKcW59Z2
9s+mWMqfT7Nj9djquxm+vmaDXPVV4y8GsR9YK4X4+rJ/DBtPR7ukIOc8UI/7tylO+7YkIpSEQklb
3EGQ+NC+ZtA5wK8a/TRXrY0kPIJdWUPc8wUTm+eK0YvUtXBaabUJz5oWjPp7HaCVseWcOwLVwknD
QfgIR+fe6GnGQaJaACyh1HWj3uL5PVz8ZszENnfxcV5d0RXQgX9KaI6jWw1ap2AXON+mc4VteiL0
jrx2NKxHrEccvXP0pcvqsxX+yuvw3pUp1PpJqjhvmeaLQ26/HdtLrpyjPyiSq0lmMBvBHHbfFp87
fXa12v3BTYA9gvq4hRg6i0ORxjgTdP9QkjPTujyQjqNAFMZnIAEX1ryjRtd2vTnR6RTQFJlboA/M
IV+2lhZzDF5rrfeUVR0G+4w95/sLN+stDhtxLOw1n6a6GFObTRREjsJHJMQHy64gUAGwv9g5HEzZ
gC00eqykrsshNuDg/55mrrA3UwTI2MTAIdaXNqtbvZCosqXzqSAs98LIadAEG5i7bB2lmd5ru3tM
o1ifSCYO+K95zplcV3RreYSbLHkoNkEVZE9XfUgpWFW+xTknFehkYPCIcj/4TNQwp5qYHiU00gpn
UBncGGT9nnF+PtOFpT/TPLAh9QcuQ8E/kraZ8TI3P/BC6Nq/6xTgz6VNlJkSJhk3h8rm2ZjLjbcA
To4deLWz36Hkjk3jkrCIcRY13nYVDgMBZmQQbDftLFOVz0mqFjf9AUiA3lsWwt1o9lgKppBCEk3K
/VvHE1nMCeglYlZdpdM/TI9k/hAut/QZzvERELIqpflSkFi6PENIPtSdWaMxEfTZN0bwlEahtzlR
+X9xXPqQtnWJpyZvmcMhVZbQjAalOn5P++KCvMFKIFnMdmlWC+uDr6Kn9OwZvd8jAdBYYXzw/qFo
/99T6QFWSJmqHW6BptlE6Fo1yYsAUICDJANkRsZdr69PRi1Kp2txxhkBN51dEpgvGM0+Qqwhs5EY
B4I8GXgGKECVW5u/Yqn09aUN6AolBdfAbHaHIXtgtMXsevauWEdpOqbj9/i/k2QARhG8eKDWo2oB
cAzuwMIlTafZDaB6vpxXgArsFOaYvrudY5ZdPbw3gWUiEq0+HV8SjsdXF9tFi41CtG38l5ra716L
uS9qH9bFnVyiAKZYIDgZ5rewKibXMF9q2R36BbY+HF7MgZBCl7RntUkDXqqjRfJ3gy18BzIdnssw
0QdgRu57Ni1zcFv/z4mobys4nYO/436RBCh1XlGHqEYflxzYVbLubuamkOToQ0zUDEtrQSw6F/BZ
a1+kqeGWWa+bf5HHuavnsdKx6ctAvbHJOvEDJx+wM1R3anwqeImt4nTAa7j3W58W75q2neYof5UD
/K1NsiAmLWp3aN1vSpreYstWyNtgXkzpduGVB1UJgupRwOKyKLqJEQ1bpSyKgNfrkEnVlHwha8a9
QayWahl0QmLmHCaiZ6lmHPqqeCPjh2zDHTrWdpEyCvZ8shrdYQ8eYHtw1y3m9h85BaCKsJuSU6l7
NS1hKvsuAR0WKd7crJWJ9x1yfTKNSCAPu+eP00aC6Fi9aM15xILF8bp0Id0mkzzQo6kAgA2usa1H
KX0SekjZDGNGFKZIV4PwHJ9aYharyPMJRVuT9fQwtI+VyuDnF+kApd5TOx/rE9v8+TMNXbRsN6ht
xHZ2W/5LxDeirMKmG9j8ZimmRbJCFwXuHZ07S2dsvlTATr+nVip+Hdx0W79IWk1uTGFr1WFKYGAg
aT6DSVNUv2K4PNnUni5/5BXOur38LgvigAZlMghLnameSDNIUFe0ZFfpVU4rjpAKzNTbIoFbYtwl
beCnMPCkakZd8Qe+D0s/ypEsntzIZFt42y/kjxEbTz1h0EiOefyh5AqR7fGfPCYU4qYcIMVx6eOy
rVwMpKVKTdZgyxNEtP+3Vb3T/hriyEOAa5ctcBRdcejWi7klTP3bnT6oEwHXT+WxZfsYtMxVDWqn
oXHAsCsZBbk0kKiKVb2S+F8wBgYCtGqOhtj00tiZAKz6bFekC029r/KrMhUvcWKk6DfaBLatLEdy
utgSuMDWmTvOFfTRaDQhxg0PCIlrXIljE0Jl7k46a3m/kLxRCsAVkHX3yAvNCLZKuk+FrVXTkm7o
XLUkWjljFJuX910hSswDJZlHKeLZ6scYYs8cknAWSeAPvM8F83dUTYsCKBRWjuvhrR0EEAbxrksT
Czy4RiAQkjDGIRZu7T7chSUyoCcXIsib1wQfK74blVNUIXAfsxteHswgY60ATlXCp6+NTOerQm1G
XdXJ/AuWB0jbKEtB9QyEWIEu2eU4xMlZUVL7gfSMWzyxM7ufdGAiuOstMhSKHM8djNAJOhTnOJW5
hQpH8HOiTFmpXV6dFj+Dt4SDhTFuyHOBkvYj6kMe9XtraZ+piOQZZbs7H07MBE8k9ANWgcFhpi6A
LKIVl4EyqFyq6oqa/CO5ZzaEUo4w3IzbSFEjh69xcGO4Ghc33x15PqiLDA1GptSdN8z5NOvZjpgP
+m16i2U9McLeuBVvpt61Yj6H+zovrpplQ5B6VEKd0d/K2S/C46dXciDzZO7lxDp7cguoO+S8r5nc
RJd4dz5gSjp+zCg9hmnzofGaQK9cMeujJb18XQS7Vpl6X2PToti4/B5LdHStJFU47cQvG+/rzWw4
73B0gRhZylly/jYz+n9eSYiluML3FhGzW4Da3wU6GbUNz1fBzeMQH0myU9GJtsOm9Q6r5XEXxGAN
sbmBnHW/mwfO3Ry2Pt1ByAums65Tv24tvoZ3F2LU9lmZkN027hUzlTVtAE/AVjbg22Gjs0vpPsfh
+ec98KKYP9tHyYqVAjyavj7hFx5nhsHQhOx9tHMlbfUEp3xCX0npATUhP3KTNtqGy+BokfVCBceO
jddfazq5quXKDk7uGnVQvzRe7ZS9aDr/Sig+PFjVRJcjV/3Goo7nj4geGHH37af0OzNqN+Py53Lg
SbtSX1Pb7ocstjddel1jA+G5fQKqFTkHCKcljwrM24c9HT8Ei+2BvaV4R/Z5Ec63LXDtunT8Ekc8
GW/YpEJYlAM7skOWGwjQxIriHcolUX34I6Sac4JVremB4WBLNUMsyKZ5iO3WVp8dEJB2UpNVZ5of
iLtNobnFg9mn8KdoNYXYogY0A4gA5YiLTT59ALfXgNEii6Oow0oT/dhH7f3nz9lazCFDm++/lQgd
NydmFyiXN23cA5/eGK2rITpynVZ4b+qIfDB5PRTXF1lXx5GTt8sWtn/3ntdynMrVi1k0yP/OxhwT
9Fg4dzplo9Zkbfbalxj+edZ0R27egYws7xkp5zbyb7Ij3Rh9GaChW4qUoMGdb2WvhG4pH9Zg8axn
u7Y9Au0p/Jf5pQ+bBmdZRfY0NDJ11HLhTRC+0L7Sy8tls0ApJXap4Y4D/NbpW9Plx+gO/FAa9X40
OQjGJsEnw7tCLQIngyKxVoaL/l26I573ofrlegDvVGLybWqDTky69thAMlk+iq7LhvTcROBU95dX
HweFMiLaR+YKoQiYvsTNrMKOiOX8w9UqGG2KzDUA3DNQ8frtSShdnmOVyh9dB/24kNY4fJfXJrlt
+NMXijyTiLOF1XESEzw5LHFIT9AeE53RV9J9fnf925LogFMfgJTCwDLwz78/sYP3CtAfv92VHFTY
vboOjLgtzfmGXz/swmwtgm+pN/g8Nuo0CT7NbYa9z8VjQNtawlhiXjJ5AzrWOZIyReGNkDW9ll7T
qXZGyZNkNzuX4l7o2TbGps7rKX2kHdwtuuX4JPiwXPHDjp8lLgJR8mswgTBHHpRD5FBB9oENuFKj
SaV15iOgMoPz8JmI+2qIxlhF/swxXOV8hcIHs5F4TeRkXgSuoaRFgWdGlTNpEVq70ElUXpGtolH4
xc8KSAdNblu5l1iAqo1mOvy3M1aM/ljknQ7P9SEaLX9t8Tbw8PlC8BUnItDtEnt5jRW+8kHipiWN
iHpYwKSHeOYZ6PW4QY9oTC5QjjpKgXTQwyBzsNclZ3S1F6nCsm4jCIU4E8MR8kVkctAJYgf/y4pF
JJGKRInQrN4PKiCk4JOA3yc6WG1JOyusfVamR1SUEkb5cHHFdUyYefIuwDysosSTt6wfkIpQnrJP
sxohLMA4h3LxXXDdDo7BWVasqTYhftBN1+TRG+RdOV3Ha7CSK9vURNwpPuXsBHYRgZx00c5u3uV0
KrK565HumiwWL9v9KlOcia+Wid7TD/PGYziRHe4zjfZNCgq9Dj8YGQKd3OJoGq/iW3BfKPA65u1C
OfJ0IJt93DbUjctxWKrQ6903NK4ppJpiodAuKcwLeRFVhHVs5xpPA+iygqCtgyVSesTZ1eJic8sb
JXoMj/xu+IogEvQ0qQSFJPPPBvcqkz2vvm0Bg3AP15JY4Bt1L6IHFYLnQHLeQchd0e/iiNlqxpKh
3cqcWBIDrW2MUwZknCG4EmfZEa0kqxoMxg7eOVNVXz2GDhvd3RjukI0fq6KwM5DqMyD36C0MM1eZ
tZnxcdyEJECTAo2Ebrn5aNS3XUfWQkYEVpRP0zbaYFcRz9l6FPojiMzCU8SuppFur5Bio35gZ+Xh
Ih0i8oQ4CrR6Bl4JtC9iKSyCVFFBmc01hT9Cc+fdhoDZ5LmbRhDe5qUaER4R8uXY1uBWbwvgPyeO
UyUT+/RS7F+Vy4YoCYZYtN+HtLTr8h4iq+tm4XI8ajIpRQsZ/TBPWaQNvvNCPdWKQBShwRFEwaD4
GnkrUwlloV5oZs4Y8mmRLeDGRWB/0LeXULxOvySIwP1enDUs867Ku29u+vqw9t29YaxX4pX4g+Eb
TmBuOYaf+jpzT51ZgG+PYOEeK+xFHF2PrcECv8ynN1llyoK3urUOasLQYAz7Yiq8a6NG90G1itTv
B/rpcOHUrcx///TcebX+jz2tO/zlxIFtZjg55MqMUqAlW1upLlsG9et36ho5sJ4246IZniYALg1J
Qw/7WHreVB59pJhv9aKTbpEGeqyis9KB7ftYj0TTFxmp1gpieWY6sukS1E10GF0TOcSGD7Y0DoyP
SlnsZkyJ5Srxrb4Cv1JQvhoiJBpWxQxg8bvjNSjSsTj57jn/6FtpA8sIl1pOVpylV3DsW/Wcoxde
U36AePPLkW/tnzgyAfgkoJSVyuW2lIYwOw+CYe8Y1uferATowjPM71QNx3AOuWk0jNl3d1vCDszP
CpX/eWUNftTJSGQ0xUe+R7/pZ9nMIOlP+3d1NrO7+5dAF/nvcYtj+2iGmx8+7RwmEh9dMmc8VxzH
fvb/PgMAP+uOweYPQOVY9HjD0OFg/5cLZ0X68VcYkVAHl91NdHl6NhSn68WFOu26mq/UP8OoIa+1
sP5+t0C4CBKBqfonJ9cBgxP2VSGxIyv7gecCK19QurB/Gd8bHDwISeWywHaDr+fJWG2UgTGim1ml
L2/kmzwAr84J5fFavRaVZN6A2thTkUrv9YtkBOAJfDFbZd0x0IVRElMTutf8ajdtfJTFfoXJrUZ0
hV2ACaWsdWeA03JmHC0Ynyc6vugb96l4D7Kp2XhGoUp1t8VhA7zIiXnOKmoAN+MjNagd3AUf6oYm
6ouKpKBMJalZIMYh16Kze6xpnLbIoQB00y1M48EYowy5FGjf9FS2UPnhHHF/wqUOi2BUud4wK3SJ
ad9llkmdbZ2F+h5TEzz4YkuIU4CRQsT81ORSbKWzNO985kmrjRUmjJA/frM4/P2gdpmpASH8pmaz
CjPT0ZfXWzRAetH9kT7JO9IXeRTe4Ap4P632GN6iAXJ1WLyUpUjSU1vg3EOcqM2ZJwADLutLqHRU
sP406sVabRjLrRbam4FOgTlcv46NkPKHN3Vl5BGkudE1KZKIka0bGBPTqZUVQrxxiTNQtpgo2niL
6ayhS+ZlB+vm+DkueMl9ffNzPnbl9egI3UhJBQgRSGIas1g9gSQ1Dr5LIYWU5OSD8xDqSSA8P6ra
FR0oiCtiduDCNPI6VT/4e/1Oww3Q44M0SP7/78BLh1zUFR0oZD9SPqy0hL7qmNcYOdA1EdFDOUBY
4Xs5cfbAG8oVqIBmAMtceTPepGjXOrgDuMUA3URTrRC/D4Dqa+8yfn4kW6aHFwLlufH4M3V0UVLj
oX1HheDd5+GpbdXIT2kh4WA/3JQ9XNQX+RXFD7lqiLmFC+8WkuWKrm+dmDWpdn+ljfIRi3usCBNM
ngSelQRDk6xFHjGWvx/6Cu6RRcJKuGCqNClIY3vXC965o1iYmVAbgClYVEY/2EYcF1aYuig74o2/
CGOQNtjpK4Ye8PNkalZPqTvxOAuoelyzWHJykgW6lbEOHfzSmlaml1d8Iu2266LABRW7uG8lfSRF
qt1x3lHzW4DTTBZRKCMHW5LXyaNobNHxbeULqX6iqORiIf9HMFF9aE3b5C6JDlFuHHvMacllq3CE
+BCP03K4+weze/NNu0IBCTEFKHt2W+GiBRwgXSs5vQqyjl55yof22drcaR9Vyp9iC25OAXkPM0E3
f7JEUZdw6c3AN2PXCcD+v/s6UkFlY4WUDTiyUVcnvNh3VSDZhB+QIv4II7a5zswT5M4U2ZgDMWeb
H8n3OgWzuBDbRwf1cdH+ex53g6TFUfIQxALW6T8D3ixkDyqOHLOD3KFX37DgVA0VYC8qlL1idnYt
YO9Yj2H6jFBa4iuAtmxmuts45SAld1mmZNiALAKRTxx0eMS2qx4iR/7RYK2+OAs56OKU1VKoFRJb
NR1YfhM7OK7ASqHwQB9NAAI9k72yzDrB/3fhlxbUaxf4+zTRNrjFNSrFgTz3ZfmW44l8vXRkq3ER
c9eS/XDkZ0WhflssBbP08hfWawSBtdGj914i0cOt7QEt0JWVyu0TDKBNh1Qu9xQS4tVQ2skc4B0N
Ql4m5x8Fa266W1dDdwH2PKXtkBlQkHQxdOro1H+gQvkHGPsmNUv4KpL3IJFpG3OquHabe1ZJE8NN
eNrz0jAXqV/AwpgjDwu4PpW0Ua8HsULjN7Rso4TwXpKM96H1J7pZyi5ns5PjQMn/3fxgAs+Uncww
3yuCaU0R7BqNvWBMtpldhukplxY/tvCMzdvhbqVTSVrCODXTpEl/e5+OeYyeQU9TlE49aq07Gmso
KWuXc2bKVhojvRLE49M90pxhB7nb6WS+0J6SI9b8IdmlQ+MCPf4NprfiOHzeecNsnOUv2QLW6bAz
/gnIujDd9ugKSLo4afGOMlmuGl/fVvTBscn0vkOvJjzWx7+EOwfQ/wk2KmYeV2eZrPubYeM/x2t1
SevZ7Vhq7BjoH6sa/m893sgnaGhOq/oX8hIwLSkKWtzC8XMEfzHmcfc9neRut62CQrO/smDMZW9r
koTbbjMJGnH/i5fbtNEUB79GXDqf4HHisOqFn3ZKhi8A2DVh1lojw1g8UDdP531qzrEApBYUMd0u
yJNrfw1ti0KNWv5vOZaBmyLjdxBzaHj5nsuvdPqlvmwZVAcY6lY34gxAPfCC4PPkIaxj7DIPMv/P
c7s50i/nb4VbnPB194RfY2tkroerpJaZQWH6bJ1OGH23vuMbXLLOHgktvZDf5VdfAjcgKcRk8QST
TYApEfAqcc2X1t6dZwZ//ZUHRiFdZKU70R++3oRMzwHhxqVx29blr5BCqgckwcDwcI3pUuSK2fqb
PQGWjgm+t0WwDkHABFGCkpeu9kV51Wavk2uutaVlhaJM+XfcMQ423uZFpsvIQrRYuEfiXTxLFzyQ
FHFIpNNcwbbS/36iVBCQKfQEKZmf47cHrTye/mylTWQWUwsW603dufAHZUU4wZFGHhl4SRZngAac
OWT5Sg3BtDXPHQfoo08tXPyXqXU/gn6qLPje3D776yyfoDZ2zhtMNe+u27qfR4qjx7XY6YN8Miro
MeWP/SODamiAmGwoGpB0543VzO7CZzJwznKejS5huhEleZf71oK/s0SA4uwc8b2hzQtITsstV50M
8MOfC7jzePeshesES/GEVKy0H5vdVN85+lB+NJsrxAhUrByHCB1T5XUHPOpbheyRxvl7oxMBD2V3
t6FnwPBoRv9nK/uAYiurwytKqD6dZLYJT+NwcU8HObcd7hX6WW/PL01a+p7FfUFXUfdDzIT3qK/z
qHjtU4F93Ph7BSlS+wYY42ELFzueF9caviVM2FyO6d87fKCeoLKTgUnk//M0NbkREtVhe6/EKkvE
fCPYVU/MHA6WdM4W4z/cKk+4UZg9U7I9JGRnqTT0IWHv0ku/PMn94QyZa8zahnk8yjh9JuZqeM+I
p8Nli/XgXFnjvEEYa6rqu8pkHCyX+2R0Wb67esNv7/RV3cuExHtgVxDOxQUgoahOEyxKCpQvowr2
dZgC6cQmBiqfSTAPazG8/iPU7IsB/9jTfZZpHoK1u/nP7Hr6QKSe9CUVv4yH0PpDhZhWQupLrRNh
KiLy2eBJ+bfMxhBXOtkxXOF/4lYKL2XDFz0PIQyve8cQkXwhnqfbSBlWlrBhmbbPwE5EaT3zveyj
gLsYU5739CVm7c0Oqlk8kmPLiQEog4PvvJ/d5V8AdkMd8CAsXAWxg+nS/diTQbUl0eYzzawad9MU
4L0yBiFG321Mh4WiyLd2ItbvP3OwZgAk8cXK75ESKj7CIcCikTcXFUTQbQcQW8/X59L5lCTj9iCZ
OqH6B1ADfiIbq+W5BvDMA9ll0GNtCEBlxBA/9bQkVGNAAUyVbpljLmvJpxXJdwMChEFFYiRbCUFj
s2TV1x3g88MZ0VRa55mUh3g+xRusXi2KEpJd5vjnZf0K65KOADupNbq8HbblR5P7SAuA35kz8g4i
R42vukL0ySa2K2omMbGmJbf+yEPJYCgYHwpIMB0vJqnMhOesKIHvfGS1KTpmEwe1zIdMLHWYydbe
KRxZHlCcy3wiORIitXktnQfArb5HG/MCD4EAYNxZu0Y8eKoyzvIg5rGLnfNERHSg82jJ/q3PBg94
kfh+ZacmgnmmrmL96K6jfsDunMdZGzcCcZD6Ks82YSxXWCVGu8KLaTCXxUDgUpl3ywCuWAkx74W0
UVAJNpmsbcwJz1DVgIonZy/4QYQeWc1No/o8HdHuuuwNQtbOqsqYIIDCycrInZ6KIUauoGvqDcrc
cMAvFMpHMz9W/Wol17DO5EFsKeo7KElLATAis7E97sputm1MGALPWkmp4adeQBbyk4wv+v9TujTz
kVX+JMJTI3EYeynyuTiuyJISAQGf0ys7ty2qNsIMjJ8nVVAlTcEvauHQkcByy/vSt05N0JXR4YrH
M5pdIWtv+O3JD1TL/xY0Wpxq+5HBMWpjovEacdX23FWMsG/1TmmcJb016ef0AsvF04gb/XsVlPSn
QnT/rgIJ3WhvjlXzoQJWtK7urNNMnxdwYQpmMsX3MQVeHbtasBVsmijcuxHPx7BFD7iAkoE/TMhV
jYc/PG4USo7BoA+iwLvG5CdmNcWRXl0A1TAG+s7fMEkpKzeLCz5AO0O9cY4iz32/tCh+Jr+byUck
xfkPnbCTz5mlOBjKgK/d2yUzGD9mgKyKeHb8szovNwMVw5WuwcPSnPBF8TxZmOCtTjexLzV7SApC
G8ptQrd5YRuzrVBxfwJKypqfJOB/Y+1d1dyDq8l+mYhPIyeSFtU3p6YLuMlqQE1FBC911S0/Isjm
bJ1eyoTYcdMAoR/pvAY0zPQxKY5t5Q36KeHUrBztQqPrA5vu6m59MChJfpsVkkCggFLxyBjCKyQA
Qpmqe/FaWH2lavHfrhcASihn5+8NEY8IPC1IhmzqsfpKufuYrMXjZW/Of9j6AKYSYunbcCXyVqEO
9ihhtkWwjkBCF/+99BQ5OIJOejNlRLBqg4pqcb9IMgvEyShfEG3K2Jz2IZxFubFVAL+wSsMzlpwe
VN8mOoD2nlyk5i0ucvShhWrYvS8yBD960PXCWjiMi0PNCbU5bqnVt1WcH+ESmcs2yCeZhnUG0Icv
BTs8Tv40Trbo5/M4XFagkwLCQ/ZFacciXNcyg86PMPtDuKfIthUpJdrTeOB9+sXV721s8TB/WyhX
aoQEp6hQhyXZ7Q0Rbhbv+ZcHd1WBRCjqYKWvlJPDxgaqcMLnhc1sVz8HNBDpHQ64DopDm4Yatkw/
hrPCv8Zn7tzOpMJ/W6XzFoIPphutifc3txtDOTcuSpIj5TMiPOiO/RV45jbzNC6WXV0nAXVFJFdu
H5uFgJcvs+wFUjgrMWcitX7cWvgW46+tMtk2NwDMmby+4KgwF5bD8ryd9MkUrgL4Ke58r4NZpQFM
zlEQBFpIqBYb4laDhkT4zD0gxq/AICVrHQMK6Ik9WzWw5xDsTRvd8qxm6Qcok9tQuE2yzQr12A7j
q+Iu2D2exShEpnhJRWHtXFCOI8VveUyOmPYtso1rr7vOWncl2MtI5hllrcQcPT1pojuQ1uQb7duw
ptO/fnV715qcoBPUsrmHAcOCEwjTRoUIQhQHnXEh6YLfK4j/LQluLqONfgVdZ4FahJCHBqQ7c1/6
DOop4W42MwerUEX0G8WCHvGM+F27uCR04bEiIztg9O9fkmKZ54l+3AcpKnqv8RO+ZWPn7uPUzjq4
6NKzzCw/AsVAQtprQJwvNPPBv4oP3o27+7X9IaeLO8AwRmzsq5nB45RH0IkaK+r17C7aVv7yh2cx
pFCwUpFkKt7ka6oOYiEWvm30SN0XJE/FgOHs0ASn+cNTjpbEun9UGfO52VLRbJGNK3MgJdEWVY/U
sbIlEFheuE31qwNr6/H2MNseyEWFvm5eDgw5eUaTBYENvXHbBj2TbvO/bBkwYJ67kRbM9E59QQo3
hRkgWYCaQNXxvHwihYrGd59JTcSUVc/CbtB7aCA1CSW5XrVlQNf4+Uw9Ylb7HI0QKmtIzb6nT/eQ
zXJWxW/OnZ9neZ67wgtSfYGhEquiKehpr/snLtDWQg9pXPwCcyADm05Gumu3YGQp/VemCobPBG3D
rXTNBAMbyeE57gRGWsP2nu9u2OgujL9kxy5NJcHwL7kEzMptEfwf51AIhnUSYi2XCpbZrDeYPS/A
rsvCsn/B2zcHdYkXP2jXxCpR4iCa+BrYlzo56OZWduCsTqCNqPTHlIOXezMRo4JzScTmperoUsEQ
Uhq3dUjYa++FvSIGvj6P6XNARtT/8selCouXUKT8X66x5Z2tvjpVpo9/utQngz/HJnWyhecGSGtV
5cgCxx5kaQkmerJZ7cfuSqyrYZR/a+JS2Gs3Pmc9DemGYRbpW2TXwUn8J/eOLPz30vyVkYfsj0RY
SPsylZmjKOJoRm/4GSIZasKJm+LPSDFcGw13IYdy7rArx7SSBbjCHPAClax3TWzJg0e4DXdUt2hj
oSZeA8DQzJAGjIu5aNh7A1KhBiOPdDSsPCsbr40NXbZdP0C8gS743zgpJuqlJkKHiPScOFOeKkao
FVJ264YttN9yuKllRNrqc2cfudEU9q4QeSmgz9xilohB6P8l7/1ckwSCRVYIo5lRjGpdpg/xRI3w
Xth5D25RFMAawjHTF1dE+o2Tel2ntx75mKuc+lwkBL+csljxSlTzX6s9ov6F+y8+wnFNtz7iAXAC
vwq3qzpk6LIkCX3wEspUcZDcU7hq6fF/eXpzW46dLTeZOpFqHWHm6eRxnD/hReo4dEbvq+NJ/gZE
JJouVfk1Y4i1qf1U9YQU5rJRI1uCvQeGwaxiUCVDrMfnaU59J4eSfb6MI0hWnszkQsrZ4Jj0V08c
tEr+rCmNgaiAxEVMoR6fjQftNHjw9Ic9HarRi+EspFWq7jVEAQ6TN+PQEJ2LY7NygVLeP1QgpxE1
XmpnuCHnZttEbaJpViW0uXiauutNKzf0jCsBR47UelEeUFlRumwS0uaPjKf+2YrNWltF10t1n6hS
iE2eIYJIyJNx+NDu2juXklEspN6LHvRkno8LfqW1mAnwEFb0Gn82hHxRaYsQJwnUR8XgQUFGLXGV
tI/v+2Te3Y8c39jZv/hTbZQvKbeZHd3OLsVl+V/DUEFtTeLqM+NRu6JoaQCZC3yu+9rT/ClTzW7S
/SEv6H4bvPpdKMK4w8/5YX3FCohF94oL+fPEIW5fRsBZZyzsavprHFcFQY2Atlk5MHfPWtaPltLu
QeKVBkd1f0wRK1tRtdMkielfrSR+BYTpl4Ysn/Lh/h5i/9yK7HKx/Bu33v25WrO0oLVP0SGJfLIx
MSd1IT+cP12fhVnaoWt+rZHOsJJa7SgMP0ssfYp7FHoOUAvhn0Na5zHcIYC2aOJR2Awds+hhN364
lrXAefXw3Mjn6wCIpxJZSak2m6Ju5ZFcea6eayynKp9MAntm1/Eemk5saUmHRHIDbfdL3Gsul7e3
zXrwcmjNpauXgc9We3lSqORjooSbm4U6cMxPfB+X/meLO4oH8kxqxvVRHlAItL1x/Eikwe11EDfL
FoQqbf2udCTasYuQinIGhslKRGhgaTEumPhw7+58JnRXMAiN5td9QM32H2wIE8Xs//j9SDl6RN0X
HGLabm/HHD7juah2nCoLGudOY8z6hgVobuZN3JMCjKbgxphmVzTtr85ESwIsBmhH3xpJ+ZNR7kbF
/u0F2a5uEVLmA3I4dIzcR6ysYAM6SBEbXPo5M3UWCfwUIXaMfKZ+S8pot4X5qO2MRGPfXPQsGZMy
10cA4i+GCpaIQKEtM7PujY5SYqO+lcZ+SS/Mj8jenh3TgXJZDRMMQ117+AA6m9KGFyUZ8FLokirE
4YkgnqwKPcJMKQ923HZsqe7Qub2s0zEVB2/O9brezull6g5uGsP3H7VHklr8YA2/te3x+JQQJwLn
b0w8Fx9a2O4xYqSs11bvit2cP9S238xicHHtMiuENfyC7AQM0ECxrKYYMox19DXg+IfXEWapnYIW
jivxyuVhX088KuG7cJGGi5uSDbCnbZ4+e3lKQ3j2Zm5oaH49RDgFFCCWLQD6zxux+603xr/Tc1Rg
r0eJTINGSBdhjMrpnXrR4Ci6ywvnr4itckexydpkNoikMooVs87LTXOREqiHS3PffBXtrNMArtfQ
MT0/edB5RXwabjkNr/ZO5BI1kZBIM/2qFAVwdm3j37AdEPtvrSneOv1MX1mb9sPpx7ADwr+zWlsK
QXCeUOcxyWMS2d48C1Odz/B7xtFcYxSg5JAJiAZAXw7bs0uvYNSaO6M/v1NqEoEbaFpvB5n4OY0e
rGIZcndrVsai8R9ZyWUIJYP+CbtM2kPD2gB4bsmeV4ELLuGFBCeLCN3oC6t7HxBDTiSPJVGyF7ZQ
Zz+twlzZw6JnZr17Epi1Irf9E/yGDRNIWsJ3PyBb/1pqjFMq9n/9zcxjGWWs8ZiWpSY6dlZb9FBh
KiULfEgCUv9glQVfHi1cy9hRT7Z09/+2GIzkWhpy8nyYaZ1eRO5EyQr+N//VDuSlm2Gmo8VDE/ca
VdSmx/h9Q9bjrHjPtk9+2OI3XhasCG4mOMT1YNHXCj8Fr7lQxKLL5ouvcnSR0A7VW4c3nB+Qa6Oc
hu7eCsZXdJot7KY/TI4JEwT6ZP8gazg+97BlbuSiaNRYNsNxiJI/P1pWdwXXQmocgk5abweqrdD/
AXjmmtcGjsvNUuN27k9lP6keLt7Ja/Xius0hMFVkffP73KghroIKd7OBzNFnk1Wr9ESqflko5QxT
tr3HCnn85JFGw/CmhEVSg2XM316z72w8jaCXTYz+AfUk+57f2d6FvdzaeFDkNysT/ZqHXrX6X2Cm
3aHJsMtVJ9steg/mjkq2is2JIGl2TTZIjzIsUcVBy3g5IZmWy4o8cXcWhVUiNX7x+NOBF7y0aVth
X0P8CsFJgyP8LU7PIhN/vZnQKJdoEmvvlLLu17422Eyc+5iN3V8MsmqOUoEvK/vBCpWXDI6IpLto
HKaGkOzQzdaUMj4wO6zhk3Oadxbv5O7hw/gCbCHtRKoRYaF2wAhT7Ck6tkV1bqg0aUdt5m0q6cQS
VJP7uxQ2aeGDdALghZdbsgI4z9nmZGl27SZ8iyV3ns/lt21OrcsSrnlU0SKRPT31YyxxHHP/R4CR
mB2BmIkDy+UPiAC7LJYou0GNxmTyyqCXNhq5ahFTzU4Z1tJPTVpc7zYXInko8UXOk5anfGO+RnJ1
bg2eviWnAp7YVDCvOY8Q2/XnJ7tDOvW8H5iLxcDqxCZ4QwkugGPaZktDI5hSJSGNCHgD9AvhbgAD
MEjxPYSxPY7qcl1r+JpTJ2RCIZalqiKWTt2xohRc7i1+XKrcLNcvsA1wkibdI3Ne+w8KRP+hZvEW
0WXaXgXy7/LawWpJbkbnmO/xxkwllcjNRZMu+MClXVVliwqbNNb1sgCOjrpuVBAuoPJhyLufANAy
cBzN/qvl1848MEO/mA8r90KnVfEyWZFTZNF9pG04hXWdxbaJjBlPW0kag2O4+a3mKCKb3UZA54BG
smoB3tO8XaCcpbDcW5KlYDiceHpa8zV5zVhLjRYoPgu4woAQAEuQuPzwBBdUOiPIATayyzRyBDY0
5lpWRwgOSoNs5532eiDyc043JTVwbGqcZpf0x7faCu9xdPr+SdXC2yR1y0UxQET9RBovgRcV35SV
f3yF1AhOXG2kZJAHQQNSo211zI/zoOG5FogTIciHtrmrTP2vbMHkY33SrXW1KZewCO9Q+aekSLat
kdWcmlxs5h7zSZ4RzVSeF8OiPZUy+5JYqU9VTYSsOTWCasrqopzjyFZI36W+Ny+3Kg98v35eevfX
P5UHBd3GbHuFTc/BQJXt9xkAp+b81RBLNNa+klnBuDYdTyFq/3Hh1APk768akK26WDD1/m66SbXf
k1U4oCnc49SXK2zneAScwd5DIu5pHcfXdaC28AdCE7wyVKwB8KcJfv2VD5/wT/8+MrPEJcFQKvi1
39yNVgtHcHHMcaqt1VG1LDcgfRH1puh/t5EEmpjKUsDyTwiT5YrebbNNL3Cfxn2R8jLhnbgtooHP
w57762Rwrsd/7YFAND+s3d+l387tnOKrYiMzIexWu/KbCMI5dr5kZ/lAS6INkcQLv6ODvhtPGpWL
PPaE/B1BIWzYc/YQMOgNxFhKzU1+zHx/rKNHs9fWMzJyHtIWhLyYfl7ktGeJ/SVNnrBM9hpLmnh1
qf9ckoJJAUnhXCbOJfJU9J2s9drTaXfeRvaiMGDNDGJkGTvux/wMjP+jHhPGMgtMoIFl10i1acEp
i7YzBTgC+/08HOU4/oa9q8sO6K1Cz1LeSS+FhAvKINriYx2yHrDzfmJH6gE+mpuv6gV7uKTlm4iy
c7rB6Wnb7HByXJlDHPPMJqLqF24qRTdltx4GJaFimPJGqJksfKtr/Zy3178KgYBHchZh28zyrki0
KKEjGj+JZuQpF+l2q6cSw9qXxbqghQw3xe1m8wsfSwjNenVUTYbeeh6SK+JXmoPV9oxr9p/1IQIW
J9fHtm/lAVW1Sd7wZ4P6LOS3w+dS1sBlXGFoG80+nv/e1/0vbNZUESe0A1FGnciKlzCQm2wmAn1v
W14aOfjfbgslM1SkPLFX5Ei716JOtpu9oyfMTNSTrsPsbg5auk7SK4CsI/sm/lZYV1BD/Ncs9JyU
cCSJsTnPv3FYA6t7oGvKI6A6DhcCb4oir4jzs3o3ZKuG/H0UIfUkuQW438IHqAPvW0xofdqqg8SU
OxTU+UH5C1fgqPZvgwAqHLfLXmbpYo0aZJnExJWm4uIwLc8OE3nu0XL1ShLokNDWC95WiWPxF2/H
yMNLfyvotZrIhVWsHYpsmownLqpZbHd6wz9JJ6Ze++830IgHA/OlbrwJ1E4lJTNA8FBbF7OfX2Qe
Y0g0wzVfsT2i74aXENVqCNmEJAcTaLzWeJ9qp0ro5RlPjr8xnMZWGeht5U+2dMPNTUOGBsef8jOp
AaLnpjndryC3dkCTDD9g3ruUQaXEaluQOaqZDz3Oywt3QN21D1Ifnl0YUQKRZDYXh6GqOvJjnVQ+
rMvP6FJ4nkqc+irXBUCvU8dco95GGXfBVpcB1WukaLHxdIk+6rdaJ8iOz8DAYcwpIYKP/Z0Pf48/
2Tg7vDsYg5ur6rjHMhWXT/3mDvPYChudV+rJj72jIWYyUEfLMRG8tEBiPPxCwyGyKc1QdfuOFfxS
Y11gP77zek/62VrUfK0ZVPc38M0xjaB7fIcahgxfTKHK54j+4A4ep7gswfAg5JNkd+TRa/Aw6kAz
JDzq35iBry6YG9vcSiO08g5pfN1zs13s2HqBg3z7AUAVqJJRUCkDUDHq2jcG4mqS1V+BaG+rfHNI
mUfdqHfAhb27zqSU+1tCd54TRRWqc3zRsLrt57LlyM3c1KF6jQ9uLU0cRen1r5JfUT5VrwW74ljj
tDaFm7Qc20PwYQY2VeLD6/DxZCDGz/b312H2bNSxFaVyi81t9/CqfciKiRhZHjvjp5oXk7czLKh/
pUmafyJ4+1gu7KB0L4bgfF0cwn3T5YaAHcGS9jCKiDe3q+cl/xTqHcnNage8uZ30DnYyJJql2IkE
08n2w2BqhkfHH3Qp8oxOeYtjDW30KRzyLHCPrBatT2n3PVjepYhQzVKNqlrhTtpcFs2qkyoYehyV
IghivFLMB49yZ9DUnQJcFVla6NkXqAyuBTmoMw7wOTRt6nq0w5l1SGM9xW/uXjKsv73lwYosRSzz
k4jC0lJqcR+2lhjjmShELEGzeChMx2PWa83HviVYzDnLNBUcMVS35/fl1/RxtIuJ6vmFXMJR6Gnz
V7BXXwmnRBtwiMdiJv5UMZibUvT0/TNkSdJh9AUvy64+iMh6Uzba6ikzi0Ufm16NtXSUaCXXqaof
5i0yy+V8o8VN2MRvbvoq92t95ZIJWl2vCNKFSMxuKhEk4mTFdqOEv0LZSpIlCxXk7Gz4C1pK+uEZ
KmKvDE0VF+Qblw8fCia7Jz/uaQPCcgF9t8KCwN1OFbLO4dApKvECk0aXN9sguA2Ly3uvhM1v3iDp
/exk5wJ7Yd1Yfxwr1PM/dxGHnluZbVL8MAP+sCL2EUAhwgrdxQBNUoAsh6031bEChFDp+8aKzCWH
u2FRxCiX7XXbTQfj8EuS1xz0mnavQ+mD10ndgLtYcrRmNjxgSxDgJDRI49YUwj+aCAIk329lD7dZ
3QHyin8zutajLbLextL1i4L+pcGwsRILek8A5h9w0ThRZxZtPnmlFer8wI3aPM1/heH8mzKSsiqk
QamzBV68MyunqAgD8168NO6A4wGnecWJIPTIVmuGn2sJ0M2kHSz10KpQXYG/7CUXb/wiZ80Ig6RV
b1Jegae0zs/AHgM7uXreh5CEarrGic2hb/R/FIQI87Q/Qd+aLCrPewSDlrxCU5K2pri2gyZTjOMK
KdV9QuR8dt+u3p8yhAAlaVuE5yHHhcL9yHJ+ApfSsJss0lUGNDlAU0g7/l/yJNOH9VoA1EvYXUCP
Jihb4cuw1y4+lyvAG5PlEuwJ7fMbjVFS/gFBLFpim1HjDNUVWg0iyOBzd+2RTl3bpYKazTH+94/5
56DUXnfovmP9F/jmWlRK8Cc7LQ0nQJWNqFnd20VxCbaHplSD7jidvsIeIQvWe8IdAttteLVcxvYT
a6Kx6ZNhWLAkDWwSM6NdZEXgXX0mRha0BmunbwiQEHyyrmBzbOC5F+Fh++RvIG22KIRNMjObwVqG
d0fbdQlmD1ge3dUyaSEm9QG0kRLs7foswwyiGdlpeITnYazV25ItTyLGgEwnVKTUI6BkyfrHFWfa
VkT3T8+O7B3Jet+sGSQJlFcUS/xyGEWs+RaBaVDfpOp3BkNNp3yOwZOe2sMTeGUec5RxTfct7ZSd
MS6TR0HIYf2DvUO624TOhwfgufqs4yvVJcx/itwKV0/M8FYkXLG4bqTbWA/askMWHlNnmUaCh1xu
ZUzkGDVb1UR/DnRZEtQOMixge41eCkHHMs7FAg3QJfM5krlpEj9WXtTwKKbLe77t5tgI2Jboirmh
pWHR/AutVodDzKODZ6zw0Lzn8aIMvd95b6skdD+7ZRGDEQJOuZuypotLtZVh2OjP64fsXWN5uTgp
NIuNqaO119QEMtH85vdCkAERkM590bRYZr0jYq6PN/lXi0KmK78YPA/p7bfeNmiz/dEWNX3KKDX2
yr8VbcelHJ89jYXjOLB30Ewq5hfzWf+TprH1+rUllsDWeQ9rAAKznlhf6LZaM+X4DYXXZ/WiRAaY
mwp0gtpdct2Oo7xsX4EsTp9eukhLTVzdG6HuDTj1BBBZdqCM+hsiCYtTCH/qchzX/ZKG2K+6gASr
HNX1H5C8rVy4cidT4c2AAeVwp1bWvAUU/WzRks9fM8CKdXTORaNFgx2rE8WzCZTFi9nAlZowMqvH
/xfKnC44mbhC/cBK9SYUQOVbzmHutgWB3/Fg1gZWc0bHR1KahfBEdqFWvr46wnCZirRHGPC3J3rd
XUGD+rz2IUly7AcCrEW+iS5hs8vCBbzBmz2dpc/TL7djOjYoZFGWhqSUfkDKT4lRLBkwrer3qN79
IMSgPGf22ZXWJfEfAJcH+OXo2lxGONvg2gb+UhwAdrTYJ/wacu1BQRzSKGTRkhwpzvIRLoQx2Zmy
1TFcYSJ4t1E1AstNCwzxQMh8i7382BBu3q5WFxCkguDQX/GhtmZbxabBGwZW0luXDyC4GKUxxPLX
vIqcPedLfff9UdAeOSmTNWavBn0GVmIZ7wNGDBkZajr+Kjuard6iyv8V35JQdqgpVSbVmN1xy2Si
Wik3KtoCxxNqtKEJ2vWLxUUYlhOaz9gA0AEEtkMRxlYGoPvk8b5V1VN+osZZ33Xzns7m6D2cp+bV
7qOEoMmhwx9wTk3Y/68GN+3J5ol5I+nDcW6Hdzhxqce/pgKwxXRuwgF78nJoQVQx4UN8vDmzIIwE
6N728ID2silKJsgHaIw6l0EQc8JGMYJSuEQFT0MUqjjLAVjH1cuLEZ1RbJ9vyC/AJ2rG9/mSefcO
TCMCtOIQiFS2YJC4MDgWSd8iNBNB91oYxjSdYA+2bd6rUslKcmtSgBhSOjhCxXsymba6sg6fmSFw
y9/ZbzIeBOYitF/HqVLdyer02fpHafY29W1pz+G2ueAN7hlN2pEc+I/aNZX3lMs0QFuzlj4fGBnD
yU1ozm0JzKjc0qO4OPKMnlOTlrJByYPi6XdRrHl4KRa4YLJpe/hwrbVsrQKa68Bz2KMlIAnf+Ixh
hDwtk6MejH8yUSGTWf/5Qg7bLNe4Tvswmd9CFdl665nFNRvcbxSfeEaXS4HMpqjpxvK9QPsn3cls
poCTd0UhJ+BwBnUX6KB1YcjiRLvAW/V1XVF8L5+1H6u/pxscCbXdiK9orj8sf02JD5HHhaHiE0n/
wYjfOMF6uMdc0I10SqyD1UrDpZJ3+OvBhKHfaJ2t3lB9BhbAE1CmDJWxna3R+7Croy8xWk88faCX
ogoLq2LCEqVmpjEOj8XxuLBAuReVRygYXbhLJ/FuFwABbH9aUFvmkYx5jVQ4US48kcRf3kEc4UZ9
8yWfRANKPqfh8l+xegLrr2ldwqv4Yp+Erfi2xw2ogI2BBnMa/iiNFV5Dx22dcrr09JsLckYGf+cK
ir4IZcmtMdM0wNVP5kAmkJheTvIQ5ewI2wGrmmU6ZtxKihPu95JCB21njPqLEmaJwfFiN7MnfG2H
PvneuYTgQeh7yjEzUL8BFTWB7JduZBTpplyftwqTyENrpp43OXeClBdAlazMFdAOD7/HjOdie98F
aajbKv8/MgxT72jHIfyvcByfjYhWt8m9to1zBWb85gviUQtaP91OzJ6uZwonKN2wjclUKFB1Yb5Z
IvjJfFTEUUgRloSMJtbeLMpoYqV3xtBSLhCYjKTWqPEdrw56VOLdrVQ+5BKiSe4bmIBRi34I2Fku
3lorWUCjI5dWM3Z+007oxzHH2NO9uwYdcIwFwW+5IVVGlUjZlOAQSw7/vqXZMdyPSHJx2zL31GeU
ujFuNZXPidxUa2L+N3oCKHAgjeu8twjCs2e3Je259FQ6z0Wn8Xn/71IbUAKxXRUGVhyUz5ggFJXZ
OY7zGqE6PC1EJiHWx9uNpgIsSOYg3So3ffL5A2lj4PChAiwh0wjtxv1ZH6NI7bcB3UWECZ9dfyPy
koRKHOhG7fOGr2ZHJLYoPpPkhGamUbuqXjCv/WO96l0QnEajx/Rd22/5LH9g8ehTOkDgSs9LUbJr
BlKqtqXmRGKZycD6qE20y4UX4CRnYzIemYUvB2j8viD1x+9t60YETobSUkGGSZsNWEjWFOTDaLVE
7N6Fjj+X6NIUh28YoGtJPk3LUW5xTspt1ajGwGp4/2MhrIlD3Ud48tWxGYkoUbU2KPsjzx84gVSH
pDfvcCZMCajAiEJ91IlnjLMn5aF3vo1jpuIDEkUXdPvr3ybBlagsJQS71QC/oN0+yZVgOtP7+lNK
clLJV8rNS1yz5vzUXCXFHU5YmbAoH8BplXeLXqGfGXniOiuKiptqjVGqUy5U11wlaDiUB9b1r4dr
fkUUMk3THR5hvTebHfBBFg8EkNxR7RqQ7sCoh4N/gsHbq2dqqFyAPYCUQmthcWbNR8zkwuTg8mpE
avng28XLc2dMWoAGnTx7ICH9l+r4TCIyo7tOvZfzGQnurmAUPuieaHkPUad43h748lW+QdiUTq4m
aVEen7Z7oFzCuyAcd2NIvpGf7plSJnl8IryDLhPUv2keIK5D8z7F1rBn6Qm47JsN+KsVA85H1a5P
DqCaZDFddbpMy7fPbTcnv1eG0zzAZ+w4MCu9uK9SqCQAMKUguqhPUQr7J+uaPkyYB0xtOnbiLcBG
WwredjJzedUnnFl6gbhD9/bAn/oluY++v+tSazx+rU9ZLYv+7rxJyEV++oVFKq6+7XxyoKaOh+yc
UXHaoH2fptkwvMA0uPXd1iPHSlMPsMDgCJRFtcS8FFwH1m3p4SGDdI0ivXqCrMdQm4PT9v9h58wc
YSqhWohyqZBMyUHCtsaIcchs++saNP25XJHM/sVzdPSFKZ1jMuHD+8JfNbjaupO8xIbsDl10PUTk
hWU1Iw2jEL92+HQlRI7/ZAFMGwKCRrc1Lx97SkA43VZ/vzkwF/wLKQn8SOygXRTVVdsVmzUt2+u1
d4lamGlvgK+tQoqPRdDZ4S+yTTQbnC0SPRvm935jv9zas4+L5sSUcNupG4Uc6Tr3fNIpBSEOib9K
yOdFpSigADkJSyOkYjCPCC+b6qcb8IrU5/4jLOrnYwGtaDO+Ph8P1ucXqjWjIBapDW5qOIVfq41H
CkvLcKnVM3Ypx6a5Cs50u91S6cQBB3razJm7wAyqG6z7Co1SmQkZQ7UBLUkNWnuRegF3+cDifJKD
2PBAtds2tFkJyGQ0FGER78jgwH4MRIf7QIGzsDl5erhf/yIY8AYJ7fTu2i0sEN659Ti5dxakacg0
uteAnS1ULdj7g/PmEIhrBf6ko+CTMeszyTCFce5LRu6rP9SXti1R46nXWO1Xh2clVwKqiaXUPSDA
v4xSzKBSBMaIrTWUtqXh3n34p19nWEfsL/gTPsEFu9vBdOFCR2JF9uzrhfdi2HmIRyhHpaBDhHth
lRC26ihqL6XnTW8mn6Qx/z/j6LudjQ+9HFXWzx/nGNhjquPpyrpYH9QPz6B5l9eAvhxcck1iX8qO
S4Qgn3B4/T6Dg4w+x/7YZWGT8PGOXUnUbk/DXYo8zp+TpkyFIuEZs0fJOAzRnFelh8JnXaUr42CS
Eyz5/okgjJEgouZLHVe4vzWEgxtx3losng2gYeTHp8jTHMj5sZqyWePv52vv806g/uk9r/mlKgTd
LoOOOIMyT+CP4YJ9XsVTJYjwNJlj5vuQ+fv4aX6LKrNwem9f3kHCQXZuWB6HreTuh+PBG9hlVSJH
zYHVZN7Vmm2OB0n+dc/0rVNXCpxz1/iwRdcirmiaDDBiKNtylmcA2yTUjHOI2eVr1iDWl9Yl3nmY
ffmna20Zc8/gpAbntJvlMSYa1quD5U6zuCycHuAVBaSTQudcewE8IWuEYpvIlY+Ndhzoxnqoj4/C
gjmlRTPd9jvujEk+pJLvN2q+7nb8SLR5pUr0itsowS/mW1ZxnySI9hR4TBHZondBE4/Hvm7JCBXz
SG8MwQR0eWE8hFdyYmjLOlUCZOJjwmbWh0SZigmk4uepeoRv9E4ab4aiDmMB36BwFQS1MDf4D4Ql
tMLnZL/dMjf2xDLMFJeb8D4Q943zjRfkH4++VeXYYWGQFfNTtkDT1F3/BMrWPaLaNXrhjc5u6uR/
JCwAG84M5fP/KCIX3Iz+/jkgm3hqikQOIy6jwVx8tELS5ORK3Xd/+/jA5CDZSE3JO5sZvV4NPtuV
xGvrFVWrGlx4WU+lQLKfhgKhwGK3ouU639lxtX/fSPbMFQS6OGN4IWtAvgrP7DLrpMrvgnbtMMp8
wvhl0QT/4AXY52I9hW2rONneF7Sq9ydyJ+SxJ8P2t9hrel2v+gFPJRLzgufXd41s2STeYHYLS+Bw
z1l+nSkmRCdgkNtACQ2NTnXeei/doI0ag+x4C+m+a0GlflL4hiz0zG5R+OwFcu0nWKiNKxobXb5m
ZMGjpfSBVyDjPuPz3Zmz7UEHq8R4KtSmvd5OLj/guIEuh2xi47Dysp1lAg0BUlGpEKwKGj+7UyoR
fiYbZ/uFBl8U556N/1Ult9o/Pa6UmhyoEksTxT7ynlM6wYdEbU9PJnhdr2PgrLispv0UB8t3co+U
U1HZcXgRkD+o8YxQrTbLU/Tnh1hxK5UhLTwYnb0gikVhDpU+vTY8+V7oPHXh9JT3jG3IeuryKZPg
e7+PTqPsuda/MGc4rYh9miDPhRSh+CK95GD3P/1aU69fCXLWHkx8uWVhqq78vZEn1ehtVcgxFPiv
/HgpLdV4ttbtydD/nO1SvuKpNNgrjC8pLbJOejgKKC5oRgXTLPbGluZitexQPEJEJAIgsk/z5SNX
Bbz9fYcHBrTr3rAY+MbNjBlGIwXfCrnadtMfMFxQJLzFW3ouqPcflqi6ud2k2B7z1nQpJ0iP/1gh
yjCMk0gUymo/HffCt3nUYo4QQbczksVeonrlq0+LRx291SHUXCgjqEQibng4qZF0BtbjE3lkp0gA
lEtjOsQHlnxhLGKo6m/tNQ4g0WGceGvr3+jyFj3p6gGVU0r/BdDPjvTavIGscRzI49eG+wHHkmwB
oH0EAwfEPTtqo2gC5yMW7NxvcAedaUlHNKgbUBh0YN/bQizJuWxbLaeCHuY5VvDNNlpgM9bMIK2y
M799KwuwqNrfo61CLcCbptmwbBbTbRXIO/4fiVu1pgVoFyDPHt/TSOiNWFTjlCIv6bL2WQsNqYAF
oHFTyG7su2xva7IQAxz8/g3QwNpQ1KcdQJRs7+5tKsRjqOxzhQHbH/zZpWU2GOnm0LWUhnkcR0Wk
CNcDFeIlJYHLRpy6/KZcsxZcxQVGO6EdXNITWp69sziizDdxWafJul0BJhs3O0r+0/aws0YPNGF9
i9XMEZzGt63GbT3cr8BFyckWRBw2jxlE6Z8NJiW2iTJE8DPyOzy6xo+UPn4QLgD5Hzu5Z86MVUhM
MzVLEzr2OiUVd+fp9hqNeox/VL/I//YhmumZpVo4FH1Pl6jwTX+AsaKzAdfqNKW6ENXCaR3nfkTs
ge2hxTAHg9TPUnURfHv/7//PhNzuMhbuvPfIwseWCyjSp9pglGsOAhtFwQQF0ULb3BaoUjXEwtmQ
o5JmyGVIdbQP6LUjrnLqi4hVkhh6pbC796mZAeC5v2OEM8rSY2nkwH1Ef+yyl2UnojGsxWnG095p
vyafdBNFFrPmT9Q8waqU6myvEE9UCZ4jrFomZJ5sCk9DupEAljacPO+2ktd3l3yyqLZzF1+T1Z44
fjtO64fgKkHYfawazs9ajmviCsXdIFIDBaRvCp0NIEm1yQTrIlUlmZ4axuSZpJzho4DQE8zZf53W
zhiW2qqZalTa2mx6cLDkRAGHdoxqGyR8pvOQxoj/UYV2r4Zmh13O1nC93tKANeKrwfQ2y8xerFOp
L2/Anj5sFQfwsTSfkLJKEX1d6RkLPgx7uTm5rWPWJ6MgZOsYw/xRqohbB2XuQKkgYGtDU04jxzfV
nSP5WGjuGE3L0giG/bm1xU4PuUcfYF2KXMWE4MrOhAnheQBwGSxKC8jelUjZYvwLZmWihRXqFShB
CHnbezkG0VB2Vz1L7s6Tk12HQEeukQ8CmcVc5+c/pC9Nh3xMTEdELq3f9Cw3Tr4i5KUMnwnxj0t4
jAhlSFADStltXd6aD1iP71/eihooQ4pNo13yV4v4yRkhmEUcGt3jMrB0dP0JNZOSXSQRYZ4Dv3Qa
Hdq52AdeG27JDmzSwPnfcB27yXmBmmx6KNAnVVNDi4UFer+A3OVRSfklTdQ7CkK6E4UcFy93NGVJ
JXryWUMYzKxg8fqe4GxAaPKWvEe8m94lgdrQ5ebwhw2jz5HtgYnvsrlF5aqnwQid2F/0AEDcJEoJ
RJZbTZcNeBX21Oa/ibJYpLnq47TS2wqQVKg/WgSmCKbi3CIIAkdTHN0GV8mp/epUr4tckPmrl5Lg
yTh2MzdRQw+CN5SNheiCyVE4SL/bHShykwWe54WzAGvG60Vj7OvqeOBdjfi5qXi9p09dg4N+liLM
3Hro87r8wYdjCucZgEJdRLAuu8HvXyPNe/g0cPyHAdHcY1GswEwsTwXkAy6lne4zzarBT+zpBydq
KKfTG4VqWZDM45//Yn4Oddn55/qk9WIQf7EiUtST4tES7knOIRWxGxEfVFxkw3qrBL7OUo0tZiie
JN6thvk4nOarhYSB1tfQXGwBSOGdzMZeT9NsV6sicsK9SzMIgITIs77/Vl5Fk15VMgrNG+z+nwbW
uO5Hv60Rgwj5vTonfHs8m6RgplT5nnK9AjkyaS0N77HLQ+SHaufJUx+uK/PyxaQgu4DdivaVJq6i
1QihRYhZr2oL+7xr/V0CwEuub6nhb4eJGaNnsvZcL9HRNTCV4HEJhWbVlDWlEePhFwzysQ8MyMd8
0h6rDAlpKcY+TF76drwtPd3zBGy6GnuhHv9+3xXKCyxZxuQs/SH8ZIihqt8GAYPYCpIUG0yMFmFl
RMJxhQYqmSsrL19rS7jBTrpJXh+pbmAtGs7w+k1hRpo2r1qVG/UD+khG2EYmZgiy83QlC/51aH2u
QfSknaOHxaQbw1tq7BNDMRJnR8KtjJ8eu70YbQHXciT5CqP9pgt5eXB06NXNtyu4GIRCMSroksxO
YPfrb5y6p77uy083kNFqkdpsMH0ZwrSEQmUEZ46VlNXf2MkRP5fHTyi3Q8F0Nxb/feVJJq3XgSBZ
hDp5DjK81O3ifPhFYrYjic1cITVqHzqFMsLCnGI94JmXGqd8vBRHoPyNiXok/TkRfNpxXIcGPf6V
edfwigyPU+wP6fZpulc506MD3R5lqzVBQBh4h8PqJv/rWdAuzWZGMfwH+fHxFr00+sdfeU2St5Yk
gWLDw5jiSvtewJl5qqB47/YvbWPVfkW04dvtV5dgr5/9Sl1VEK8ezgi67FvSgFj8Zs13SfeDmaQC
jg8O2KsUGiPXKTZJfCfj+ffapgj0KPpAPNBS5zr7d321WQKkUPLf99qghPNMrQQDTdsDhoihAr7s
7rY354cWQ18vTnvngfOEmoyCRT2UiljWTKYUh7MFqfVmyUdS1doAXODYNDtRnA87fi8tVWqc7OTK
9dNVKZPfnjAxi4x9Jf5yjhYi/zTGdTMumUfgCTgOfpuZ4RpfueASEH2WhNAMdDbx1zjNUuKPMluC
4iv52eiiezEIxrXu4fedeH7p0E4U0DMGMFurRrIi8HroD9IBJip8zPWcXh/IUb2f/9Ggi++GntPv
/nb2CJal+m+qrD7clm7h29oOx2VOSsBl96yGTLkIXQ7ZO9PCvmfxsi75ek5npUo4R67D70tMrxjY
WupMA+c2swfYDeaQK6cPZmHOoa/7GAc+vHrRYo3vCcjdYLfiuet686h4KIPVwJUXAcMVkIwGhhqo
n82Gg4uTTC1IC7NOx3QDFFFULJuGXkP6PC1QtOySQKId0hohSrjcfUjAnpTv6zHGS1AgRx87oXT3
L2fkOvJlGc2PjqrrLwzzoYoEaF5oYvz5jzONKtgPzM+PlA+PrXeu6UNKhdqk4rqWvxCA/1APxUWx
LfNRpV8+H7NOmLXT10paqO3208I+XN90f9byALATuA/FEIXQk1rGtLVYC2WP+YIBufPDd/pybfHk
lGOyTU2Yk6SMgRI5a19OkC3uUrQs79E/VYIqhFJUyCPSXQHMNIBa6vd4TNteu/JUnRQTbN34o+HP
8EXeqJUEpVSs5gmzgi3XOMGjRlzNCzHl+KPkwQWHjIy9SXgdbhXEgc8irTp72pkoj2LUMGE+l27R
MBaVrehQ7wZbSu/56N0ymr94E+ldlLWPnvsjFKZYkimSIpfFixt5ZWEdFOYONRXX9XtsaWsdUNDQ
kTwhAULQmf4E5BxXXxevKpfPkoBSgQ8kyKyqPhYN9Cwd2Q6QLRkaSyJVsmJA/bpXlFCKpNNlXYiu
F7O/em5XoV3St8nIIozwhMxXzo6+jrEFg/CH/GDZNfjnVxo4Ue9HRhf8FFaWgDe0PBvM1hbCeAmD
S5Z+pahSOvPOK3RJDAQQfW+IBrGI3l6Du4N5BEGPBm8EzOwqG820edv8sellNjs4KjopdOJ+qzwx
jxupPwsJuYtfzKpkoz2YIGsuiG5EzfZ/N4lY3ybWaEr/nNZUa7bK7bcrtwxO5mWMZQ4Wh0U1rwmH
MCE7diQK77KcPoBiiijAIh7xldNA3dVi2FOYPNEifum8H+hZXJMtp0IAfUFTwLKQeTmb87R/Zpoj
kk/R7SzUfbYMQzbHdwWj9Jb41XuvqxZTynwmK9PqiUdsIoveuqXDv+CajAFiFaP8hvQT3Lma79tk
Kd9Qf/ct5MMnsmkH1LoBxj4iGX1w2O8bt9kMizCoytWOJLJVcRcATFTk0QlGoyvbevlMoFRytkCx
tdVJqTgrK7zBTJRyfy/LSugAKKhTLYLhGHAFvEViPBiP1lTcNSVtutguKWbSrfBvAGF2vVQWExJG
983i3YHxsy3htuLN9nIYz35eszkagLlfKOMsvXdD90XvGyw8h3s23OL3EHvu6SmX3ycUwb/QWK6h
blA1kOKGfWkOsS6Y8buB/qtY4yt+83/ENymLhIryIleRNDdhJz4gWEgzgZYAxmeFcbsv84gnegLT
EGudKWDqmDeBJxXGZmZZdhY9gNtY80am5AqDbmaBoMLXFa4U411Ccn78XGJ51R7W/5IRBtTcop3z
JrgVfvopoaWEI5OoJChmBQZ0ETtUV02fF/d+ugRbeoN1tM/DXkk3EMVsr6LD4EePUVXJRPVLgCmu
WkM/LFFF9ITqf67hbD4eX0+S/NFuijFxyQcTf8rO3QrZWHw8RKdkbf3OfLaHSspp7gY1+K6mTbNI
shHZn7ZSR7CiQGrNdcFMmZGZTOH/pw9E6zELKyzoq79eWdGxR90tSlGO0p+EfIul200gdrqwB/Fc
MSQd2iRgYhws6EinseYMAAL/ECBF/D9zydRipWKsDXc54SvPEAYZ1ko+Tq0f/bCVKd0eYOnQxiiv
S43pfCGapGNA30DMfR+O/OtdqhlrPxZYh1vX8Xm2AKLQ8keFUtzXr3YB0CRU2tNH4T+ZSDgeiiHc
GAJjZsmXGP/DiA6+7oGxQqZmzyPERXMmYDSBzm+mz/ZMtpxRtrSZuIBnFycsCou3hgz14uAIJocL
kHr2B1UCiFmRzh2cWh6L0jnc/OSkeHZBPVdwd3SHfnwuFtynb6iJI6Q3TcvKzA27aXn/0uOOrwzg
+DwfBReV+zGjOdZMzbRGq/9aAn1udXa2hhzD/J4znp9e8U3a8lDo+ARxh2dB0yBRgcOijT0hq923
EJu7CQcbIlu2x6bpBpJh1qkd78Z4L2chsJ6HZMtIJEVqsxgwH94LWsbbDaEPPtKi5VsQ6syrut7B
PL4YwOtoJRIrJ4NRUieOLPN2rSy9HA45xLkZrqbKJ15EEa3NHHgYRIbhjXgFylxf3qszVTQBKwpg
J8UNWuBLiwUUvTmbcqAabIlms1F02NqL5bfrUeCy121dbX6ECUamtWrAlChaJ77s1IFI7hBB8R7t
6iOOvQgFsIB0XJ4mIYO+9NyMT43s6NkkjN7lD/tzRd3Z2qLFQmpvewJPfzC6RPaWxV0OZE0loGZ0
10o04ElvOe41ntE9WBtH5CeLh1AWek6ZWKjdrRCuLk+kwEMCl4Djl1ylKnJlLl3YntUYC+g7MTL0
Aq4oRIoQ9DNMBi1yN8TPsj5YTnlGqq1aSokFsX6bDkekF7/htqjf3YJI2kMLafTdQVuHAnVp53xY
/jD31YyFKuTxe02kFsYoHgR3EQ0S22y8anu/QS/PJlSigyrMWfrxvN9OXxggmPOx5hRgkGmUpaEA
C8YruEuAKiz14jt09jzU8vNF+HOqSYcddvUrSaD/nqoA7OUhLN9yBZSTTcj3jACg+COXkqhf+SGg
BdpG1yogmXY7HW7Hamxxm/Z2+FxvpfEWJyh2m3d3ZReCuwn4nVJyGIeeRoV/8fI25Ea5mEwigtjK
4SZ9Hy/Ehc8FuIHwyqWMP851L/mP/JD/0gegS34wSuEtIB8ZWxu9XtrPWkI+EHeDWk5WL41agJBj
cXR5HRg8tUuvAJsYvd3g4l2nbhM4LRcU0sjo2rH0S+iAPuzZ1CdKomwZUrdsKRz5W5lbWz07uWDa
4j6l/rVPfnuqdyyJtewLs+a6gIYOTAbO/TUjtKMwp9YOxECO4bVppD/JBn3Mk8vnVq728ve3MVm8
iVhYxI8jKrewa+TWlS8icX87BY2mvdr2TZR8PV+ncLU6JD2o4kdXK4juyi+POGnMaNkGZQkB59QR
mjgleHnuoticK0cFLJpjnfDSDSVM3qtIa4ReePWpYDIc7poqHxRm/ZnyIk2/Z9V4Ys4ICQSoDKuu
8xrEzc22GKHtFaAptZ+hckVElkIVOmzIQW0VZon6FECRdR0juSRi0xWEiLodzS6EJ3JI02h27dj8
l8+csjPjw3WanzhudmrCuHPmCG7tKTDEjPXA7p9hYgH5naa0xyvJvuAUqT9qg0aAvGay8VSmms+B
tq/GSJhmeBGa3F6MIWNMdbIgtg3MVVvROE0SMKkKbtJTq2TGqGrzdvJMuyZ719lGFpRUnNm4j+lO
p8l7eiiLkyFEN9gjSPyN4T8/HGP/nwg0xHH4nnwebc9SyEsCUPE3igJ34ezMS5Uz3LvxhpmedOiN
JDRREE6BeethES0tBrUHXfzKAhdMtZ7ORm18UNIdlULLi2DTzwNCPKlOgP/n1qR7BewAIN2+bMv3
nPZcdshQUO7ArJsZ/7O5IwbqZcxkMPR1tujHbDJNla58SMexO2+4n5BoeAAy0qy6Cb0GfvSqA+OT
XAv77G5ZloXpt/JcNw3F89JpU+FihOZ3YlYsVEuyrWsifSLpL1fMt1L1vhhgQcauKZyPx/xkrX1l
sFjWRoJNZHhZhbnmFEallwGExToy0pmDIcfT8hpcybspZO9x1/rkuBbQchTWjmAjNWvXmKCl2Lax
whvIaojHsQPeuDuRkdqBbDYs5/wn+8Yea73TRFFoG/dQ2ilXVlRO8rQI6ARVjHpGBm1SCFSkwc+O
payXMnMRk7PnJUeubLcTYyRTHGZVsa6k1c53T+f4MQtJwldtapG7x5EQISTba5Gl3PL8fow4cKZm
33lXqYcUU2rdJAAkmm4k9zF9DnB3BTW7oifIVkvSsGND0iWxfqC3szRmvu9RBkhVx3bj3TaGzPyB
jRpKHMfJt+bAigGTOpJsrcmmt4mIIyb8AfjP+B/jZyt8ovKD9TVRiHMSBB57YR2s4/AITp2ehNYl
bqAR4zIud1Vca5yYq+OtxCwg1f8jciF1ziCGkoumcCOvV7Gb8028gsiXUBkm1i5KHmjR5PTs2GiE
nAmpWRMh5DhHITOh7qqC6QbwczVynZtFHheU3vyx6F/w53/GVkYG2RvXwBp1ueMbslGd2/b9ksmJ
+mGIfe+lJ0oZIChf94EImXrtZRpjH8lksG0OQ2EcCr3v42rqKs9BYa5QZp6nDYHFiNifVndr1OlL
tW/Qm8o80Sb/ofDsJcUclneI2YgbnzppjNxNG0N83VdaDT3aqTfbdnlxFhrB/nN5vYCp4O0XX7f0
f8K3n9G4lQD+HcU2O3sqw7+8WWLe6KHcxV+UtqumhUAez27GEbZ6ZvlMbXTUry9Hl4nuyhO7J9kC
o+gr2XztHw9w0LpKFcd3M68g8bpjPJvKRfmuWryc282PHsT0I03dhRE0VYLUb+uX8ELi+dVFlBkl
zLj316JZBPHhNBQT7kiS+wa4sH9iaXzpYhiR/OfKkPs1eVT4Dkg9nSkx2QK4lMJHW8MoqBAJKCK/
YHROfs3JJROgemmHunDrMsPXltyWLISYebuUfFC/vI16V1VPZgEvKDaU0z4tE4CiGyhk7PKzFlbo
jWUFNC5tLE2H+0Gw0t8LTljrgf5UntVU4vrYwUIe5ck8d+mwmDcrM85NLj1Wzk2ZVGnKL4Cv9pKP
9K0pVf+9inrLiVBrygORqADrgYqKgFmhNVjU4w19x6/V+z4F9CjiL6hAG/puN6t5x1FRwsvlXmHq
8d3T2bdkcxcDMN2cekmEwIpzXi1TgF4I32aLXdrbyUuFoPJe04D48DzrLaIs0YO2FiywZuWEs9ej
IHBi5+t+bpdz5TpQTaTY4UtSLVbRZomSJoaBZ0rW4c3EVbitvPoiUwqZA2tRwxXZJe8pmSP0+PRe
4vhqlKR9y/tMmXfAp41y2Ss/ewBDTrM721yJzq7DxHXPh/p5N7qJloTgyV/54ENriwl5UAUAutNH
Bc6k6yOCVQrvE+L8h+1zSOeRRmQmWJiuWRJslPeSTILJu1BJ0hdUQUmkbWTsH3mTK3xAHJTFu7LV
/ohVQc5q20m8lDxlM+jTNKWuum5TLW497fCAOUJLVZ3EmGhwsRvzUbIxbMo/X4x1zYrYya49kLNR
iyRFMq8vKwLYghZqsuv5FmCi2LS0XLhaNQ92PmKbq4a0iEeo5wLTwdOuQmB/X0q/+QkIWDBd3dZx
/AE6y1paZ3RrEZAgsUo0Ep3bF33/VMT2E9nEIwMVDIS673ojE3HvU4wTvtLH7n/hf/gGnFxM3I4e
Zr+5tjIZy/0XPDCEx67EP79kibbyEsZxFf762DdLjqOaFQ7G5qO1iObP8rub3a9fdKKvW5LZHSqq
zWaRUzl85julhIKV6OIMiAAq2zY/0XH7AVcX/H5A+6fhGufP1zRYJsOzucMdwqqmpAnAahi0B87T
gR4K3NA5gmg7jxRZneqdJwX+rU+RODFj6BmIz9NsfO/FCSnnbZmfXEVwT2LF+CCauFapZaWeoj9E
Mxm2HxYkYEUlibuyP42J9RUaP69EFjnQd6LFxtDwECb9AhJA2o+eq51RflJEPfyp799cHuyGaJ2a
/tos6+XqvOJpk/XGEilR7jnu2eZnnqw+a2hVS6567GqbcfQ9iUTkpQbBQdEsJ8rz2B8zM5/vWwzA
iLmnVL7gbi919jSBMZN7+aOHLPsblg3fSbhpu46mUdSQ2LhiffzA8Pymhuwgi3VKgX1q4dIm1kH2
HHtV7CzTx8AnMd+Hnjzycg6IR1oO4FdSspD/UdBU9XlotNs5Q52C3mG9YfwQtChUDhAbKp63KWQ5
ohCeqecED4AhMhiR9rWI5RhsbxsT5H/OU0jk+6agjkABOB6DG5F0Z+p6vrQjQjd/XWRLkB3ay7wy
PSpegq8C+jYJtvYy3piKvkL3kqNVR1/TY8aQZcafHysgWIGx+GD3uLcCgwksO2yYUDtdN4O5Dlre
LyPtL7YDulaU9qmXn9NLeOZagWRFqpin/evncfv4Z0dlFvCkDURQwXEJFSUp3xhoVgEcxT15nkds
/s70jJmR8Pg2ZO2Zw2GL65UZaUH7htbvgWYHECBxV4Y3TpqBVkMHfu48itlFUtw08DWpRvHCzK0E
A1D4VR5ypP2REKc5A57AI3aPY2bM+Mur2LNfAkCLo5S2SaU71wmLIRNqhE5GJYMUituzMSl/ewrD
kECLYE6KOpX3TCYJBnnnmBcfHOZ5yOXNlYeUApwN9Tq6cDSk/E/+0wEa6RhoSSWv7UKbcc6bcj9b
FfJtwvW7Ish/28d4SLTKPo0R2QRAhs5505zmGB4KOMyg6EraAFYXGVUMFCbTVCLs3G6n+lgL60Sb
7WLPuODyvETFaOgSoSDczJIExHdyn7+R3ry+MUcRgHKxhq8kPSC4OjlSPBmDtcEDaQZo0PdPbK//
NvlUzZDvOF4R+61DBi7zdgWe4sfTOLKilajrSJXGtJSpwXT5/vjYhjzNo0hbXmm39BTcCT+PfMjM
AK8IWeRwJb29PpHO+eC/XrIILRShSDTS87HiHHQrJBgty82lzDLvAqXQfiElZa11Mrni304bXKoN
HW9yQWIiSRrPa1mPFlPqW0HJqHAsa9OqIOyFmJUtej5z/AktyEJ0lGSxz4S9nEuJK1hL/v9Q1Wvr
t8CvSRhGU608B3QzyHbyGBCYW1rt2DypZA8ZpONstRj9x1aZ/zQ3pyuMLgPe0l7J9NPAkPZcG9ZY
t3UpUKR7nrPzYDeEvrL0uQMXlOAZI0ozQb5lUoyzM44ilxnxJAlmSbyC2Mnfwaqe5PybphP3jP7p
zFobkDRlHhRwpXPKJrJXhrqsVWFlxFMa++6B5SF7qW3qNkS6MqZfLMJ/zi5xbLJURTL/3Ir6xm/a
0YHbJPk092A8TnkdftZm7kuk+okAeW/+78NAj0IaJNrKipexYptWNhNhvi2196AwJ7WRTJlVmb0z
zbQWsJPKFbE1sItt7xyp4WSAfHtJh8JCffjSBBzzqPI6ZXc2UqPwA8zWV4h5NCzDm6m/0zFT86fP
VskGja7bPIgtpiC8Su3ApWIQTAsV1bFi2FYCU7QDD0darkWF9MQGp3k/cHoWT/R38/WXbQpolLsq
B20x6R5oX4HMudKOOkV0280maJL03Ulvk3PCAgWKxafKOOwVBrMUZ+oJZf8FSsIstwCuM7NHdrKH
MRSmecdo4e6+hZO5LYrUKIgxLXVnYciZSicGU5sMaCXlEsw94KKmUM7FKIXJ+9603ZVaE2AQkua9
t7henQG6xDOW6hcf7O0CJZLSnPpQ/OUlr3GgfhguPDG8L5yKtouN1ShTjVgvJGs77rPGogyt7JWY
Pil47gjF93uUJvISYQscBdnny8/J07zXOTasDRBfDvMW56rtQyw3hoBmNrp4SnkGNRZnh3+hg66l
xmyjXrIKBFPUION8QuaiQbtk+aEUDrxirzsOViKf6GGg0ZN8TDJ2M/V7aQDlyj2nDLyP521MXyFi
m4EUEtykI2vULaGC9rf8I4o+LD2yn59jcp5ljwBOpm5oZGda8jFqSsBYkuCT9rgENa6FloWxwUDu
nVkGh2K6H5bz9vCDWp6VX/EowdUAK6relA1UP/FjifhkevEH2Q6zpkOa9eZsKx8lRB3bamQHrw5y
0QK41YWIhw85FxGzMbV9hxvWn7CPaQ1HDNQl16hR656uRYUmqHhv35HTg8bowE1oSGq5iLjsJe2v
BgeNS2eUoZqSWFUDlnoiXenvmAIOQ9edFG17pkuUE25zepnR5VUd90ggbs/zGd2wjHtntqzx9NZZ
iPU9MSldDY/CqeoPRy3xu4KXE+0VP7yLvTFr6d1nRRPu5b3WmQAFJmRgq9UeGW2gE4RaOJGHCNOV
Rs+jzcvoqdst92lUtOlh5xmB08TnLXuooCzUOKhYLzGZCnZy27s7QOn4Lp9CwFwXHLDQTz8rHMww
Pylr5AjY/pL2cRaWmOOAXnOeK17SX2hMxBu6XgulN8TvIWvNb1QJMMBlZJhLPzXBMKLkxc94V8gM
TrgcaIG6hvBrgrobsIiDih3CymeT+gm8xWn9FD++2fZPHKFezlg2GCq4mF+2p/DOns16xmLFLkGr
T+vpwi1ZOayauaBj830ljV2kUS4eRPToM8a/g3FfqnLxGVli3NjtXiydPlnKf6TbHVKMBrule6Tx
HzuQ9Etblh38rEjeaG64YS6EY9kCn2mkX6hK8CxDRakeWVqSYXqGx2myZEOflE9SWMeQrUpOvOKg
4CqxzTIHxkhWemwyc+2GtRo5ilw01YKa6ZxcEj35vQnRKbrI/7giosmehRg74vp2Y9V+JaHl4rYq
aSYTzIdrLBtVqXyqd+JgLTqtfpiMU9ngjpglFKvXKuWPftXQR4mSRNGbbC1uY29KqZg186vjiGD8
46m/kE5WOYqf3bA1CWqB+woOfs6FhS5uImvK82UDCeEvmGTPfJEZ5kXEIQYaAEAxmx2yEqBmtArB
Icfkb/ISdU0TrlAysFF/h4/tFYyoZbF4NEv60pYb4Up39vO/D3xnzmOQ+gw+h64l2ehH8H+ej4Rq
CnU4nYFdMRvCTTpUNuFFy7FPP/tZdR3+yQRjCiVD7yUls+hLTOGZT/O/n5BGnhfkAiSf6mWtj8P5
ZK+UruVRBpaL/HX/t4wThiASncHvEkn+mJG2Y/n6VLuMqdw5vmzA/jwxCJoWrYCzViF1KyoUQVWV
lz4Ks8twRIsVv81w9gdZXggzn8WowFM4b/QOgOcbjwSO1kL0MqSBLdCq3Saa6j/8J3XA5f1flb+p
HDa3EibH5S6tCKGEbFQvJ8+SQJEVBnbDQ0EfPof35UhlQ2mDOe2sL2qgN3D4rFeyMUBw44cXRbmU
xZfhDLWme7nAi9jP9gKhFvgkW3KSynucaGfWBm5MqweTjxjH+mqtciaPgD+zDOBjQ2foMZRBSxI1
QDR+y6t4CQsl7w0o5SRdMoyafjrYwnP8iA+iCd5wOgoaGTUUAlZU/kJ4FAww2HDzzFhy53CCmRfj
5U7g8F9Dasvd02Gq6QJ62S04Tuw01GQqL9eAQn0FevdteiBXexiYiZtC2N9akoPw39nD9u+oBG5/
tafWcO+wx9S4QpNBV66sNMB0bF27N6LSHKp3UP2C6k+wFc44nwGjNzxkXUp4TrxE3dZB1/cILNii
T6HUQ40XYinUOJYXzgdeFQs//X9pf+1iPjTc68kbezpP+4rHm/4/5t+ROeYDlKetcwP848SeusGZ
wQ0p93kWyMD9vd8SZwrr6YQDuOrknWn/f/jWxQc4HKGzviTf8IOd9mFEKKNWLRfmSjo81lx5A75N
eSrfI+JtBfdwoaxZOnGcP/UEyUOWQYNFIa2wWwZJLKmtr8/s08ww2otxBRwqTipq5C5aAFYG8uSi
BPHO4E5l9bpkL99fgUO5z+unzHHRuRk4ggSkAtLDJNxARY76DtB50iPFZ8324EyJBVrI60yTtwpG
3U+5i8rlf7GSfnHy/V1xO1eMReHafAadEgOLtylQD5Vetk1omC8jAfb8si0aHtRdBS+4DNNwx3RN
349XlpdDpK7bezRBAjkMhopyHXGRmmiQYjrr/F0xCQTLeZn8vrOMf1s4tqwKSyU4C1QEO59Q/cvN
xIoLePDMh+I2BWzV6ABpENG3eG+pVUzmeko17VT9Wz/yzlYC/bXCxkRO7RYAtIn99Y9j8uKSY0wZ
7sNCKisBomwi0fnaNj76orL8Rkv4KlmeZYbfq/kSrOD6wI0C11pLBiQLeGvcR7sXwApYi9+AHKQ9
zEfYoJB3hr30DSU5kFalmOoSG8yj5D3OtNsveVYCEIy9Inzk0ULhO7P/ZlQfO1PcBeJkNzv2N55V
AeT6bkRAsV0CeczYSAgJc9OhoDuV6qfEkpl3ASg2svji5Edi6scquTmnKpurCirw+qiHaTv8HIJp
q7Ay+FVJ9tUb0rA/SD4o5RLineee87ilPFBd/A/krND/DyfbS+tRP9NtbzR+9u6pmZ/O0wfg6ojb
ZWnlxsJSQa/ernXYjnrJ7JOBREX2yMIQkb3ZkXJlKv6o/PD8fiyU1hafZj0GoSX11MbLozhxuVl6
EoBpuXuhgm0ovk39UTtfRCc/+niLDlJboCwFSdAGN+lO4bBjoYaaJVaSrhhdYbe51SEHus5R0xaF
kcaTZr5WHyXvwb9BMuwPY7EgZzDx9TFZSYxebS+IAxILVMTqWzclvYJp2Y1UqwuBT6WdeGYDXxHW
Gx23ALp3n8XWkYlrj43vl9vHw+2IO9agTVRTuQrGMkm9EkUMOM1VpUbkkftTP5dV4S2TtCvPUBf4
QI2MIGGms9mq4Wi+sQ5VoE/4HUjXSsOjFv2AydiIJckQJkGYfHjTIeD25NZf7MPa6k3vhmGY1XO6
K/RW/8c3umyBwZVw2QB9oYiinex7bXRVbJhstRuvyyrJhgp21rqmoJMZN48hvixOS66XKpUAPSe/
1REDeMuEB5QXupO13A/w4jy0zWw9JlNSzC2XBKYw2nKqDQ9if7yKIqMDpCb9hO+44pjJcW/fASRe
l0xfGL1+WOqmHir9gdyNrVTF6IETTNl+WHZj2x64SyqKHcLtQYp2eu8kVnxy3cQR2dN8ISCUCj7o
BdtAfGFVyKkgt0yLTl/XHTNPXGCjkz0cy8vd1kXJhSwFEJplUykx0/PmQ1k2EKGIccl1EqWAwXGc
y2QD1ybAFvJpOmPHo9yDOsIN5qZeoGS3E5QSJk+Pu9d020Ryq2ttIfA20mUqD7wdF3HsFO8zn5nJ
eD9fjHno1vECMwsxuqWukNt7idBueQuTa7++r7yp/qFQPR+tg5FRH3vmr3N/5Ny9nXB3rfvLhTmX
fN1Y6h+r4YXQMcGJYhsSnqTwil4k2nQ2nkfB/TbkBKklrd3e1N3YOiOtC0wNdVDZwSyqcR5C7KxE
CgfZ+PeQ6hqqDwngoBgZgO2b9VXK8FaB9LARqsjsWUkf1yDc0UiTo/X+Ly9Ipt78g37I3JQ9eBXo
1MFmNWtxoVR6Pmz1vjJBi1CWMCJZA610Nug1L4x7vK+8cbaQST8wJ3NmGVXJ90FeIbmSk/qVCjg8
UJJ9P01oz1xA/kSG6zVVsH1uFw6vHS+NyZcqLYjJNge+bcbRpEUg/IEBsHeEYLUciFtOQZAwkVE7
3L/u5qUvFhGEPkafbVoIFZZOgFiQM8dEQUoVvIDu7eZt8Rl8XFYNDY2unmSmekuu3cPITO7noqW2
5mvJa5JHemx2akHGkxQtcoX2uBQbhXkE37hWejMUEphTy8Pgwp53cvliFtyI21rIqoi6lB/b7PGc
pxzN/JDCZxytackWpoymZ5W4K3ZbHCxL5ZzaUNjrxuwzGGMzOsWToprlgbscx4/FYPBiD+ltszXl
ZWpehsEJ8DlHwhj1d5opy0QrAT15fGgJT6Lb+W4JIxtI77riC30ip9qWGgdU1edECQ8c6YMZ9u4w
2Gs9lBCfTBTtWKm+eudXs1q5juIlUHVSeEfERdsGhw83ZDUvN6j6lz7yR+3ONrkdRAzw/m2pK2Lx
3GnR2KD5idwsHX3dvUUgXgH82j3lcEgnQuBTZyrvN/fFRus/0aCSO9IEmUn/KF8UHSqr6z5q1zIJ
ZYu2HUha3Ro4ZT24rpeYzgtwnBiglCp92uNYg2kLG0jsigWArRF5qaZgnz4wapsTa1EIgb2DatZw
9lSTFO/jxR1EbPrfNR7g5dQWLpOHYS0lr6S+TvTJHuKIXKbpnYEnGZ+D0YSYFX600BOc1nD/eDlM
KXi4MTUnLTjCh0Se6aN1htXh49lYTBgVL20pckyjBzvH6IMpuyQ/ynJN5gp0snQ7N3fCp7fBeE3X
eqScR1CiuQ1a7cF2BX216fn4oLZ95cqvT93BYOGfbiXt4GLTRrJVgfGVoGz1C6yiyZb4HSCeWpvB
p96mk1wiTh4h554GGNGUG+qmNMq5ouHyTufCf2VyPTpEeByN1DNKI7h2Xp+vDDNXIWsFdDA4uyKk
Noh3z+gFptFsyx46khROm/b/I8O/YLuGUGZVQDO405dQucy+k9uFaoWMv8s7uF60nCHZMRWdrZBm
eALA8EM66WsUpBqkIhVX7nDg99U4nGKXm2fJHeV6ZQ4UPmCLWE1tx8jb1Zh/Ei0C6LEVQ7I5a9oQ
e2YbrD+ML9D4u0MUhTZxnS29pagKeTMyFBV9drM/IcviwMBRv6vCS7bQ8iOrmmUmq5KsojSLr4BZ
ngrCPY/iNVQcKy/pO/igxpIKZRO26DAriaE8QR3/qTuXByMAY5nGIu0NaVrSBdgGCmgZeBhTiLsk
hW93ZYqUoP0MEboBeFW0A8+7K4+hih1i0v+C/F7yLP3knhIieWnDDeNazII0NYtZkkkeCxHMN2c1
7QrgYwZdXA8Q+FhOsx8XG0Co8JtMW+NoASHEP4Xd5RsGcPbuqFKjavv+XihicpwBMgGUjGbRCm87
PqOf1N+ojMvSAiWWhvCGDulBl0//yIioEbC3EvLQ/1R+HVeauG1bVQfLN31dtDx6NMiR9MhlzsjM
BDbyMuJmIw25YKsS2rnKC54mls/Q07JYOEg4nUTD+CQFREAGHO/EIokg8uUiJ8AVjvBWjH0xUO9a
SDeffQom/bRLG1WfP0qWnd/HJijfW6Rmn1AamxBQO1eyWy+pftI5UCIYMzlwAGn11AEwRHfwbhnb
rGRq4EivmCBMGXjnWM8xXEHST1Y2Z+V/HiWa+m7ptcnWVRFYsUi29K/2GwU6tpkm2//fNIpqWXiI
WLxCmpeDOHQ6BTV79fwhcHbRIO4zYoV32Qfi+NUEpMenAgQxlN8fD7MBej6+zB4xRN3+8z+YdCiw
5cXGe0ShJhIVoH0Rc26mOMUPXojiaNaOXzGFgeELktLqZyWfi9hKvTjx39IAkkBYcXbMnIpuqIUY
+hglbNMhN97bw//KdDFZCghRp9J0UjDjZ/HD16sMs+1Ia8PgX22w/Jj+NtaPFKtqjcJ4OAR0RHFN
U6bQ1uuCZ/c8pup8WSEKREvf/a1wseZjJVQ98O7o5WvNVv5aYpo/ULo38UdRflqETodd4QLmJaJJ
keCtUAm+En0cgRrUd2wxrEBmo92JenmagWFs++rrbCnBk86OCl2/JIg7h0Abf+iPChYkCbIjIx/u
WZ0HbEw66c8KRsnPWaFA/mZWuukR7sBjbhBhtnYcwAkw0B3IPhVGoSXOt18PmcXB6P/RBL3IJ0cO
8Fg6HcsFebSPdytl12FMhxfS9GPTu/zG7j8FaJLr/CCsv7hvIIf6banjBYzPFfN/uwFa9RPvFZNb
YFyqueSBbPx90XGLvU4Rdm2oksA8HxO+We/sUQ0KyllEMrhYcJV4bNK12HXM9Po3/Kujh+QQA8vn
ur6VGQVjeo01DDAr8x6zshZY0+VBI9R4dA7o8N+Gt6i99ABEc6A+sDC/yz/lkdsccs79x1lLMML5
2UK5HyqVpdfgAxuzdX5jZfixFsjo+ygLA8lBiBauS7gOxBF5ncOHBQVLcQHVtOq54hGs1obr3woN
oEaHtt7ERqZ0qgu8OspFM/aFEkZTZ5VZL+dp2PpM+ecGjsq5G6R/kPjcTV/fxJj8w4BepkmNrIFU
bXBgsIxcwevczdDgUp9nLWiXb1k2MpsHVcBy8nbx96XOl77eUpYA8hEvEzmrXTx4fRAbov9AMJT0
TCivWe16KMjtsjJH5GMHPBJQPT1VZ0Z50W4w81JWrvY2y5yUPaUKZBsCy2YjLMHvTTD6kOwJyhj1
+etraCd3zeYYq/BIsWFMiOfLwWi3DAVG215Oa8GwArLLfqAenhWel26OhZqvcpJwsRqkgNp5JaAV
+GabSJ+ssPQ7eJlk5gcnb+fwcCI3Rj24QTz74QhsRY5fO6JFz6WsKm0E2HfT+fYmvnzxqayDFPpu
VYYxgestYk+KAAds+vOG+1gQC0TffwfnII57AUQKecHPpoSkRshYj+m88S+qENCBLga7T6pby5Kc
RUJH+lU30u1tQh/YfwYFJsd51NeyTBkNF+ugc4yXsRI/JUD2HV2lAcPHrNBDCvDEwCMI1x3M5j6/
QfQcUC1xCH3haP5EXoeHY6nm70l04JSjEZkRrNTEFR1XdZgxKlIvVBdwLn7PnImuIB4iE5pdA+Tf
8ynoZGF/rVwr291FLYVgIxsIGZi16Fb+XZfb+EMKI0UC8M6VPnoC3PjBxspULsrZLK477Ncj8YvK
cZ4s7eHxdacFzf9tu9Uit0Bt8ljVtd56p0yVuf/zNqAAWeDljAej1VUMD6ZieQf8S6xoG4ll3eRG
RaC9IxLWfmeEdwyPhG329JqgaSvaBvVrQh9wEXmHc//LO9+XkmWgB6tjiOMogz/RTvYAofGnYu8C
XyyAVB9icmRgKI57wbLNc4XwyxUxt0nwbtttTCdbU/NVvF/4ct1m6VDVf4l7F3ILv2et3SGF6MHZ
kappfupGS8mxWlMQC+2two3oHJTm7G7N9sZHlmYViwUdH8YnZsM540ViIxkN4b5BfWrEpzoGKmpX
6Mps6lbTqK2if6Lkw8LPA5NgwDumGwhuicn+cUhiftJn9bZXrwYHxKuhfOMwl2MYp3/wAGf2Y4QD
fSzqkBbq5irT1ozG4FcrqTa8qCIGdL9vbGYxzY0MDbabSQS5DhRqDhzC72LJngQW43+vvhpSKMdg
8S53mU0wG5RbAZefJyebGbxmRn3rRfNPVD9CuhvVtkh7GqumTjtcCAvOQ/hLWukVx+BWbRs24j/T
d/cKrJZRHxrXGDEyOsntZnpr1vKavcvAZTaYWZidNo47UKkW4MPii2L3QisT0NfXY91kQ77sE1Cm
IiJUb3yW5wsgtcUhl3kfQCpRhE8SWyrI9xrHhTo9cbfkHEBUqm7YtzMyLXLjgcATwg/EbXjysPyI
myJUqh4kdrBUbmPWxZ3rqoGJ0uJgFfCUNvA0Zq5wB/EuZ14Fe8sUmAcOz9ww2PNLnEf6iO3/dlWm
lw5qF+buubXhr1YObO91qd609A9XLGWL0x3QKUuzkbR02gkE42ry8lh6xp7pvaslG9HSnCPhWNsr
Sg/WwNBjVnkKHzhs9SeiMXZhtJndKo7hR4ekyM3UkcrSZq1dKz5j1H21DWxqhSYWDrlvEsXALGbZ
Xq9tRS7+HTwSFviChu12EPztQbmYTzuowFXiNE3yk3LYINdnBeIcB37KjuTSYViJmPjGpD1P1SVp
P3AJfc7zYpvGq9xDYrVcdvzuOuWk0/AU4qnoTeY2DuiNSPCCGufDzjHbc0W1pnTPYs21d3Q8GB1Y
YBiXIPen8GwSxAC45qLsUEzFq+mDXd/mfPjuhqI/WmxQjDXszHxQeRorWhtcYR1m+87lebc0R5YT
J9Ecs5Svxqy8aaDhfR3T+bVkAXTuFeJho4AOb/KVFQJtQsE6x1rqlVH2l+M1tCuLojIdampPPctN
1riJHH7irNGmMjpEdyvT22Fe3vYCUm66cp/e611yCyUQPo1kZU8OSfK1Ysa7rErWV2VSwKunYXWO
ZTURgK5oLEpq5SGO6kwq6kEIH14/calVVqf5hzodznPAw/o3YTAMsqlyWzaOL0oG7WG/ZZztkN0D
xhDatZELJjfEHwGQzgPnr6L4hrchZCNPC978H5ASHxK8epKg2NAmOe9O25z9oJ/pbc5Lc7fi4NHu
IKAGa12LBIxO4mosH8lUSxRYXl1JHncheUFETOohUFD+Ltyq8omP3qj8+OYrmet95V6q2qSxUI+P
evmseJKG0+dbWZI6yKkQZRXipr0FOcx5FA+I73X9scwsvFfi1gzon5a4VKM/eDdrz7kgJYy7J4M7
RcZ8gY2KyuPRIu+9Q+yRHeay50WkBDDeLrGpzLFfOSnHFBc9J9LUz3upzeD7ptemQbWlUpPR1KhD
a1izNMZtKqGMhQekrdhy0VC+A5hmTmbKwqlFA1FvJpDp/7Wy8y90yRDVVLHiVFdbj5v1ZnzGprxg
JMcE8Ce1O4FdYnbsbb2N1SIuj2zpDWfCQsHSD6bG3lQWjfgQyIK/mlzMe4ZnYuQwLr9aja0wNqti
To6FAummgT2B0UOMMnrWPqYCXD0qA4hHOY+zMU4AiKgYgdnuFxeGpmewIeCwE4K2Rekr/nyi+Fqd
kfKq1K5guuCsS8k9W9/EDSZhCJBv39O8BXa+5KWYp3hnpUJHWVf106KMNC0iT5re20DZzzP8QXJB
W6gyYSUPOCzzyaF4T7Fg/RVoQ4DU2yLhhlw7DXexafytCGRkgCiYKpYNOUdpTxfTS/NpBTDTmgVm
88wzdATE8PM2sLEKhsx2xca7unA5nTPyEj9e8/9TXCo+cZQ4cNHBrhvw3Z3oNhHgJYJPcJqJyOmi
4bmdtM3KrVDh5NdglUg2RtuSlkiJH8bzgRYwqSTJDCdmcnk7G3OM0FKWKzZVh1gLIIvUg7VVpOAb
0MjyfmUBLNKNRzlx0+Oe2RN1Vohd4rAu8E7NfVsnR24F9k7QR9UfZmt4Ub7ijdYa5KeXEqLPlFTf
Btm3a0rAtT4LF/3g9gXCFTC+tYbcLaKgnAFDcEPXpmEW6HVxtjnnCX0baWl/dDvnLcrA69TZ8ae3
IJzfZCCuev2sfgIWnpOWnVZ9Qu019wQc8goYdvwX3IPRwoTdH8dcwFeOCXqorQTU/hlu3qX5UrF9
NMzVRnJAnGtVUPcypULjli1xf+vhyCToNIoui92RGzpuJGp1C26bwB0LcKMJGSfYxyuzo7agHtMc
aR7yTQOnGCH0VgMrfmbKJmcX4aMQy42gVKJrqGwE2zXs2cZFcnlKFTq0vrIJUlnDSwzRhOmtImUU
9WRDfZJzOxZMYVC8jcV8XmZ9NPIm9o7Ir3kwcbNrU/q2oPfQqvMhZhRZUrOoL9esWb8sfrca8L6D
69mh+XFurOiRNkbNvaUNFepUDfXESuRVJvfBxwA4GY8N5G2+xXqcuXKvPyj/3DI7BuUnfhf7KJ7O
UMMoQO/VWzZRhnTl7Iz5LtmrbVKWjC0LrU4MeTytuKRkO40CBHnj1ch92JrYGHRneZNPpqbFmvvg
CyOPkhjyx6mjtXgphiafQTPpbprO+jgMykl9rzYxPJxdOmkNTeqQOuTX5oDihW+0hq/kHHM8fgm9
IxJmjmuDJ6KM9KuDthiB6mpa5byyOzxa+DuTUcHRFWMGob5aHfnA4UjMVLsZEMcilWDmMazt0XSz
qKSqyYo2JaDZVteRrP5fEx9q3kiw8gU3f9IqogE9DrEytyuNiIc9Xt6d135uFFuOFhB+iNn19iO1
jBWDcG+vMY0J5l52Yt1jmRFGtGn9Nqfdf/EXI6k9Jrsgy5ysjW2ahKCVPd5FCbQ7QPSulLnbIRSw
4EgmMV2VkHIE9cm92xqEWIlVwJ/ixSVj7PtI4errSNk333ZVEkulJxY6pSW5a995kjeYul+C4/ti
UZhL51uzGb9q9RTNzaI1BLozkA6kIp3I5M+/x/pl5H5TCSxOueZ5QA1+tD8XvPM4ZHpNPES337bE
TuPOw8wDX2+tc+9YRAnjmFKa2TO8WJxIdXCS8k7VmFKMHCJHkWL0lranZJNF9VgkvqypgRlwgZv2
QgFZ2Uu4ap/hAC4AJjuR3LJs/bcsVJ/4pS6wcC5gx1MG+ci02D0jKq4hF7upJi7c7G997rJuNH1T
Jgq+zT1VXZTw6Fr1R/TLpfA56/rlz5wfO12B9UUVZ2+lQJpO8J+J5Jic5FZ0VQoKHClqn6knAtLJ
Er8eYCbIM4nUjGo7GSLhIJbNa9++nRPSQyzmufpYAS54tuzJSTAdk+CMLbQXF8ZsZQcy0Mu3CYL4
MYzFxMtlVPJr8I1JG7XBHFQamyNEvTkvQv3IPu7vV16teaTR6eugN1uUHSyBZGd4VhfNJ9QTw0tb
1o/6kb0ZNgxMEp9g8a1pq1stg+xfhmrhe3pNxyVX6GfGCP39Lj56/Z0KfJtgDlGDapLLtTtSvsQ+
sqoZSWyKkF6VJvRr/OBqIVrzZ21pFhYkSN3zLnDnVEH0vT+1H+Y8TrUa+iG/sEkaNu0pGjVcbM53
RwZ/4M27QSPC2qHrEZZ6K8/XmnLPqE5zl+qhmniCfSaCtJdzzTsIg2PU/kKWnRMLjyaB/qDTxNVp
4rvhaXCMFZeOF1k/jPnCiO/s3t7LgmuSVCxeqMXG/ThzbpdJjerp2M3DLaXAMDFRvkCP+99WqhTq
rB/dDPpiqUGOhSLY4Nn8QDgQUxn7TmjOcilpAAJT5/itH3ct6XkjxJV1gh41DsFt6RiKtFdgpMpi
T25jQnPwC2Oy87SNzXSRfzG56Cdky/5z7F4ibA9pq9ka8h7h6egPfGQitxj/U8HV+b7VZlz5yT9W
bdmDxLAaEfJSg0TWHY0VyEEsdR6HL1/XO2J+5/k+dHN12gZJk+n1Bnrs6JaleCToIdRg9+BoIq5Q
JuAaP/BTUXUjegylN5qoCQMVohP/JnDy2v949Egq+kWoew4RoZMs7DGOluJGsxTm4e5tEs+NSO+V
lDAkqGifdUsvjd3FAaf+iWNsFkSiIAPLpcux+M5RZqA3Cc/1O3pilPeo3DAlA7S9FQcDRF6A+iMg
2CbAC2xwVgb+kFngfLjN2ZNMcrc6clKpl1Up/LpVQsMxv28rmuqjS/91vz4xmeSq5QBLOK6G36bt
HxUWf2iOaif9kwuU/eqO+3iA6j9qiyPfc3TmHxjI69PVtwStgzwE+iN2z52KhxowrY6Gin2KPvLH
l1B85mc3OfP+Bi0qvoWVO+ianiGTYsT8sumBdgw7BwFPqVF5xxByFKaGGMnAuer4WaXgjs0aDq1w
anFpnsQmWEcjNxh/ConbRQSiSPti4Jl+kcXzA6GvUqNje2zL40FUt2RrZvyFZQoA8Gl1jl1lYiJQ
O/sk/hLt+TLwXBH33x3IZIO85hypTm5EezmnKI2LKaM9Y/5hC78DGP5nAf9Hj2Y97f8K5Ea9RC8N
stMFnJvbyaHXP2X9BAK7O1tg6XLCrdKp8QgSRBGgNt7dge5QKhwd4fxsymYOQZFUIaHSqE5M7Vs9
4WKDXy1XFLoke64YHZfZWq+p5EIGMpqaIuJyVNEEHBnDz9Px1aS6A/sbb6SKA01P1VZ70SAfkyCG
dT12pb5CM3qMq/oum1QKn8BNC5jPPSQOslqx23LLi7ha6oqwbR/19TlIZ6cc/Xu81BfQeSi/n/vA
M8FTpSZizwtP+ynrtDNBLO2TRChrMSFm5RovbXIjeJTG67Wx8ujACyebV3GAx9XdxyT87ZWaDJyY
Iy66fr2755bJtSaLHklH4mTpESmsmCXS+lM6vGSbMLX4ZLLEDLIK0PaDbjak5slxY3z9XtkIWgZe
C6cypcBL4GqNWgsj0RqonjVpXSqDr8uyCvXqFbRftZaBQYZ2+3cWJ4OhlCWcGApvPHonIhpKb84H
fX/ViTnUNlrOmEdNaEpr0XLncLDS3ZPB4Na8Ttoy6H2RNzOo8xg2V0E6ZeBfly+/udwANU7wnXjR
BLu5R/dkxExTXxkmpZOQqZ1uuln3xi7gWqhFZsQP+qxp9b8VckFHpgJ3z53M6BuSqP56LkkOlly8
rY9xtBaSzxmsMVsksGW/Lnta/Q9bM9BYyPY851oO2+38isySSh/xvSGjG7ZjJoafQKvaheD8w6VD
blKpNuohmVZFa+kBTvbLQgdxSzmlmkEAoct+6wqrlaIGSIlHsgxRrlc9mk6peqaeW7o9JdET38Ir
jVEz9RlJFv6pTrDrShQhgrFdmu5PhtEyN7VYQP1Y6r68Ap8i9iLOjJ58ZlglnDEvRaHAnsLZSdWm
RdrCiXBV5bYTgZUFH8SWqnLgDmI9OHCgO4VwE2Xk7BrwNiWlMzQTtJ4f7qQL3PwyrZaKoyEt5p9B
0HZAFgdaQMjFM+q/lcIS0ldO+Zcc3xwc8kfLN0fuUZGOuo4R+S5wnhVILxlH7p7SqqEBWQbSTCvr
DEFgl/iVRGRP/VZ/7g5U5IOMIgFdc874o77PKHYB9/tTKHwgglr6Eg+Gq5m+mVLWmXAUihApvRgN
WkkYdQU/osEDRqD0PYJhVVZL3ObrF7S8v2WjLM6L3soeML+CaygViUvDdhUtOVWMtEe8b3wo2Vr9
b6hZabdnOgyzDT9HQvHmRbAE77qiRA881/UuxnlCddLh2gv37XvnQtqSDK0n5WX4x7rZck3pMtyr
tPwmJVpHDUi/pXJ6Yt81Y+EjGA3bngfNzWb6GRPA6nN6BqbkqeaayOtbDbd+9WWA3y7/Kkslz+Nb
TvHY+R1xBL/cWlxXCMcfLmIXKg2tzLszpXEDh7PkDOcJYPxOltRaWeQrNG2DTx1UhMfQyajKNrTJ
05wOHIly/+BLThVa8ygCWo6+D8SHsTe+N7H6rECGuntpGAwGRMQpsIW1Pw2/SU7M+x0R2urKoO+3
88Fyqy88c5PbrxP/cg4ITZRJD1ecQCQcQpH16NUlHZTCRXc/ZB+PYP70XzXMukCvOX6RQ6CjO5cO
eTPDwTsb7vK1A3qImqFy19D2xucyXaS62p1GMd1nIz7R1IDM4hNp01a91zSXXEYEQhJRDdhTISkb
h5BeW651pE9gCPonfKHYWGyNdEsYa+pYqyeXM6L91A4GhSQqelCGWBtMRhQgR6k7CQD//0iutgjF
HDn0i33glecZE8k14ybV0lG/ZJYHcG7tRdAXku979ek0RF+fd+tbuPEjV2FtRdWzA0qhdCf8At48
T1Y3RxFT0Uy9y0cKRwCGPXfmtWSBguyhIYK8ffxJLjHCLGB5hX1Z/lqoV9eumySu2YQ5XA1iu/fZ
EvQKMIht1EOp5lYzW91vqIKxq9yiuC+L1oYMbW/CMF1V9IOlJLBo25UgZxl2rm0s4k+E7TUym/HL
NtM4SV9VOusmx0kF9BRgk0fF/LHM7HxO7icbf5fdQPX0zwkzypKIjs1rLHZj7xnZzzLIsf2NKirh
WEjvrbmhK2qbH7M2zlsdOznfTmDOjn2EP9+HHjDO5TBOKYFHszM9PYwecL2T4RuGwdeOOZF+DAcE
sJId7uwJz8cyIY1nCyUd4BRMcSN+LBtNYZo7plr96WuBZj5Ty3D3f245lq8ocJme4V/pycfbN5ji
9UYRe6/W95Shq2FlgpJlHSG3svpkKRGLHQupTCqHMDEcbJdKVE8dvLzUlwpKiMo8cjz4mE6W4f0n
VERR1xtFiWrHXVGmQB8pJAfg2eXHZEHovAFil6WpwwSayQcUEHUBAlCOvSZgBOFB323Xu1V3dtCB
+4BsPDRL5Bk3vG8SOhItFXVlFKzPJW+YwVlNzlH2kXg7URW0Qgx/6X4m+R44mQmAjHI7L1vEgH0C
0Gj5ZIkVnE1kPeJru0TFzYdH6vkNzWFcVdECpEcY9/TnMwn16jEwrTauZowC7HNxfLZe1mUDQ4M0
Yc6dqaOKIIvU0fDu97mL12S0GDpsejOiM0Ed8b6giFgS07Gj7FgWWkF6kT9nXoZwI1jVSyv2XEZk
5IUoF2r0cDIXXuelaRSPrrWUbTaKvd/89ylQJkiGnMw/JMKDDHwg965XRNbjfb9QpWBAbQDwikqZ
fUkrT+HT31PTtHYo+muJxvVBXjYGZwhRoodynL9r1WmSEahQben+lMZIg5cOKGDKmKRDYFpl1mPJ
V3qr7uKqejQy4nsNCJwlM6Ry7vi73Eyygb7yQIHEHrf3YUVBhz2OZVOyCx0ZZu0manPInrDFU2dX
FjilVVBt6bLEjWkREYaT6A9+Rv6V5auCWnlaorA+MEZ+v5uA9BI2KKIa0nw0O/EXO2NJ4SBXSsgN
koiZasIlYILmXzmLuPYWq7alR6fMh4DFyNYWBST6RMzah1X76/rJ1+JVAfdUR/FSWBmI9Q3Z9bCf
yFA11KIw6q0jCSWMQQ2ntCGMylJdsYtlo8wriS+T5/LxG0QQCUPOcfPLqkBdU+YWJA6q3VWdi0pO
H0Zw/s7epy9mw/5eoFzLu/yTE0W+9TybXBye8UD25ZZy5z3DYdJ6COWF4bVAVezV5P3Osc7NIdM4
1AKcUn1MRxY8UQmYxANw36DF60QUYGK3kVbVWQYgv9kxKydqe/OIO0GuwnEifLgF3Nb+gW8fy1pe
MQhUeQqhucZPFymuB3llA8x60e0/GZReHy3dUV23Yi0C/TJ3U0me2gaKOGDYRSLkXDDgr0WQp/4E
S0hQLE6CANxr8toDx2hKpq5avJRZhh5fTZ3WoYlgDQL7/HzOZkiJsqwT7EqwUz+5YH5wj7scTKxR
4xZYFG600t2EY9jnwGuJLsuMztN+LKbTT0wlEC+jkEHagGXuADFbiYf4Zo9LKZvCFcBa8FcxSwTu
VjCmby0AKTqMk1MUnIqf+OuA59v60EuFMPq+rEHuUGuLI3b9ThPfVZN5jux1beHFFnwPMM7NbzKr
IGdfgaYi1ZH8f+rkTVemMYbqOjP6NSVp9RqkWmR6/N2kpX++AXg7dGN3qMOwI2jG4rQvEK2Dcj1s
yL/Kgm+ggGhq3gfp/kAENYmCIpKjZn2FiaAAz90Nu0opJUyUYBUtLFBtWpUoNbdKRZp1A9Pemr1D
gxy6IGlSxcJONHERROmiFk8CC2tp5LPGd6LwmrFKock32ZjgHdZ3YIVDVzDaP6hpxhMTaOzeaQuJ
r/3Yrlw5liFxv1dyqLslMYcNXKtC0J1c2+Bojg7hUec5Vcfd3d89OL6L8DPWiMD9k9dXkGO6q7ae
XcbSA7SLMSASiInQmnqA2dShWlFSXZbRcPg2OXInWvC7ld796TtEXr/M3rsjIwV/6qpsf9d11cur
Eh3Ia8ZoK3WVQ6A1NJV1FAyMVXaZcFq6DcRqdJwPSRgfEiZMhmfJWzikxBWWNile79vK2jR2Gek2
2czBcO/qCJWTyM+1hA5gvfIiJ99HWyT3JsPy62mqtEhKyD3rZbcyAgrMLLRzRliQtUXYm+ATj/ZR
OSKXWRE6MdeAq6qyhMxsdSA1nxmrzEeBKkS6SJVlpBz8d7n98f3tUiWmbNouJ4Su5FTlgjQ451dk
5PVe1g0QEB0QF3MFV36PIJUqJ2PTt5xDjx5yTsn2paN99ibvNZevl1Xwf0wrhdb3c+Th8EkwWuKx
Pq9vkabjwxeCpLOgCiZ6gEQ0c40Q/8YpxAyZ1Aol+reGWt48JJ01iA8KZFzsa2ZIZNxnIRysfxOX
ueqCv5TAVAuO5jkImcos/zHpUTkMQZVacAGXoEn4JYeej5PVu/UebyXHQTjBkOpFvMUWruk50oPy
ohANVcWXngh5imYKIdU5JVN8QNCeqP0UP6qFl2qhH/xsC/Z9yQMNG8xrVZp1lEj8eqB6C/YM5Pxn
v65TiPgXNKCvb/qutU2wM+BIsGl9CF6/Cy+4d/YyL1rqjOILLXYRYeABuqsmoR14dA2D+ZPFxXjV
vewNMNB6QcX7QeFUmQ+eUAzXwbw4kX1KKLHBfbSL9oar1elOd0Fyh1lfM4CKRmajjWm50ek1KrUN
x6tz74qY0jFZmg0iWGb3dNQkZlHQmaJUOc52r8PzpZhqsgleaIHYeun4CWIckdOrUep4PFHOL8rO
3FADoLpPasAILuB372QJ32AYc5DFkwibJvspp9VTnXBoJSD4smP84NUDJgmYI79Vukc55fbvjkS+
dxNRsF7IDe74zqKIwLEMgpM6MLUNNEroeZeQxk8QN4HEBTPeCq2JTRFrw9zxX5elHbXi1j8cwonT
tFD1VMmHTbqdSCx2k5JBaFfcKtMZlZG2FOsO0aKElN+7Yupxqr2bDk3x5mxlGEZD1dDu2smPazhi
qhI4MH2oB0TMmt6tQlCdTWvrv3Ua+e/oYGZHM3TQz9di7jfRpFlL3Zud7zcAGmAn7TTLOxloyO55
wGxIxMxznFA4vd2AbUBYXSLLzVhp6qZeDS+XGrrFORq0AKW6kTyU9MdfHczU7j35OvWpSOlqKlbV
WcX3YcnxQTeAcXUJcTVrXtvYUWOF4hsomi4N9YNwi7s9QPkw5Avf5KwqMyvNU5On2hI52X5XBWNv
4r5v+++yJe6jw4v9BH58PUQ9Qkleh5tnWmbVvcG5RFm3Ov5FFQLceuoHsYQ2HcilMSS7NkXgToSf
JZjgre9WB25aQVUAyRgzEMlVoGNgqNVAYS7RxBFR9NEPBhCMrovQPOAjTyaoARN8aGbyKqc8eOPd
Maci+CFS/6r0ci8NUk9jQEMPigAdCVb0hd5zouG6Q+kN4Qs7igIVOl6guO8DHxMGUYF/XTLIBcgg
C7fr4AOCs0klUcLfVqOeLnqZB2ib+8BSgii1F1Jyl1+R+EHpIrPuAwX7ZcdVxx5rJ4Quw3jq+4qG
/OpofCaweb+DrVLvABvJHg5yzQkciJdink5kIA3kCNps6j1fpGEaMQaRXKrScP8E0dyHDmfUn+tn
Tq4TbChA8BnhIBUvEzjNrtR9EfHItT0fwIn/NCJ5+Zv38H2cM+Di1sErZK5JGoYwll0nG2Ays+Ly
WXxbjA6vIeKiOAepDXsn3ELROXPMx2wPNNbT2ygWPDd8Ig5ruW36L1xVNkAw7TUgYMKLTOm9z8mn
oFcc/badylgR1NV7YZmPbtd73Oz249mMRS7U9F098Znl+UzELW0aV6DTxmVYW9VjBqAEGQEDj8fD
9q/yIXQU//yzS0NwqvCvlCE65+hp/ifiv2W+w/rkXTwCGnAWITPUuKOw0iwVoLZrIlRc2VJiVkj9
4ACvGX/SYaB3VkcZt7RkgyQURChI+ip1/lhZkujVrt8iaq9HNnqUsE0GlGR3Xj2+Y7a6VP9L1EzH
9jdYGwxZ+2Ev991DU0jABZWVo8k4psMPix8tgjdOzNSHI2VKvKiR0+j/f7p+vSO+6c3AE0QfUkqU
GQVYe4sux2uVMAzWPSlcPLBljEkHuFtph0Rksg8dobPjspexWps4XXLxUDaJtlYpcTIWBwcbYpnS
dJ6BmmDi3HPm5UkSIAylbl0g15M81WTUf9F6LA==
`protect end_protected
