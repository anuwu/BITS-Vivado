`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
grYpUA5jzoYp1LlWmdZ2ALEfyb0iZaBlbu2Jn5TWbislv0ePefGNtLrxAsy9+neVRtGKqzd/weQY
1GDOlCD3sw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jJRJFGl+freuRUOkHi4uiJXF1ZSDXCZnSp7sify5hay8gI8WQ5QHE0Kl1tU1VRdOD+ovbKr3K+cS
UqWpgUyeIHMS2fFsOi6SAu6Aoshxr0Vl9PE57JGCyWYxhIS/bFj42inspCVQCybe04fBzJMNWaUp
2qePZYRz32xbymT2jPo=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tu6th/stm+M5ynB/TKpquW8ZkolQD8eNSgYHhWrx1S0Oj+qDq3ifkyYP979H5aZBSsmi9nhkBeP5
00SMQNL9WZH3DTym/hO1AOEB/vZQ4iH5QuRFIKccEqDq2JtY6+UDXXKzO/1rIfmarsHX8ltlRTV/
zcfaeOmCAj7ywQc9UqYmky4qV8fErTo0+Sdz/lesSXUkxz2bi3RdkWlaTaVx6gglEIQd+UT3ZYt3
+UGswd7jIOxS6vlCnneyc3neS690RMPIIoNUnxysnaeZZUGvdfZpjktfag6rjQ59uaAGWliO4MMi
6ToA8bqievgo9dlWIHZ7qHH63+ZPGm4+ACmZLw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
anxX3tP+OSA4f+Zz3xRPWpNr0NFYOEkjWa+yDywi9ewNNEKmVmuybI2vuUNyxHHqdZuNWtw1fzH+
LvHMudDHSvrqUXO0i+yPr/b1uULww82dKZJhMTouZXfSBUYYR2R6eOUHlkc2mpuJW1b0Yfgqe/lL
U2cURbnRhzUDfX4a8/KZsget317eHUxMWntDUJjMnFKpxAe6rTs57ljr+47CKoyVApxpFRtXyva0
iIrl61ypfwevW1NM+dbuq0A2ep4qpKF3QXqu+5quZRKiS9wqmBIWbGIwWUFzi9jVuDlWbiy7K2/8
HWrhgAyLQfd3aizqZge9Kid8TFg/tOAzl3/Dig==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hfg0jhNUSwZoyKs+dkGwZfuOuLOYxt8dUSYFBsXNe53zJQUTW2+PTKtB4x0Xb2iLN7gmIGI0MkTa
VnwntAtFN20kw1KSsvMMJ5tmSswwrxvHJwEQEUQ97ZGqSWO2GHL6Y1M+TGniM4GhJ4MqrJ9nz3bJ
lDbNWHgjFGsf/h3qT5IiPslEewuncdt89+9yjAvcmXEyKAI2nU9sb2+Z/dYcbWohVAJhqZIShNET
j4MueDXbjuGAb3rviJH30Ms0ITe492AtvNh8bbtTcCumEGRwdxdBrBtudooM4fhp1QOulK1MlV70
8clOJrGF2872zCxai4LigCCBOk0uSW3ObDKbXg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SbPUQ56CmxNuuFeULNmdtP4VI25yIuTqRpQZv4fdI4ab2e9QChHgoTeL8pKVO9WcuhlNTx166GsZ
+J7LQgSi3dQSR++PcS3u1e//zfZcwXePmh5ndXtuNKSeOT1YlsZMy0NFnCR74oDcXIAWozlvfa3H
+Ha8zpAYNJlEcIxIlN8=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iBM86j8TSZyV5DU0rYA8Io0mzpNhxgzW55YqzBpIYOLzQUiY8G8WAdKhnnqwoz2tPjopVirg1TR5
tvZKebOq9UC6KFo7vKxpOX57N0cp4fFPLdWGp3bfCI0YVxBdZnmmB4Oc+YtxYdI6e+BC82GkMG6d
gVuqFuf9L0mulL+yXuTTt2uiDajwZIcjyq11UByNJFKgZWndCJNV+FkUL21qP0t0BgzJPx1vq9GI
Xcdhwmaqi5DH7ZSxtXWYHzXgMDV5w1iNgDI3RX7uYUR/uvXUFc8tvCukL4SxyVDekPuhO3EOq7lP
gm4n/MB66m+/WkJd04R1OsrCyFsGEkoFVCl47w==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TDm/CaHzF2sRlkHDDHosS/V53FzLYAEPesCrg1+oRNDDuRD9Xb5WpyqcNNNidE9joaps4c7lrYCD
3nRf5x+Z12x0YPF7kaiPnyDbXkFRv6Qy+JTaRUXeoTs54W+jPqxDrL1x6Wv9yIyFxShptBbnNkVI
e+UMuxDyxwcdq81KmTCZc+NgWtBB1VzY7ity43L6Zk/6njjEpAsUd275HuhcP4JW4NFW1TZDaNnF
Cww6OTyrgEG5hWZR86AzBS7yjfi5vJjN94IDbGHICM+1BbHZNAAylzDKaXvbNdWIsQbt3lRVnU+z
u9i9+X1Drqb7MWsOo8jYLXDlib7Gpm56+SqMOg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133696)
`protect data_block
7iPv+l449APEjqvJSEcJ/iUy2vtbwWuP6RMcvdjCEq+Ez9KTqM2oACcsSKnXqHsv+Ocac121zeu+
yIdiPJIuqi/50X/cbvcRh0PEQbQOL0vxV1NvYGRWriHoYw+zgOAa4J97aebig4hAqKdlGXID8XAV
aEWURwW8MpwJbPV4/lgWoZk2Z4xjugToxmufTuDeGhDI8C6pVhOBU5CE7GmQ9sNl1bgz3ODkw3I8
KnEwD1blGp9ZuG6opajrJeC2zVJlawj44FVxbPQ+WvhgBsHyg4skArK61JPqt7bayH9tBP0PobH/
H/Yfo/6Ke62nRLzic99MEunSAEhwL8yFPTyWxhk66Cigl4wN2Mlu9RrmbTITGYRL9lAZc0b1Brf3
Bnpj6Er8eN3zwjyftOCZFb1CTMyXbXapfeynpQARxIQkfApjYXi5TKCKVrGD0BxBJtOTmEJcobC0
00PWtOApIdNjHdo4dAiwWr5S2rjMX5LQug+umrup9p75KYVSuqTPLb/9MG5crMXrhyRe7kQQyEbA
Ju8P0gQNsMZ3ZzYZTtMLJhFnUFT0NkcmLbEMUyQ9T+9m61+4OqFmkP+6Y3lVo2YNBPSDEVGrHwXn
fRdH7edihhMlJfqGn6+joe8GUA4ZMIIxz9O+YEPTE0am1zaNdG9ZYj4jkN2f3YRa1I+FUeW2zefx
PuAxAnrml2GpLrRo64+7i/hdtrXCpnAIf5rE/lHNNNoem8qudHwLVYdePzTO6FtRz4SNIwYfAaXX
9OxIcWcikZm+9VmK7GbyF6hcOAwfN8eo3KDGqZ/QdfeB0hUhDCVp/TaKMkQqj1CRpER5yWmvq95v
rikqlWDexouc4pW/AkYegPX8XrUR6ESxgQ3QBZ7zZZS38eb7ebY4VRsxJFYNGPVRiHj29NAG8s0S
eXpo8gocxFHZqtoxn6LC68prEHA7cMqhSr6DWNZftwx0p0DTwsZWT5HVS1ApNyOLn7JbJUlG3CUv
RFezMAEGIMD2SzvVezI3e5jFMWYoLnQbC8rOvcMSY4efJdv6d4UbcPRfb00uFvFt9apP19g4xaGK
EAXAwJuWxJYOHS9wcMGZD37hd+TYCHMkN1cD1CHMPtpXPPmN1QYkrnHk3B6V/MZg6YkRkeS66sjx
yIxqUbCWodNFcFnexWQVvVy0VG+Au5OmXO91eBiSsUJj+xGPcIkkfjKVCsr/g/EZJjzhpxgayb6b
YT3KLYOLiLhU0qrQ9ATtUPnK7CLuJhJIObDjFTHuyxShOfcSmT93Zwm7bEkHGU6buAvP2ENYg2jW
9eSDWd1U+/y8y7y11ZdApJURfDr+TSzzNbXnChcd8FW+pIQcyPkbGHi52/g2uIeWZmd3XaFTH1Rb
FVejz+aFGHJzpfjK3FoYc2hNjfH1cGu2iDO61O9YKKjqBN+V0znjyos9ON4qQ/M0a1cJEf10SKYH
FvOCwkpOKy2HAOI8OAQUW3GypSQputIREn5f2CEC/LtS0LIIlpAIvRbgXd7WahF+WEgzbHB1qFfA
ykYIaQyISkx1nQJ9P8zJK9jiicpLEjvPw8rPBC57Sm82zirjKI7Dm7wWoHmFpJFys61cRavvzbxS
q4HNm3rtLJxIVgw2bBSjDTvTjgUTYFFBbvNBbPQMSKJEN2FDRK/QIDExeZFf2PHIo+6ZwgdJVOoU
cZyE6CnpExywncolz4tfI/hobaR263uBi2XZg5H9xaknHnyiZCt0dQer04Ddpkit3theGuF0EP3W
gIujGIa8nd2CSeQnLKbp5+UVkeAAPbXDaCwPGnrw3LRhz8mct1kdXIV2clmpigpgMo1cTd1Y1P6H
mVpY0icBquiraAuVtRzYJTIFvz0Z+kHbZgsajKS1l0+c9SLUXKnKwkwvehgw7ASvyNC3KBx8fWKZ
hfkqOo7MB/11unF3fn6U6q0tYruV4ulONdXSl7PlSRznNgsihUaLOxlaAvkWSMDYB4FApsXvmpwJ
ema6Oej43loC3AdfpYtD67oVyMH8xt7CfTIfptocDFg5WJg+HWOU9IEyI7O+/KAnezI9hOBnTCQ2
RvRVNvo6c2kgJkKLzNmZIs3QSC6RvgBejwniR9UYP+ZipkZrPN/cnBuXWOtgKDbwIvRBEn81PrbU
rCXXvm/O+5KnVGkFyFXpO3mvW/c1DPlLyBLmhCBKpUBF+gW06Q4piyQ9I4M37x0OFcxXwgo2IEFR
0EzUXlgApK8GliIh/0GKCFCa/IyfV15Fg7ZhlLiTrI0CX9XHoEKXnxjQL+jGI6ccoZT9S05rKDJy
Jzgp6jz+XwahX/WMXx+83fGJqp9Mu5U9/eLbmCaCF7+gk/a36krZ/CekFCr7V4iAGjT3IN+DGwPb
xaaKKF/c/9Kr22BnXUkUkrXWpN/XNljTQ8Eso+HDGQMqlt6+NIZ6UPlGe88VBKUmXXIRbFMbfeEq
XJ3CtoiSg41vn85nwmMrq4aInMVZD2Emq1QSEs03NWYchCa9WwZYykA3PvlarxTrmUt1Dw8gxfz+
Mb+NWJoceBmhmDrc/1z+25Y9OAqV5QDypMrgZqtjJ1+Maj3k1HOpH4PFwbwAN9FQuRPX5F6uV2NV
FhhUW9UPdMhrbuf+VA7/ktNrpGL3WHYVi8IOtg43Mh/azdEL8bPRkzzIJQuJp70FfVpeTszq2Fpb
A4SdghmcYDQ3i8uVfz1Nmwzofz+u+XoO3oEG/fNlQSeS5mTtN4p3aGPWUIb5sRo8vvm/pxo8mtUb
zOEnav+KEmFsr86srGNBWhHerPqanMSan9kqHm4/9h+UaQU4za3pUyCYBv2Cm3jZM185r0D7daKb
uhvkSq8HeLgQfGKazMvtDbY+Ij9BvGGRkZCcTftciSn/uvEzH+UeC0PK9V0rZ/qN20sfAiDYJTAs
E4wJGTggmBFkoh1qV/1eQ88Q5zWe7lQCGn8GPB2SriRHOjbCRQ46hjGr/EcuNVNIEdqQCtMUiB7I
5Fb5oFPh3R8tl8FOWLfypSNFe9UtGTEk/qeVxQgS8A11lePVNNk9CONFJ7wJOPzx3ARcpcPZhl3l
dQBoDiG8r3kxFYID5xThwBZ7JYV+tq7dy4U0tn7UBu0StRAU6McIC4f5ZdCVUNEuEGX0TR/m1xi/
nfqbJLg6PJRI3ws4imz98l4C7h7kbKb3qtCwCK7w/jcZf5WYHOKT5/btXz35PQ9vcOwOnH+IazOb
neIegIQduOOwa+h7YGO31gl+o8972jYrrdJbXr9nEb556Pj1ykMjv0cM0bde334YP6kNxQwrgLX/
p+pBtH0f9WGUFshKP04m6VC1HlUZAX0l+eXLTTnMyftxslflGV2q2dIYASFMo4To+G7aiEvrorFx
CRQQS4IY3VfkKoULqTKlpcATAuIVGBX0GC40S6HU+kIfiVmtheN3tSe40wSGpEz1OgidlRjFAOMW
RmLQYR671LsNOoRKRh7mJ8U+MQFvKGuxj1OkYTh916B6bu1hJsEj7hq2JTp4BJ75FkYW10Mw1RZX
Hhqx84jAjO9kn/NfD3Oe83sl09AdwneRO1MUreIBnWvQxpIn1Bhf9wDe7e9xDrSb9XvYP9YjfGZ6
uasCl7nwshCjViwBqjSC/aso01vBGcE1dVFSkiX2z3Afb9wwquLWN4hN2piam2CRUZH1+X/7uZqj
/zyT79Nwa90a/i+YfuIQJs5/OgmqO/pxBKdeyKCYBbP6lguiYOfrs6bt3iq6TiW72k2L9T8zOaAI
zJsK/S0hXdyYkyOloNp0lEQtP6m+vGV3BKNxiFop4B2VLSEyTJ6xuhR94wE1/hteJQi8VcLGQTje
FMPJgbQ1S50Rw4eceKLqOdODbbmHy8OBEybHAZSrnlkWvMyAl7/3vAh+DpCnESPqg1JMdIFcR/lE
FNmfbSJ5I7nGlYTW0PaLtc0M0ePruoK1rASs6f9HXBzh1iTgDYiqalZz9eCr1e8DD7asPrVnBIik
EVUloUTkKLlOwRaiI1dyj1BN0PvVi/Jbnmm3TIYm4KneVyhE+fD/iA2WUBF2nlz6PBJluh2GCk0z
v85aF8UIQbBVSd6LiWIkFLzHef2XotpCmAceemMQUMzmjXAa6egdF0LpDIDQakmeY+t3V7Una8s1
kghlJqOp92n7KNxh2He7rbAmZYkWilpr94t6EvYfBu/tj2V9yLxXF7sFnVjLwh6VAwjCHrDJLJb8
pVN85vP5H0Uvrbgy9ZWTfSSmlsnRKOdDCXIKnwxs+WPPq8phnrMwBwtJTTqEDMA5hJxucTm/Vhxd
+XRF7IPLoGkfSY8RkuLo/oZo7UzCD+ZKxG/c+v2dNn6m2AW+do2IMzyzAcOwtBw00hmYt70L9KsB
R+3fP7kIZs1OzhaqcTVOUFY8Nw9qZl31v4w8Z4ZkhrVdkdffwiNEGNiLPrfdRxLCx+Mq0zq40U2e
2OW+DDEvhJglcuI2DQR3rMujanLRWmDeKubWyaQ87d1w4tycGNImOoWfodAUUWM+QBAKytMGiRFl
AkO5BkXmevC7NTqxFKno3kLKTTTUP52Gw9LlemrnPkB3pd53AZSpVqEvmDFZynvZJv0sxFAfxOfG
l+YjLP6CKAi4DVb0301RA89wPrbrqK61zPf2ZrINE7CwuEGc/gbSu1O2PBP7Jpr7vGS4iEyMwMQn
A0SUHxDDKp/E7jDqTFwX3XNDQ+8+DjIPKrYG5ByFFXB++dq8RXFadNFi0ezh1eCwYWpmtkFvh+y9
IqZc08Df6K11nBUXz81jQtpbr8qqid/IXXw5sg50JfpA2brEKX0U+539HHSx0U+oMf/wZl1KMFiZ
EC5UTHK57rqkOBHU8kgCAdhvNNI5V70sLJ5eqqzPpgjs6bOepOCHHE/BOI1MKYd6BEqmr8cOxuRY
i/AhuUtjvpJipIAh2buDJOre1fwN+4uLuFHWdbSEKW1lBL7Pl9fF641yz5pooRdmb4P0r+syLnGf
es91659KD97DFy55FM9nJ23axGvh/qGBd72z76x6r/6VAKwCOz9owxIMIxy8axS66sv2AZ3ICXze
+InXVTeNLgasbg8QYbkkpiN5vRXDnW8SoIDSNlGJ68GfRWPYtkoHM2WSeV4FT1aOjVVgEFmXVuWm
KMiz4UMk2xbO6Y3TVkaP5UuV7edihqrdHpbfw9k9JkJQ+VrvcH7cboHUyOXdiWZjXWuCHMX4WQgQ
NRujS+O3+DC0aAaMnYke8fVqGKV1NE51/GPcHpfoBuCPJb3OZfmTtwfkdPYj40qjdhGGj0JBGoJe
QmCR2z3q0UaUCG1SnHWEUJAlszn5BjpVq6JOGHVJfK/UgM00VMU7TQZAbDhQ0LD3y7Qnb/EUOIOa
xthf0z3hwu3gCLXNn2e92rIGQ8jffU5IymQCzrny5vDsX8XRFtqqtXt0klnoZMk3eUePfCRmB26w
d891RXdDsXmx0qH31le/eBgqzH6XpL8CRPwDS1Ct3FBMPQyY6juaLsfFMJ5WhGsN+JF4CzYaD/hx
RoY0PjvB2p72+H3RADJk07xgWoHL37jQOdlMwoK1DnPoAqFQMtJLrvq2BJyza655NR60/E+lCEke
q3Cd5MgiTUbb/RRwgQI/0IbKibrZYMuI8Jfj1dkuO8PlL87rEZHTWZFANvj8cndIfiw/5cMhYAod
tZDefxqULGHENtFXzZwI2nP5O1EAVJ2IeYAmOlrvHkpH3BoI6unNg/BIWX7HENHNutT6CtCMIHhp
TdbwY8SyZIOjiyku63SR+pzg3k3URH7dE3MR/3efl8WKFl/kQN4UOTjo0d2Z+Kwrv2LP4V0Rv2Kw
TGS35cEp5lK+OQdIggf3sJ6isgfSBaMDnsRMCWwCv+coU3ouy6m+5lx8y5lPIyxZb7fo6omuCd+U
NPHZIQdNhOhwumi4N0ygZZdhWzcqCMfKIg7TR9cU+BCcjnlXEzNh08Qb/JEnraVdq3E1PyYy+4NJ
RVKUiSOEi0LRxMkOFBDsdtp1Q904eJQS4Qx+gy7E18JRPMhVOwatV1oPXYs58vOhH2g2aV46CLqI
uRli3yPUM7eS3O0dt9HOvoeNTXK80nYG8o8aPRb+s9GwZBVvruHMzbRhfArfn9B0jBbdbVEpqLOq
EU4t+im4IxyHPnDNEp7I9eGJyABMEaR2cGqMFpNSo5p5dFKIu7aRObxzDT1rbG8PRX8j22uMMgnG
nw2WJo+94VxM7DLPgaFQ/+bexV4m10x1APfm0f5juiA3oEGPLNgeDKY5yH1NhXZhjYHbIl0JVSg/
Ui93yj0JTiVC6QYP+RHQ57XSfvlYsf5aZs6Ih7FEypRhSlcpEenmU5HjWPsk0kDo5Q1AjLS4V0Ds
c60+6HK+NSzMrmDFS/6HYtwlxYOGnEPyKcIjXB+IP1zScJOTg5bEzasOeiB0YrNzWakZNlUJmRvX
s0pSEK/ncr8k/CSkni4GCEj1zIRGWQaFARYZ5MrpLcTV+hV7H7MVXWF7837oia5Vw2BXPspzD7Dc
3+39S8CaQn9YVpwr1o1lk9GPC/bZQJHuayJCb9NsORpQXY9K1YfdysRBLA4esyxrhg+JsrwRzcC7
lpDWkvtM3bZdXsyh+7jyxpkgj9EChKY9ooyDs0Wq1PiF8GrVLFKSn0dZf3FCUqfglqQKuyENC3ek
cD57rCaZ+MnlCAHDvvvPsIIJaJ/APNYTe+Ms6nwQQDU/tbtHA+473t/7q6IEuf4DjJxXUNaTxvD6
ovKkkxIC8VTRUqUhGbw7NOnbhV0DMhB7URJsn2yzDT/P1U8CF9e6ElcMXbl+BY6xoWgNJZ4Ymetp
GC4aOk2RTkhhVvzwU1eMrgmFkGfGlPBtxIPlREcE/ueKwEAaPax0kmGQqUceEnQwd8FP+7R2HD/p
U2qi6C1Vnbf9baUo2fsvz/knixnHtekACQFSESm/F47GmplGuXb/g2P32uqb+HTmWmD1arFMBpMh
3omZVP+Ypf3ehJai9Zg/XiK06Mka5PFEzVC5eKl8xOts0/C5z7ltuigif/xoJ6GTcSZRseqsp0vc
DpxrkR12MwlksH9+2VOdiuYFVgnKmdgIsyaGrs/3rxAMZCvEmYZJDu0OwylmVVBGmoY3euHfPAYj
iHxueKkD6ko+osLvMPDXm0hiBiar2LzjPaBcJj0MhqodL7l2eR1TmKV6I65Qx98bjV9FmO6KN/uu
aGPET018HuL1Brh48kvhhg2pv5Of2VhQBOyOV2HWn/WKKb9LZWPA8c+r1JBJYayIg4V0vl4EaXGZ
56US+WuwjMjEnf8nWRI0X+KhfK3JHofgNLnDjmjl4M1HVhYYqtrQU/CzW+kdzireYDHQvuq1giho
RrkrX1e9wcekufowU675Hy8KFVoFGNpJ28nfT8hiNnEBADYMrYWSqlg6HNuihcQxCpz716r1mEnk
BI7KkUdMSLiBVzUfOFHIEdg4YHumIO5POk2kDk/jwTGVVEjEv6b0MbM6du/mSrGqE+EcUjnnaIyZ
V3PKi7svC4RbvYmill3yLwgWh042JngGYRMJigsjTjhlAoTzJPEFE+afAee5X2ha8W3+8YjlaWAF
tcRCcXFj9nloo39KWu03oYoODrLmaI/mk5V0ZKu+Fr3zb0zoPaByHjiObpa6zcvura33GNAh1IJt
0Ljngl4VPKoTpB714HWTKrn1m1bZxTbV9fkn95pMnNd+nmd1WNaBy8cRlHyQUQy313kZlhmLDxzy
rqOJBAKEnUo8t3WC5LO6KM+fvK4YmKMqkb2FIBHZYdoDs/Ih0SlfDorBZQWJkV/kAdHbRQ85Bg7N
hep/khcT3ZyyRYJW3Y3QkabsDWJ6UWz/w0c+DyQuLWNteipDu77sJ80zxVSDWxw1uR4DPSpy59Vo
1Y6SO0Ff9gE3Ar68YPsn6WTzUWLkaalTDCQHZGemq+k0JvCS+m12pKQ9c7Xy+dCdp0P3HCSuNy8d
oa8v/eGtd2FDLbVhACK2nx4uIa4UjZs6HJ8lFL4ojdLM9BTLUWjPjrlA3ACHOTssYgfB+lZLAisd
JOxP/vvkF0RlOh10XGaa7IxRQp2EjP1E9JYZyWjifbjk1NMY/74DUr5F2KIDKAADSd8eqKVdv4fr
XTW7NcJZ/d32hEHwizObGz2ly/l5dewf1r7GWsSFOerQfqo9oNb9/E/txHjzbcRZRNYFyquD8zMQ
UJU0kLyPYVx970z7yxK8kl4QACKR+CQo0twy9yKEqmbftXYN2+f2jEjOfGpGycnc9gEZ0rnBM/Hp
KMlGK6ZDtM/FFvTOfoySZcshcV8Li6TGu4iEYI7UxknWPUyrDdt9KeX3Vjuot+zavEpYmdCp1eYK
xX3ePh56kCuh+xgaWP81VP3/M8tj9B04nsVAUBOby1//+IpaosduNUMBRQmgznODCurdjEDQmDdr
LJZTUImVpEwu0T4zUnLxqJcPtTnCQxOrP4CZk+O++Jtgh1a+54HHHp7CrnbVAdiDkZZqSgjjuj/U
PbUETOpl/HdCVd+E9qhhS9f/MaveB8kuiEAsYlZpj78pdtbQ2PsShpyNvgitJ3yTLZugmz2HO4UQ
NF0icfCka+umJPb2Zs4p7eVB+muewo0MbsXJ3EX5TV+YrekT26DQnOEuaCCytWxfe+FVl88U4zMu
MS8e/cq065MCMY8j+KhVc5H+YOZZdjIHFLeKR8RSsDfQD9cAy0TPyYfFWvyTp9VbP+PR1PnVYeC/
aiB8jHSEVpSoeIDh22SNI3QqOFR7EiiTFsa488fADgYfBi7xqID/syVoMqvjgiHcFcr7CKHmhLjT
BePmSKg3JflCQcXlqFeWLMqlCHnofDD31Y+waAw2aK79KzIFtJ1pIQOymQ/WLxPYafH9o9aB+pzo
oVlSxxQ90mbGvL52qCvk30wG+mIDL6SK/cggBzK/jj/wHD1zDu2uhXMJVTg+7CET64fvDSqgAMQS
6XHjPaMMUEgZw9uFirD7sEJES/Gm1nbxuQtC+zvrxK2O1JnxIqdQRzLPotv0geuisBV6G6qWIubn
QTHF+Gj2rKcsg0521CPjpJiT1Y73be/lulduV4OYiGFdv7qrTPSrgp+IBt7nB4UtUSpdRmjPB6Km
MKFtxNpmgFsQ0KgE4B0b/QuA2lN2UkhhGn515Nhzz/nanCsXb37/T7RRkQjkHTGuOtUbU+jIH3xv
Si9rWquBp8gfKdiNtAlQy8yWRDaGUNxFopHnH68NRMMlf3MZ5jIYtqrkB42WjBDG+uppFKd5rALs
wNosyoQDuPEZwR1RqB32PLA5FBP3HLCdjFJqfJqsuYtjqIj+DK0RtAdcSx/zGdV4ydCgTKpTAZqb
0KMWtdeOLljJYg0Qbyp+ils1OUo+gDIjbLoO9sVojWYo6Krq+kE2xlI+ICmeXH4+9yw09g1XGh+O
fEzCWK9ClZqhuVmlaaLBlaupezkRAEBK7zQ31QC7b6kruw6IPIR51NO8f3WijeU14B18oqKoebXL
HiMjoAqdk2KupwnTaXSF6wRQML1XD/QVlmE0IThshDPGkOXE49MRypLawCRUAlfOFY7YO1cHTlBT
o3Cl/+e1od6n+/9FVuoROvZ5W7s+K4EG6MAN4E7O82DQFPWPNbLwXJt4HALt69zndQekIQohGoNw
093JX7Df2MFSOhcz0gyKuAOfFnrVjm4s6lyhMcRKNeUAzFGdYXIL05cEczuX92CXaFxiNAvTEMuf
nKfd+ShtYhV+9DB7ymwW/ygtLVAAn2ykGroc0QGnbTqJF19vlht7AUxcs3OulowA134l3FqWqwhD
P9anX5Ak/tfZISpAK9M88+c/zLb1DeiiqbRBWvDy02ril8mI4Q8D5J36Atg4ZTGOU+yxF4TvBegU
FLeLsgYGQuoTfm4Rl0OvW7yQDztS7PAlBFe4cZVWif6/5M429ixh68uynfdEiiEAtb/3eyvBmRgg
qwmBCAHyVJaW8PzCCDGqIzYTwdfuycySS3yzKBlQVHUay4wBgxbMrNkZgrclTk4QTtWCWCdm+yqE
g5uAzqkAh2HRk5MKSrzM/BHEPlLGT19irmFvAQ7UIhPMoLTp6wsjDcIf4llMbwkDFuzX74fnGDVe
hnPvZRNTmXBzqQp6CP98i1pBoBu8jQzQmtCS1Zp7mjARvkfL8ekStFbC4gixdFnr2QVflIu6Wi1F
eR+uVErKVhYwmzk4hShoMUX5sXSc7s1LvEwM0RhC2Ap/ts3pm+hSVxzA6GPhfPwPDhz0FEJtB5JV
0rd2kAOirfzcHXgV1IbdnfkrO20MDoO4oAzijdqUunROfs96H71YyAzpdbW8N7wleekJhnCv/uwV
RCboqWZQe7hFRPAQ3ymgNsEz5N03ge4hsIYrnPRQizQI2fFnWRBG5EezKNm5fmMeBV+3w57IS2oo
dI3EuGunEU+/lM4TxcWrAWTPv/GNmcFntyVCU9woTJXZwR/0Rn4pwxJdNWA4e5cv/yxFfWU1Qy9v
UvquInl+3WshWUrOKdwPd4beIaCqo9YWQBylfi++IyEfKWXe1k+gw1BeFKsYFHRhuH1O5V7Sjr8X
Re1iAUDABa0TqkSdrm/ytpJCHenfM7GZoyDzFVoh2apG7I3cOjXQOf8inCrFvLyu4LIz2uxLNrt3
tRC0k+jd0CowbWkH4svUtD6YnFvqSGm2BOvXUxLw+JIOLiYh03H6uAfnQZ5NFqERsu/UMfCyNw+M
RuPK9Kw+UZAOX0l4rWuFzPPjLNRo/oUtRaTLRxvm5a6l9U/mCAcnranqMzJ7JcXJ7Tbo/+OPRyua
nA/0mRsyPePirpklwVDZ02idJYL2St2YxUwLn8VKCKJ/gTpm9ZqD+rHEf725fWKRviL8o9ShVQUR
XHubdDZMghhVi4ESdWJYIyedrr5mZapVPICuXRUACpK8XTDlaHSmixtmA5L5xdd6gRWGcofJ6+SR
RSZ6K1U/j+deTRfmzjerWIWS7Ydx3JOJ4FpdJc9oOrzpMdQgO6UEQod1IhxUJgzsMJdM9pGxF/yH
ZSoOzxPhjFpz6jLUNqv1j7lIVbv55k+vhpjAKpL4MxUQQBT5f9bIiDmE54dVUJTYQSrlCnbqQYPa
EE1gpNtw51GRpKZHjaYjw4aFljUmHj4KzlP4t43IFlNFtZ2MscrSMYOXfjEB5cqxUEicHA7jBaDG
6gC/kqOUYiKmtjm1pZ42C4S9wRZZOd43putFBwTEcCUwNausJFljaP74PcSCUXjX0gZDNk4CXjFy
2OHh4sbQeLgMc+XROQgXuceVbgim3gbbjy12Yb1wtsSKlDvn0HNMQJFwwwfdSR+pWoBqJo88rKaJ
fvKjohs1DLQ7f82VO6d+59pp/1rR1T3vW1vOlEhitIU7aF0/YGL3LX8mLfYkVcjEmHLRnmNEC8cA
faHgIb3k7Pcx/vyeP6GUTeQq6tPhkIGxWeQu6hkVucjyrvwxkKGrCfkpqtW+PTVJ5rY/jSBB8aKv
b4njFRkV4CBQ3GwwHJJECj3jNAEwxuNq/qdM3dYs36JoTz3FMdeOwSwJFIsCoCT5YP3fT9sxPoY9
1+uQVeaZ6WHeLT7DvPT/DEy8MXZynJ3tPy9jeQcsVQY4q8X5T+Wub6A/ELueS9BjGWYGO3Ureq6c
cyb1g6T0+9QlrRbR03d2KuA19CXGVvBDF3U8tnGR1WB/jHGC84MPy7b6tknS3YRtMmH0TXKPYGrG
yDlG344xnUT8n7V/sHM3oyvFjL2CDFv6YFyHSoyVVTmKZbnVoaUvpXEDd7Mx8EYnLOONDTKHYGbN
WQijQ/mo3cwaUJQY6I3uwsxbultlTXEBTLLR2ksLhTt8UHPUezSQNGPNVgzuYObKsRHVo+pMGUOA
kdZVpj3uT7U0+cJUlY6qGyjkQeYxGFH7dboyGcgseKEFkgo+qnQrODKU4mdul8Sd7OyZ1lTqR2Nv
M9fvBWrRtXwYjYibSfT5Lj/ilreykgnv+VAKNuxklJko7c2M2GqC5gIv+t3ovBjBGBl6Mq8d3Dd9
kdGm0yWQTVwJ76LtER3oTk7az14Z9hYUIeLftsiR0JRm+8uh/lD2lR3g8K6vp9umskpxXR/EjtRS
8g5FZUX9AzxUwFognlLbxZsnkJ3J2JNS+gkC0xABOJbUydwkljOKsDUXO+Z6T1FpJBx/dCfqdGbR
9SvasQbM9X+aYvuP0Gqe4ociVveGFPeXomTE7/qjvMcDqZV8aUYSvasG4ZRqW4VyWTpocYI5prcO
LFzjq9VJW6BHHCPbPVrSc4LNeSnhycyXWZ6TgYgRiqA21CmLZpAM4eKGOjZsuw7TCiQz4xterFDJ
BikAdxRZkFBsccFnJeHm9K45cXIS/LeVBkXGSEgEf2OwCI7dmuM5iSTdQIu/sLPFr2YoxuPuureW
6SUWwpmKM5XbAmuUlrkRaA43zdjra9VC83bGSc8lFktL/U2qrKNH5z40LGRp0IinABVAFSwgowHd
OqroHpmgeI5BXnsIH9F9ctLj/uZArLDxFJvRctoQYdzqf6i1t/RhAXtuPD2JfNXDdjyvNa0u77gd
FQ4YARvGgTInoZyf6RYsVYOUPlm/FGHkN4siT1B+eU9oIqGr8talLsWMibCnOSs4V2y3N07AhcVG
H1Ta4b2w8n3pQyyTLDWw3cFp3bsDietNRx87LaZFU2Hc8xUd3wj1c4PMdlwd5w+nHJCbt8pB0RQY
MtW4OV5fj0UOSQRmpzBNFOWZswNEOcbHjNBlYxFPampI8S4J8cFlrcPA0tQ9port6pIaokZop8oV
qLyhxxBip9GBoxZGbBq07P77TtlX+HzXOoCCDHW70HS0mImFyATUf9CH8McxI/fJFvKm8qUdMfpz
aUlMugnC4rq1DZg1pIXryYnSJrwXbzaV5w13HV9NVhygbLw59qjasYHEMIdCIR8t04od/ELh0ug/
4sRACz7iF8Nvvbrj3AfWbuFZG3gMqV3yLHVse+Bw7rlHo28l2m82a68JHXFFYCFL9HZo75+nC5HS
9Rpa9GjgcTEvVqB/kJXHDf96DXmGjGRbp0PZ4/OF+cjB76jXD+JiSFPPePA7XAhx4CSEboZj2Qy0
eu4HR6E2A349dpnVTuzsWnmvtKPN+cK1chkMFkkueUUOlseA7hdtitm3uoe1Pw7vd/St7I/X4cK4
mLcI5dIbIbGGUdNCUmyBubjKWh7NoDxWBho1lR2NJrP4J3sZcq9pdTo1q+EGFouktngEiAKWI5gi
xhTjV3uZTMd1DcqzvADlv8ZH8oSzgDnxfc99TczZDwxpBhFQlSaf2VuCRqPaAeQmVQQXfeX+PZyH
Zy2DlUPxQiHQEhwWjZTpOUEjU2Z4gs71ItydMIDWQUfE/+aFThMBAELG387yC1U3dG8E8OzPtcSZ
86y4eufqoIYtEBfo8h4uJs6K2KXMuuGQI/fhClscRkvwdvUtRTJE18hu/Kzc6PhouU2s7qwsOq9R
4BLRKiEF0QtqTWETLOO2M7Us5R1n1VNgoyp59ZWV2GLhRoLNXCQ5oL9T7F+8427BOKr+5oiiyQTf
eroXAc4w8PAvTGJKUE8cj9jIIhZYCEBDtXr/n3cRfjYLbRNMGL51ZMQW0hyBgn6ZgyvcBkHj65o2
+c5wLXB+eEDix09Jc42PHNV3AwnFRXostaJBMv2tqZfPDtA6ENeR0gge/E7U5obVfKz+UmLGzkea
a1bIGiqhDmHs1sBOKK8DSEW6984PrCDWhp7cR4IrEVLDqJMMqZsPrjf22qHnS4ML9vUQSG59rArS
s5ACdLEYMe5WtAHivsdV10AQHDUvvg5n9oExYti23M2MKnqRIKkmiwPk7/rgupi7hy9qPMHL9Z+m
jhVTp+ywZluOmg34tXFIYouu/KxWSFNcIwnZEaYczSUKTPNPxn/WrS6K6Nj/DuNOXOA8QGOXe2Cr
uvtZak0iZTUdOmfpwkbN3Vzhptl2ijEqua+PXZGUAyQsLe3H2yXWZw0p+rvT7Y8NqEpmsuu2ORiW
U8/MLPM1ULTj2hD7U0qNiX+oPCLBixaBUUNmch540RaxKG/aNnBtx52y1c3prDj7ZNQUBVIUucw8
1oOhoGbgzBjQf0to/gLnhic33FDvVye5S6/POPSN8WxdoAN8fS3U6JwVGgb2ZpKh17OTaDFYZ/IH
ddUv6cmgR1zEIiHbuq2ZxUuqvom/uFXTh3XDMwM0CRN0KyuzPT+j28/umyA76W8dI9iWj65HPuXc
FUe3fTm1+Vn3hxDS0seKG/qMDgoR8SvwH697VsGcQnkY8AjUJmPP3/jHtuIVy2cVu+dtiHfF8R8U
3Tym9Anz2OWAQn2mGv1waa8bd+tV90JRo+tN3dZxon4eHSX6QFUpHnCrOmH/2IP0I0XcSpSitJ0T
gBGOkZGTzyYe4owzIHHse+UiUro2KAIG8cV1ZmU4rDtS/Aq7lDA7vuPRM02955QxkBIAGneuPSv0
gqjrGC7+Fxqv8r1DPmMxmyi0KQPm5wB0aQgXplTK7a6F1kyRo3b7ofH5OUCLpecCfLoBIFe+IJKT
t2VmLpSna8f8Km/+6Sfgcy0VrJkx2KBxPr48Dd/UVeTn193GYFqbpagUvgeFCIXcyIha/W4Fru2q
aTEkneRx65jsHA7nBJByV70jcciU8IiRWNvsnX4u/CRaJpUjMwNN6EuiAf0r26ZRDPQ+PjzOU4OG
ZNfnrDajjwArscCUdTAitqExLm8ttNWdDNSP4YOYBqQ1Ade93MfQk7/cahRnlpmmv5vzpxtwrjbT
95MetLv6hwFhg7CuGYL60lsD7iTG3j/muuR88hCs/9IpQUDEL9x13xOyAM2wQoGdYbCLoVCVYRVA
jGNePAJPy3d5c7Pk88UQfTAwtPA0tU/3g3bQBCyqsGreqhZH5DjodGO017lNoSpjMotz9fN6RYRZ
uJZw5U21s+yapCcmejeFoR38VJQB4VmFSvBlwN1HKV9kvfqRuLwLVSqIXU0XvtoOyPKJJeBEmyz+
HbA/DybLHanO2CDNLc52SZqyrnTPXWJNQc5qWVJvdngtk4q75XKlO8uURhFMGucW9F79+C2G2RG6
axArygwlB2f/9XicOKx161BZ3q6ejWZe8b56ZL2sCuQCSGLGzHrsdw+Mi7UADrdS5+47JvSI+q2N
ohALbL8v22VFjTyeOS/b5xTI/ZMyEB6VkxP00gS6xybf18zJ/V77iOCvy4jko0/UZr0tOd8gRYF3
YaTLCigUFbkoRUf18+pieU0sZLIll3VbQk7lAwqV4XgMs7CRHBgqXSzGs6hFQg+01pTxYUE/7Z/C
zotojZrDL6b+/armrosJD7WkDK7k8sfMrF3tX0eMXXHl5m8GHrpjkdrVKe/87lpnJktIeSbhNQ8c
nc93jIy8vTGlvYk66jzPfkH43QrXkKXkGk/etn8G0WVSH0+KOfgQTqSmS9KrPMwKnw2N/J6GvxQI
nZrk9PiKV3vX8IX3vtQPqhsS+ai5FLWlH7j0OlbjjXfdv1Z8IjR5iWl/SIknTEhS8jyW1llLyEOk
rpENN9HQPREYaiZU41+B/qAbxe/jB/sWUeuSOEEtMnL4wnCHkUNG+RelWVfcEiII9XZS0xsC+vQM
zt8JKd373A0CAlQnXu6Si3Y2iTHantRDEtVKFPMXzgMDIAUohZskB+jyCA09+ppxI4YkYEsc8a9+
+liaVBOX96vPrJ0zXIjYFkM52KR00iS+10vf/PKulXgiLQoB2GxyPAOeU9T7E44x6tiA1bN3+bPo
KnMkXj9kzZMgOCUSC2vAHW+VKMVVs4pL3uZQ9hw4r3n8TA/3gBycIcjdmEHfSOz1fYuQAbCK5Pj9
SVBDwv9fxBsumjxU4Na5u7t5qHmgevktE4i8hvSLlavQwOLoI5LJMk2MG7vy9JRIshtYXKoA45HJ
pNWWRCBVtH8n7g+yS0SBPP1/GBdAagqnCRirtR9WGNgE8vYpXvtQyiAw1jw8DnRFFM/eIET1GjgU
tq1G6kesxnElE6pw2/Fp+ShVOEjmgBjzfrOBsomGz2BGwLgGNvePxYi4HE1xBILJpJjbRKTRH9vC
iC+FkFFf5+7VyB9dcqatUrtKeL9bJhvM0LTifhMNil5R5N9+l3QcZuzAAnAHUd0Oo6Z+fHkFMoJe
c8fYcXd1GKKSm4HdluSjiH20uw+Rv3LvG10zhQmQD9j6G0DIFJV8yMI3CYyfDyzE3PBsmkoD9/vK
GDqegBSLCrt9ynf8FAreVJvpYoEPYaorJ4jqYnIixtWuQ3au3pEjQri5AZWq/YHkwcMrH74Dagf/
gFXhUVZ/jJPFMvM3ws6UOxbJPVqnEkwYFzcVtDsPC23qFn4OlanR8gsVHFR80AnI1DMngJ9rPVB+
LgWf8J9NeKzBraKS9zX2St2DSk5KBvAOL1VF9GrmnL4InXxQjQxNZSIjngfVaMZnLrKxI1dO8vO/
yNZ9YByJ4k/CbTzN09oscFC4YzR4AmcGrSEs7ekO5joA4v6/EkXCbr0FYlO75kG2cZrXWbml1KU4
jFPxV1dxVgMFYQrnrZyeY1EeXotD3cMOUAlr1az86ANGhB9ez4DXTa5Ssg/x5NrKvKgEbNIlTpbZ
gtmycQd2JLiNu69FMT7btV+QurSvaHrEjsnXnLZOtcXkDUmIkQ2XOqGm8b4Ep7oRUl7TQn74fWMR
ULLEUpdBI94vVAAW0melR6uCthLVFGeEgiJV/9SQnepSIutibHjn9gvS648fzTWe1/w+fhtCGg3p
qLOvgiFWFBny/VqKz8ayaTzlObgWVbl2fEiyg1ZCaSKBw4eku1OcyUCIiqu3wvDGxgSK/c4vvYkP
qASTX2ydu36bFlS1wiUnXGAduVgYZieDjiawlBkZ7INYB/sAnkFtuQsPfEhynTiVvcjf0UUvXLOC
wdiUkkmKXjy5ih4Ar/YrhWhTWfAGTKrOP4iparKEPhULCnIDCdkYxheIw7910q9jSPl8xQeop+w6
/Q9IkaFRTDY9vEF82HayAJbowXjwc3D+ZzP5pUWn9KHD3/d+K2psdWRWNXvDtIRBFK+hN4K90TLk
y/84HxuBS2GO0pa4GUQ7YSXQzPAApHjb7HM1j+ZGnDvztIVJVku+mPbpJfblabiMTeBgoMKkO9mK
KKh6SEDNG1jNNfXjpDbGgL6fCmVo/COEi6CAlOHkQG7WArWD90c9xXQpiqbD/XfYUkeVn9/n6kCj
K6s+Zhs4XSBPIl1mGkN7l2TuQGfg5fqE3PHCtBGbHxP6w03/2Qgn3XKX7byqsj1nFUzTWHwXeDNt
uYREvQ/DdiEb5MWlHfAFJn0aVnNXH6b2QfUzTzxG4KoJ5h2GsSgLwArTShVEUBT4IuhdXpmQlzUe
emEgTobUFRMAFd0bAUlgICqqngsO4Mw4zjxvHjFW+jw3eQgNcncMrpeKrlzoJf9cDGMmCVmtOwVE
biKMBpTeMxLjLgqCminTG/ExA5hW1lsrqNGN0uH2IGZjag0oMuT9YLsScBZCZd/fx6dPeGzLz9uM
HSucyhg7IvS2kYMECc1nOzmSXP+6NNza5DWfcL7OrTqERN6G7n1a48QtBNY/OrvZCYm3RTcwPPjT
ltvsbyrk89n/v3AjZ8we/q73NIFHPkeSkr9MkbiR1Fqp7z4lfyA2vb1LwJfAtdhSqL8l4vaiuw4b
MRxqv/u8YIxyINYdfdmpjc/OTn6MeNwe9MIRAFobntJROZyd02MMDs4hB36xIecr2Z6dOCZVhyxr
FV9wqFgfIQxm+d6G6zftwyn03p3fwnPhGPx9q9avf1kpBnUIe+AgGt7iOmGaGatyVI/HzzXnpL/q
jihuHbCkcQmYwdovDYrfz/HKlCIrIDPM0oaAMSTlBMfQSdRlffUQ5qh+DQggSRLe9MEy1DVPk28m
kbOFuK0fkL64EgnUoF3/JaHitpfO5TSM7izNoUyMuzqq2HkOyP25mL399AEquXWyYLWvZWU98Xy/
9ONyPBYHIbiGS9ZTYUiTW2Zjy1jpBcZ2+U+Z0wb4Mf6c45HAZfxxtpxPy9PSjtNavkM/eNUTFC7C
7m+hxgHYWHGmRfjoURauAjFpEIBnPU8CKJ7g8SufhPmqIHTnl0EE//jCl9DbSfNd8WCJxrzhMoQF
PwHoITfBr/ysTLYTflrgZvmjL9MKCs9YrToxUtVf9bMkGrGbQxLZfTaQmClE4uw1lbtNMgZQpEMT
i31N68tp/hyUPJSTtf7qteQLduRELOv08+eluOu3yAaPuRzt3eOYAiwxiCyCSus9Jx6iJF5yQ9BV
znkm28Aa1JFroTb2rilxQyP12TIoxNmHlfKeDcHMxGfaO8m027Y+iNg+FeSry7Jz1rwiyNpK36ks
a1hiIyDzHVBFW4cSuUqwy77AYhfMrQCYHlMSA5DcdrB1fy0J8vCH+WV+CmBO3jXnU7/Q+pOevAoR
6+kKMsyExB0fFXBjtWxZIlCuTHFCVE9qZ2e70g0H15QVeqMB0C8kBOVaB//N57JPZYraporB+pNZ
jup85jQkmeenr34QfGZswLsHCTxVUoJb8EioIn7s7H1nFfzTyzIEEVSLdQkWKGw15XXbZnbG+bdq
UI6H+URq5ODIARhC1zDvLgA8rommuYB4LDKYOnRoVQSBfKbyMWENHb85e/5RozgMJiZvl1ztFT+T
KX/tn+gjDIiOllLby1kCVE3AGUZHChS76TUHHOv3OtLgfQZaj4lMtt15nDRFt+VDf3MQX+Owxmqt
huMO60sQ6fRs079AD0PtsHAnFyvHSLq+45YYi0KX02/NrzNs1B53dgXrP1iT1UyR+UQuUYwSJxLq
aIJKC9za3BKkyJQBoG8HxqIiOOBwQX2iOTov7edXHIHMzOWZ+A0okvMKZyo835eRaWzxlt4Mi5v2
uyq8ddHSAeqEA8r2C+LvGPwtSXBLS6DsSYzFV5t8V6FslZgENC1D13sSlI5YJKze93K/AzTVw/LA
35E8eYIhpDfABz3FzBV2OHMxUG4C6fx5gIKzCRwjzyfoRslLoysULIGZ1dsjm01Z7EyQfNOCtNro
MJ5FVe7IfISPyWSRI2pl8p4GTmZHXwmpKjtIpTlE6lP10DafLNx6QvJQ1GJtEFkPUzYXfowIdjOM
midCjcsjsudKkbMZNyXksZZPR61a046btLtsz/YLpGd0xrJpmYCeMakq0DIKW7yq4v3XXR+kW3Mh
kZSo3JhD+ZiuZIuuul2+QiDGnqoAu8bVx/xdt/XivdOvqrpCEHrCvf4N2NuKw93X1/Z3TeppSit/
N/mzWC16XbBz1MPr5ok/W2CHsGypAI14X6Q6VLuBh2N3rzKD/+v61pEyuJ9QobYrl/pmCMguYKrb
qzOTN/IfZyg4efKMI4Bce6xnEeL8OfXURPBVo8J4PeD59XqmGqMlYPKd3q+QW80K5JmyYm0g2+6t
gAFzlgvT69BUbKNoWBMfKKOGei3pSHDjrB5FBsH4fWbh/5/YWGLfxuqlJ2NH5iF6WgtCqLUWrhcF
2QA8k9NSdb7PDLBkEiF/LuXi/wWjqcHnMqUAaZ419oQR612dpDrbB+yHqn440LO7xSo09CS61BYy
5TIgvgWpXjMB/2Ah6/0q+/cFaD0SOViIvyVwlmVwMsTc5elvd+WwInI/tp8INNUp2yw6H49V+ZB4
PW+bz8ZimwAoxEpzAZBOx06L8gw599bp5ECVR73zkjiI/WGGBADQNHKf1Nn6/jrqCoR5eP542FvD
psi+bvRvafcfaFUxb46duPq99YiBA1nI6l0Y+M1I15WJ1X/znRnu5T9iM10MvKOIi3vRIWG6mu0j
X8BHHaJhKa1RJeVEo54i9UQEsTfFQmrQ31SYWPSdztC1rT8Bfz8N5LlNTudFn3M1usbIPmX+UPsj
WfoMZaOPp1B/wvPjpVbwevyuR3tXy89Yv06QyJdcu5UsK9JCeNcGnRTKvIqOcE4vgAMdNpY0yNCR
/OM2uVy95UYdmWNBALpmP9qRRxefWNcfitd6rRrniEfc+BiJZM17IeQAuzkYozIc9NA09t9dhaCD
ptBClSvoX31dCn/sZMY2yEnJ9tDHQBoUXhtaNyzOyXL0P6Aa9mLae7Tq5lFpB5jNnBiEN4/wHkKx
1D691v3xjRbw7D/qcuKhlPSyoc90PJlu78xzMlQINXLs3MypHMjSj0+abyou+D7FRHkH0Kn9NKoG
Ks2lA/acrnuwM5FEEoPgyWWu+i6ur0sUQ2gno/7F8GLRlAZ3jaSz+g7aSYTFOeH47pbyKUjFKYcO
s4oUo5d9U+PV0fi57ApSzP1lw8U3YxqgBcNCNMBPEBEn434kbbo957ww8c3KxWEpeZd8q+/eUa2d
nuAfKkn6K2mRtG6/bu7o3McvoS0VgdKMBF2Muj1rYBKyCT10u+tkBOMZo2vMbIYXU8alrRkY5Q6g
iHVUZ/pL7WsJ1Lnl1BRvIPznTWPry1585YA2tA/NWNz/XZSH+46OlMoB7Yu7WA1sj2BSTMTk4WkS
wAYoYN4KhDP+7kLBE3W3DENJaRvN6yMwqtPjy9+OtFQqSew23UXS4hsIQ2vPHnOy8heoQgQbobJq
g1fsNoWwTaz/7fKiZUI1AoGbf3dEFrHsVwnerR06go7+L4t6J8m5ahdxs0ybJY7nKIoXmJDhxpZL
QE3dnPrIX/ouU9GHblrii3wAM74Z6pAjED6ttf3b+20/rPFVbu4nYs56h2U4mZVN4IVjMBiZDBY/
xKshE0+lYVTPft7dy6pJIlDxh2b/JRIvLi+dtGU/wGRNxChsPYRrdMdueTfH4e9morMNRTLt0DaC
+dY/1sEpCZh04TWM+kredp5Ldx4tEXOZYfZsEfcKHJjxpj3MerhqYj2IP/FrLPnEmIkxIFhfnzxh
kzFfrx70cFsWE1ER/VQ3LHwN7KSFI+PutM/RpcyqXfl5+eNocHRPkpzhl/gnK7MU9126k9UUEjqW
c8zYCPiVLPXC8cTHwDlJ+PpvWYnX9tUNCTef3e8Xey0w4MRJ486xbVkbdHwHL6L1mR9zVZN2THPw
rjR6jD3CwfKwIpVJZ+6/GSMsPaaXmUIULb7pqribyKS14ONcxj29Bsywg6aT2Bwi7KlXc/8Y6ANG
V3JYwXrAPt6MMasmg3jlqpfxlSh2XdNLt8UCnvLxD9XjOpErWLCdciCRbEq1KwEfBAW+h+WJn0YA
y3B0YKunhuiTNKgfCFtra6wKV40QcNcNyPH7IV9AVsOaoOA7W5u772HV/m3hUOmhueMT7FrtKJXe
0NVJ94PckBJz3kXofnxrL+StNyfcLSUL4LYVmqhSmYH5EGKdnujz68VPvGH4b+++K4nnw5sXVhlj
IDiEo9hiPvG6KBwOTSMq7xNBhOPTGuapAyGk3IrlZM+Lhru9X0Fm7ou0e2xxcgIgYEurUHvuvNil
BEWNU+hu9+ub93bD/IMiouxOYO0p7uazP58xRtzDgavRVA8CBsGUCUe6IYPeJLlikJOX5hL9rK4J
9Gvzkz4YS4nVW9dKXHN41EVFq8O6zqMqltNuEyEUrRu2bCs9dyWzJ1BugxFZtsbh0wqmlzLFUoGS
48BhOIzYxklb0STHdzbXubdi+Gbc0Mycyl6KmErzm4WAbO1N3aDiWUyYNb0ee4MgaQfNX8DN/p9I
g5YmOEa8IwGlm972ctOwMh7PT/2KEYoB3iymYkMTwDomftadXV24jGbR52E50gQ3SahlKsKUU2/p
ZskahKVdX5cEUEOt+QgNZ0nXmyEJFlGACAy2SKifw3jlpzep0AsHN08cgHcAbchVa66M6NAce4ZT
vxVLPwYWGdy/nzJEF26pr6fRh++ubChhi01lfqBbnwXffZE/FfxsEyJCIq55Lj0TMry5c67EEVus
FwTo1y87vqISu5JGFv6/CiLd2a2FGKDrq//LDcrRaTXbagkdATwv3c6VAagh0ZDSSJn7UdT9fQCZ
nH127a6p2CCTzDaJbtAm5BDjy388i1WStk9XrtABfm200/nLyypZYCqhWwNYTpantJrkp5FyunH1
awmg9yZD3fbxkPHLYJsFHE7LQ2uYnUG4PYx+R2D9QUv2m011Jj2rtyUAqu/DqNRyxoqT1C40oF3x
R/CAQTG/3/G1i+LDJpS6gZWGN/nTXJYNK45ZBz3tSnXtlZ2kNA0Os7LC/cH3ibxzair8XDPcF0Ih
3fT5UzF5OCdCEm5/fVJA4seBwY8JZ2a1r+eosxeUtOR2FAYVp2sorsUYt3eASznk+zAos0eO0lso
ZKeKj3CGrG7JhnT6AeQ4toPP8Yy9ZIJcMuK6mx2AlqjBG7VQ+ULOX6/hp7YIAcLa2mjqdVjEyuVU
qC4py74AyxhpBBX7OhcZZQb52MgzvueinED0jj8mMezGkHJHh5B9oejLZBqx+W2ysIaiYPewOV71
c8tz+NQ/Cc4E5Kcp8sDyBm1IxEXjn87hO3HDvxmc3MBJmcq82ww/WFDot1Yo10Kxyopw7MsVldFp
nVVoP6twa9M5sINSgpgjJM8+ZkWRynAlv9d8hkIds+ak1jeGwhIcCKwE9iDlQwmV1gKT4JNYKFZt
LQ+BIuWQfINXL/0AQSciR+xGRoaomzl/zE8XHUdRAjGem+PhDt2/KJAGivUs541yBpnZj2mtGww2
E/EagryVnllR7y4D+tQj79Cu6tcjdaabCnlxzwHwObblfeaVlyQaeIodpZ+DDsiJdSxda9K3FrZh
tb/zfk+84r2pCUUkZlxIaQi+j2lakagIEh1tjvlrEOsemTOrQC9GlVogMzU9RnbiEsPPhglbV9Vz
VAnEswDtHHQFSWeeSN+B+ouvs0O2BKETmLju/19nwwUKkByXMh8lxPA74W7SShN+07RYDnNCR9OU
V+SKqwozBQtzWq8Vs/yOxQrx6pTLhgCXvqQh77DO2rVa/CPDbVJHuW4f093YnGq+DvnH+ebRLfpu
U+MwSesBvhAtkzurHQTR5Tj6qOPgCJ05g4RqT+XWFT23oH9qfNMelHquzsh5m1hvLPQ1C3cwOLQr
/qX8b2iFrAxmboUX8YliJlp3ghBCRLXrb3GlAPo52oZR2pE70rCVDx5DcSLJ/JoaUbvsKiocLe6I
5ostjrq59A1vYVzEdcyZ1t5dScjIXNwYvViHtUyXBO9Uul1CX68yu2Qg7BmBNnCPZAK260ZpFFTN
Mg6JryDhllDv7UxjjehP9SSP+VGlBS/wfsQDT2qbN2IdbduSUcQO+3GuvPkH+myvQvlpRNuMumEV
eIVf4AzInN15fBCyRofkeHynjepSW9mloJ48vutPIvkMSgVfI1uv+PsDTaMG7VdsCyVMqQZyjEvL
5CYJheDTeYQH8UBB71Nf4afNoztboycZswE/nGNIuM9AS+NC/MdSt4TLBFZJtkO9X9qfczlsVV3T
D4Jr5/twiNQF9ptEOZYwiXI/bV5oZkp7kc4S1finGCthDjXMLIMiGF+WQdzp0um2mWVbw0RakdJ/
HtNSQJ949wyS34hM9wKt4y4t01xa/HB3h2Duuo83qo24+0yVZd/a3yleb0do+moel3tFw6/yUowm
YybgdxPFdGoMNEpHnJDgigp+dm7B7poel8eQJhY0lLBBeZfiNFvVsO5fek48YBWzzdmqaNxWF3E4
MUW7N7abKskEzk1XH6c3WgzgeWSd0IItIgDIq5jyGon+1DA2hZLL9kRjwg2Yfv102kI8WjH+/0E8
ShZgMmqSJOUan5KNTHP5yPG/b+OznA4LfpWVyvztnnBQZgcDEaUaE7XpPAgR5g1Y3tvwj5+bP51k
jOnw4aQwHXVXutFsKSBPwCR4xl0MRhoWMlZo8DTSUyTkFuuuAjlmJxwXJODjZ7WY9U6TO6xAgex6
ojWgYzgXxI4q3ONfaqJJ/pI0fC/pPPyXzHGjksHXV7mknwmyu4NelfYw4AuUhzTs4rBMwniQM5Xv
kXmdgKNikbscUOS5ufZhEm0Oysmi64VRpVnDM3LGm2Gr89mN9ssX/iajVM1OeDa9t9F9ORugfrqy
9OUdLIh+ZY5YoFEFCKhpsBqoysR7oXzBsrLmslq273/auwJPoFicVgoys0y7RlpggNpqDDC6B0iS
ig0kvQ1lafhkqMbmtQt6cLJPVs0TRqx4PPPlGrfAPLk/24E497ZhE5guJneJiJkknOOM0VL686AH
0dni6ll0jFawfvsKvxEoFOgELDRilB0Zjp7GbmeRajiSZDAoryiw9OehrQfGg2m81sYpzW3NHNtT
bLmePuVs5PiK1jwVOIIQbowRwreBM5gVriiEt/GDGmbxbo/px+m9+O3GURW7krv/Kbhj80o68w7M
jBZsbKKUdzFsyrMyIPZQBFNLpjoC4SdHe3EMTJTUiK7GS5WhNtjTnoLO17XYKDVwkXAjT0oqyt05
WTEYOKyK9KGGlJ2T+apdo3STnzuNYmkPsoSFrGtnuHRk1rSUGpPX9WRGyz7WBrBnrDw3/FH9ooWx
/w5mT8kw5fi6sxoeCRf3MoLn5w3j9mYLhmIuhGdKmm59aYGYzb6h1VklahDze1I4wCXzh89Wy3Jf
odSVSJ7cp/wKfLkjeRJM8r4Xm6zgxz2eAuDVYwgJaAfclJF2mK5YV6Wnatg7cOdlTKXJXc4hk/gu
4avrm8e00VJQsHveys8ugaga9dZxBKYiqsS4eo30ACZ9Zz99RDD4hw+3HrCMiWs/QvY+59f6KjSN
82/o1rj6e5rrhDC0TOas/v728h3aW6RbeXyKvSzHLf+TFNVxKmYGuZKiXmGEqkuCQup+XQdaZFHn
/KuwvIexA3kcB5mhUsIPObbztDdEBXd3lIPCA2ziz6UTLFfucYbRQV0ZmIk6OrZ6s6FBxfNbX5MD
jqzTxc9u8bw+v4J0qaUB1RlaGDm7HI0Ln02NWeIAQAPJNzIhKzwfiOjTh2e3T9O6GJtG7LdigqNw
MSY5yrxLBtipPSwOoEC4FTy12MHx80LmMKk3jYdq2X4kjyDheN65loJkC+QpS4/62VLpgFbpGZLB
/yVMdl/fxhfva010U9HJtAi+NmaW9e2YUXuEM6e8lbhmUqOeCBRbd1YViOXUNgHlI/J1Xutc9ome
yTszf2t3AEvMEnGhzumBqcY7W45GslJhwyt1405wUPNsrtvUAZg/03zDmqo68hQUbmD2Cimnbw/J
kUdIRUijhZeSEQXhZnYbVS+ZftNNVR+ygjYOzA2OM2KRTzRXMsvn5MAyRCnzmDga7Ir55FH0Ul5Z
T5ALTqKix/xnJUL8edsQywqk0LsYftdBf54ezYzksGPnjIhE+G5RBqErd1MvvBz8yWXrfaqNj8NW
P4YhIbc+KYwqhDC/C2UJqA1uy5F+pUEobB7qFnorpL5L+4Vk/JFIS/HKPcREwz0siPTWLVUVGZsR
maz6kC8AbTceVZxuI6Jm4BfojjmohmL/wX42nKx33oTV/pWajW+05dS/jlLfj5mPM7NsemDpT4ce
VJ8+O/xaP09UmQqLi4HbyTny8bmyL2UER+Mo7PKlBdHIPQORkXf6eIg3hSZ/bSyYQGjG7mSLwk2V
Iq+kCQ61iKrmpwpTYPJHW9vhOwqcenbZ+5PBdTxM5Tb6e+TnlovKSYcvtU3J+Arw8Uoc8aipcf4U
+H3wV8Z+QjCz2g3Ue76mTJ0HjIGKVW4rLT+rRq92jv9kVOQ6e46tibWqjlWR7h0iMVQETQ/ACDAy
Q+C+ZH2IxN2w2UsK389s0FNw/HdBhlXM6oCHDCQhywKf6OZxU+c4nFZzgNwvI6CSKKXMQyo74lFM
pnO2Y4HptB2q9a/TYRtNb7LJUXHL7gY14auRjkFQBkIOcHbpb2nCwMQbDs8bO5tquztaL7B1YBRT
MdcbzbzFovLdlfVTSE97YGzHNRUnlw+TrFYUljYPH/7/aNWC4It4qhwd4jJM1ZHybimxKwAX3rtj
YNTPo2cQ5KMbyJ3Aw2IJxt81AG+jmDEYICLhXrRxx8JrT3+WHlBvMR1FRGhd6SoGKryzFBAQC7zk
i8kOJzJisp0vPQeI2TlwnyYvHW0iyJOVmcXfx5vqTXyapSjQUZljykli/qRkaBURWWcU9w5lHTtj
/T0tknjlCXFrn7+CIpoPAtnyk8nZqBpxNPBKuutFZlwjbUZlCVO08KihhZOalAi98KPO0K+psEuC
KRebWLmFzjZh+0EBBr5ZgdmIDaRXgT0zRV9mqX3UDHdSusA0sMxU3L61bXEbWj5pGlx7qM0HYqml
lySvPzqNAgkIPb7agIkraC92UfCvddA1jBUfeDdOaF7NFOXCXpdwQ72EHMBJ8tCneEN4O/CI6mrL
vQ62t+P1aKIu8sRB4cOiEGZ+wD4gX8cQ0RtRn8K1zYpPb+eeuTEmQurkUsuvfU2Fn4WTrCheNQMB
E/mzzsvztSQShGAOAnPCkIIX1U6a80wUjuopaxf0eFL5rCsY/MzGeb46rlQmK+wUCB4gA61pvlsG
/JnmtaSouGJWd/4N+TxZg+jpQkKmiYrsc1AQN8kGNoBv0x9Xa99HWsw0Mm+3NOU4sDUoBj+cG5PC
7FQwai2iF8QMaSZkkMOgIHCThHZ1F5/Ymq/wMWoG1e1BSehBOqZDC/j5nTUWaWupnTB1h8e59prD
6DMJlTd4NEsWVE/8YPz48K8PQ2J/ewDG3upKGl+KU/8OWWdOuG+UrjuSaZT1mn8fvoaOfehVA/dC
8w5x+nxx9ep3Tc/ypRZikC+nhgKosclosCaFuDKY1R9LPn7slsaFY5xczN4kEiaxBQBbt4LDtZTH
+ZqBfpYHlJXd/E6QL3Xuo2yOWGYc+QUjhhWimGRT51hW+ai0HCGgHDSrohdpCiwIX75fGcytFsFB
A0gVX42/0qotSUfs1RrWFzpxmvG8ePxAhD1Xx4KCOnsPsywdEa8gN9Q3xVjfQNmwLKfFYWpWY8Fn
WOJ4j22oEeg+3nx8BiSaYKB53Pm/r8VuFHS7K081f8HhzECYi5UVf9UntWlvG6sstn6vl8cX60H4
pZRGyAp1wSkEj0dU5c638UtPOtG2DcD58d/FeFhsnCtfjQK4OuodRoudC32js/r5sA0+lECCVZ9l
EBAExWHnr4C9c6iAMfb0gczFKpvAkrVayPfhTDKqEHPzlIOtsvPQQe0i8344tBlqUe+x5uDKbkGC
9GFYHojajhAOJNpdKW7hju89q8VvbgRCOJo2VeaNAvAXqqnbNQRwspDhwg/aekaNKUuPdvec8kOY
p9flK16CqrjLRVvAE84agHrxmvq2cPJ7JxTVayrc/nvcA0wjqc7hp4uu38VRpCX/xv0rG6HJX6la
Jmyxph2ESzg/3omiiW1CffGWDvFGwlUl6seVsyTXPRfFqpXZbAKKukZhgd8urPG7CEe3p05L62So
xRYDOq+5C1CBZOv924AIxFLdnc/q2ETeNj0QiftGX3lYjXBlxEj4PZc2MQHlCD9XpNg3441sT9XU
EJvdMGQQwhNkd1E9dqMKIqgX0GmilGebc2GxX7QaQiz7bmt4MAx4c/6hrkM7D4UuJCg5JCs8yJKB
7HEzWG3NnnK0ciMoGK21AMzJJoa1lvd+Xh5XNrpfLRKmVdJ6k7MTZyBsZ/W1xEW2hhkVtjSExLFX
ZXUOCEC9dSByTNXYRaknVi+SSwSuqR+3tjdB8WZYgPjJhjWYKk5KNcwjg2TKtkfg2l4mTdrZqdmo
7q6IbMYhGYt8zQbVMFtBem1PcCZrwjWzcSV0dy2Vi2DrvY+ZR3uTWdkBTjh2twgfKY4rK9Q+6eDw
rB+cJDpjh7Yj6WuGu7SLBo7sn+vRpbOrE9QFqyxaUqVZVzputRBZWeYH5vhU7TJfLXNaCAQi4Ih1
lFn9l1iock8D1+tHpwlIBVhhRa6P9wzhvZbWJGPD+sWP3gx98zIAz9hZIlYnzQLDsdlBK2n5UN9s
ELKmF3elq7y8ftPuBlLPzcW6+T22RG6f38NUo0QtT/UZzCRIRkYGVS++1FujOkVwnsAEgYwNUK1r
zFkHeLUSCxHGR6IZbZ0YMjpdxwYmn9AyYsq7jImqHN67sMM8jHUSGz+ycu1JoLpTOIlZfgbBJDmC
Jsz66eUPTlYCcLYDkxaDND9KU4Z6ngMqQo7nLQQeu684u3yl7HHliDQYHIm43UoGPlhD7bx9t4m8
b+4sG0RhizGmABKzM9oYi974ACIaJlKt7GeYeLLVMcv2/wj/oqNgjI3sgg0GC7PLWogUYM/4aXBU
toJJ6+jnWsXkOCJ8KJmxOcnuPntCG81Zwx42cv07wCzMoO3zmLLpQx3DmMxeIbHIrraTZljjBgiZ
hHZ0q2IKz0KQzZ9173UUlAt1kUKYSHbNHjVTaWYQBWtt7X0jBeUQA8aPQ6xJu6htEb2xfO4+o1dH
zGi79OhSqWxaXdyyPYdlxji97IFsSsS9G2BimHJUPBr9h72DXt+lNVbLhdaemcpxF37rwKU2Gfbw
nAA4iPTxLc5A4otWc+k4p82AJ1UAplpT8OaDqg1qEmRRqGY+nvdKKc6cvMNYsgzBZnm4pI8/Ii0Q
SImZ0D32IGnlGx3/lHP4yQlAkIUV5AqwKkbLKv2PXD6BzxmKtfRrFfUg86VUDBi4uJTlJEf0VDNE
qaiDsBRC6tEZt3v7pgxAnBqKAD44vOyrNKYQyNZu6usXWIqaKgKPfu17kyaOrLIXHe+7Fj2BH45g
zqxhv1eFBrE7fGL7BUPiaGyi0QtWAalw1AQldfLemY/OuWPz6a8MmfN+oGTH+KZKZ30lH/cEjXdj
gOKJcmXhKvtk1bedKQ/lkLp41A01isEFVhGsjNFOxY+qg1/Hefga6HeLmbpqQHpHpEWWmYxRJh1N
g9D4nDUkr5XGfFkD21alo+6bO8/i49ZP0zVVHKs+lESDp7WB5+QYEarmYaBcIM1hEvTipkE7SkXE
5FjBbFgW9ACiyMjEMSROxIs0AnIfY1APAofywSqIc8SN0DbKfph3MKOcrHEFjoklTXlw1Z2yf65L
8A3o1rUGB9wUaMQOBs1kR1WyvpOjTHnCsz4eXlHNMy+FE6B0AzC7viqMPmBAoMuY0KU9yulwIIYw
YziPkv7wQKPcdWO19o5aQWIRv+uEuWnF8l0W/2JxYWA73QBN1js2Nqxu/w4e57fPomP74cYMhK44
b+3ERxsnEFo4bstrtRVN3HlwNhegpPA0JvJLHGoMtmIJS9nGC5C2WRPjuaSKT8FZCSDBPmHLMYOu
HSdIazla97S6nD2xyNvd13T22QA3wtpQdHalSUeNiSOhY24EmjPxxQBkhPjFP4IxS+o3hpLEteEL
Sab+voOR7RUUkp3D9AbhH+QQSt6b2ONNnakCfz809FI2GlDERgBx9mtHvxT/I6YMkt7xBkcGjtmZ
NekC2u/oMjR0xD2n/LLyI5OQ8NlQNmnjo710XEvhSME3WC3mLw6V8K4i0Vxaj3a3ffgX6NAeIFCB
TJUtNBREznLYy9EkRcGkSZrDMGKdIOI0Zw/jEo1OSZmhHfPBtvkQLOXrLSuY1Ll3PDspOYSK5EwG
PwxkkCa0otgNUNeBJsiCK4klPm2n4VtP+uuF1t7+3IYOkCWPDezEF+As3DINnpMtxTUSKXgt4JML
u3uf8T6iBqlvKF04580tzvIH95QUiuVip6tMp6W4HoA/zQjtQ6kVfbCY4sVfsJuE2FNLDPZwWMiK
zQiyhcdXdqyy/RFJIBMKCQoehMyQW61wjj4VliYziUyqJwUQgcQbzCJAl61AdejHE28xZE86CtOA
gqhX63EXhn+GTeGjyO2cGPhOLlodYGVbXTVhESvjDRdJRyfdX3l9tW7fjKWgZcVuBJ/susRBwkNp
d9ZckPS/ihK2Hkqv8ZComRZM4PIQQrrTfzlxJPIv53m/TunzAUC9308INtjGt8np7vB6DN/M89w2
4gjqn8MznxS2GtCB5h6gphFuIx9MZ/3qVEgdTHP4VDjJQ7ooBwI/QZp3pS1VrKnZ1Ep37YU1czhX
LKt3d2uBI0facc+c9Zz2CPb5c9BwvveKmjyeMyezMboIVFU7bEpGAO7fM+P8KnQBlIswXIJ8cD8Q
TfFlr0/Qd8sxthgzvJLLVHVT93U9QB+cgVNVue5kZWFby0r0+hokmn95bPeVVewoxLjcbLPxXIT9
wdtc5gApuUN1GvfWUe/sSxkdV19SgY64p44raObjp2bdHEuLnHZBogUp2R20y4X+5XedApUUbg8r
Dpw7bCWx16OWiM6k+BjpbiZWhjnEyo9iNNPy1Avx/hkNVqaWpL0H/leHPG/tkEkpqo3s6bqH/OMl
dNBVEnlUKp3r69TzzWxEjR/bBhxlbA6RBfVx0GJ/xxIjAINUdOrptxBfPL9I3VKqLaDZKXys9Au9
Ih8oYJ2hRE34Oz6JhOxqCHuNZboPLXspkHu0zJqoEkjycri559bjNOKdeLyNG4uTZ0b0U0IB+RR0
dFdUhKstqiwmMRHnLYCVKZSMy7WE8ds/cAc/yuk6WwrM6GGd6lDp9JQdpC/vYlTEJBfQOCB5PPkP
cK80RGLKw/paFdQXx08AxXdKNRfvKxEfcjWU3SPnlPkF3yX+d4xaxBhoDAXtpNfuzcS8H+0QGUyZ
DPrM12YzH+b9bjUCh+lMLPvWyitlDZN0DD/nLCwLCM/g67m80RR30JjoIJjNjqSetnwYMXxsXRFO
KIPz1dw+uj8ST8ha4QQ5UMewHy6BmQGYPlcD6D/LiXnIsc1ph4Hcbh/kr28hecDuhuvzSRnvk0xz
hPnO6u8/l98tXa/lHZb/GDNzwEXwejYhzu89TdtkKE6Oaqqg1xrj9IkRHGIJstnYp93AwGTexZoP
sEWkYDKoNnnFmPi/i9Y7O2K+Q/yKIE7lIpB+ROpVrisH6zt+ss75LiQ5x9RfD2yiUNFdmzsDT7U6
lubWeCFT0ha3rp3fvjsOQKXko2E502UOBBev5HAzVK8LqhJZ/I6UQGAYqV0ftEWzIwXkk3kRbCOs
ahD+YMZmCdKgW/2834X/fAsd1bZ9Ufz+bJ7bIhXJUVc8kZMHAdeo/GIAyc/c72MIjgnbjNhDcMUA
PueyGeB1r/zbWKGR1RWQ9aIiX6C52Aub1dvu6a3ShjAecilYMeBY1AiiRja11sQuhPBQUIq5N3V8
YXOD7ffK8M0OvSXHA5i+WdOH2cnLdxQ39tetYM1PPJ2o+AUZaBZFAY6FS2kjxt62Nq+u2e0XG6uF
K8+U7+zgFTJDMlRvI4EeEBCKHLDNtRvfPT4r7lFjkcJlj3aIyF1o5Lah0DDn+LQh68KFkuzVRvEV
soPCnbRZY8dRXRKQch72RGoz+KgcAyaHffMx0Ia5E1h0qa6d8Xp9QAjY8CIgMqjir5wMv8AkP+V/
HxPjNT9WYN+GAWptDocHqMxCJNsG2Q7u45wvesPNKvUBPvdnqLw8r4G580ly9rUnsqRGXOmLF/SY
mxctj5ZlfxqYmTjS/VRl4f5pDNzLVZPP59lzvmaotvFC+0d96RNJgf06n08bfs6GKb0QJ4MvZZXG
ctmhZVeNlXC2kV+pbFRqrA+dmhkGmJfffaLhASEZlpZuS84xRz9mlkAnGTYMGWIERo3iaxE9L1kw
2JbyWtSU/oQdCVvpOkyfz37RQXaqLiEZb7LGwrCPx1JUe/4Y9bobJpt2cIhJWLXM/QGxs+MFWB16
VLtnC98wvmJOe1Er3WTjPljYQAynNaNBue+ufEWTRzneZxVrTgQrs5qu1bZKliEQsp+939JC2UXh
VgaI3jesj2WGJazwk6UCgJAoi+9Mtz+XAAI28DyTK1B4QJtt+6wVDVu+C+hvmXGSmN8GPQafVhCK
0gN4idowKNqUvgUAcq0tQXpowKTWQwi8gfYbwiNwGA92MtlS5XwgVucVKY5XAwYfe7zUCXUczLlO
OGr9woiGHpnIlLzV/x0xyuUYxfkSc8l47hPknXT2HWBk22i8l/pEnC441qa27RCGHjfW1WA57XRo
8e4MEcGOHitfMffAnUpfzfXPzyhQJcNN3h1pIUJrXbkDVEn9hVBu1wpFKufLtoJvtkx39WjnLSCM
iJ8mFYWIQG83ygOmAnMM8CUwXnO1KnOX/9RAZQCoNdWg6K9KrNZA/Fv0KgWWBc2sut+Zih/5YisV
BY12GPtKThMk5YHUTxuUsyDhwfJ6QoLC/JmA3xTeyNKkAW+o6otZuZQDviadjFsmGQwKm1KpCdgd
ReJe0mv1yxBEFaiMdoJMUsxakPYFKikMjuIwtavhCD1ZmlUnv4WnrI6USs3//OjZYEp5YiTsjaGX
YSKg5HnLQA6izKu1HfQW0L88NzC0VG5yVzdqBW9r6NSJBTuKH/tXUDgziwstaVv5QcHLDmV04r27
BsIj/WhzLouKtAh38UHkWX2MumaQ/HcA9FbtZ6w3Q8jxsX9RuEqirN9XlmTGrcENgy62QeDOKO/P
YpMjFPPEwn4wW/36y18ks7/iPsnM6m1DI9iEZPBSVSw5M7VVJ6HqMNJQrvUEA3+DVC04IOJiiwtE
OrQ8Cy+CTff0u2P2rwUPwNjD2Kb+3y+H4/9BVWE2jNJqNiGzv8lFs2bYn4W5hN2NqPGiRf5XSmw7
V1z+qSoz9ZaRl+zqyhD9TuCab6c+8F8kmGa3H8b57X0783yjCaiGeJ+2oxuT6m93fqRZAoP/6BiA
WOHdWpfYh/uBGmEx7NQ0X2C+4KuTfyjqvcqUPWy8z8Wu5se5tFPhwc1izDKmnD6w38eZFdqHvmxp
O9E+K4JIvyLJ2SSjU/pMW5UeKf5ElX1atdyivUQpWTKFE09u7356+omrRY7tysy5ouN2FxpKemnc
qqCX/ktRmka/NjatcNHs75tOCCaknvr9qUbOcG0AUdBYDmISpJtBkbUEIv6bD+WOP7SUhR67xR06
X52oBL/n586o8kRgdA+VrS6ITJItu1P4PnzgzLMikyN44qBxq6WUE41zIISPKXmnn826/yq7i1mF
TuEAzuyI3gH39pBhm063yJwGz0CUzb+4421mOMB8Ghkfa12hlqYBPCH8rOIR/IMFRts20PTJXLbQ
zFzeYTpRjb7ezWOeJAdLWtlf7SswLaNpEhL54exLpi6gpSASJ72d4GqeMUI5+rU4NFdjsKjSHLCT
Jtu3lHH3vfZivtUmQni0ZxiON5m+faZOKhbriDExF53zUfqOjrSPcpjlUirxbS88zJE0X+HLmjM7
ffeeQty7dW1kzcdwg80JsPJjrJOqy+hmA2BGLKq3cMOk8LBTHUn5wFs6EVI8apvOYUvVYVgANXsX
ftJ6FYJQIZl2aeFbGPUw+FfGf7gxlETts7IcrLdhl/yEYkRYtM9U9quQfK7VcXD7EZEFPhFMfiXH
Z5jsFNqovhtN4LsUbSsHfQ6vMk34Ht+TgVlHzwBOfrcTyvSS6AuBqVRdw5QiOa4b/y50km9z6Tc8
GKkmOrMhir1y2SO2ctZaGO47BbHmrSGyzkiwL+2HnJNT9VQkNllmZU9SwYs+W2GNQIHRa8HzNk+k
yTpP6VPyocr2shZmv33XaQNTtOC1dNkGaLW7YeHD1ozrc+OuCdSBuVHC7foprrHUliYiI+IzTKO7
/G4s/5mkgTFtLijrWLDXJFZAPvq9YE6HTw3MZT37MQqTlPKT1Hb7iAgw7By1yOkfCTMmSjUMUfXa
8q7w0DYvRRrnhWV2wnWxD2FfArwl+5wTtDR0iwD6rMK2q0Co2aj2zzSumf6OHYSNLB9mb13/30FM
o1W3E57RhsqQKz4hWGPLIEJOXG9pnG2s55VldZrHKqkxuAtbOhxQuyHSf0iElkVI3voG4sG1acbW
ESwpwjCbGf5hp+OLIyMrGL5OPInLaxNdeNbjc10nnIweV6NynbqJSS4/IQVLeXHxh5JBq11su2Fd
Se6lJoBrVlx51BiM4H4IOZHECzjxsr2yh1epXkvzdEp7v5ZfD3tmW72QxglMfPpDTer2CIr8NRl/
LJdFcwuLKtjwsske3kP3SBEPdquuVYJ5pjMge3VgmVREaziDPXMCFUInOKlWMpzIOQ0FFrwEPsMz
B87iUmUGmht44U9Yb2nKBNValtkqzU/GTrhJqdM4Bbf9R+Uk2M6A63UJNTyb8wN6Whq9McBuQXz0
RnXrRniXUJhoJTXQg+6HmP5lCdfLpK6k1UEDUGm+Bw+NwGz4eWqEfdLmIK/wKZrU5lctLXMhNKhn
eB2fFy3+UOGb44nw1R691akA7DqrTmTHsoyDryw+U239I+wnP/72EFK5QCS9zI7K4Pme//fva3Zd
2F3s1u90L3Sr7I4m4RbC/33dEQWK7f0I2FfCpRcnW6/A26qdkXfBzmNZHWANvd1/W/GcjUNXw3Qv
mK587ddNGPAqG+6zMsL1lgCM9cgRw40ssXgWDUbLrkDG0KVTEokKgYMDPkRZaAuP6zoE0KIi5W5X
iNXwPVD4CxTPKe24dGSQrRTlDBL4/xQzJzdBWkX5gllkDYJkSN0ap/j3tZ69EXh3MwI5rF0H+u8g
uxy1NFLru3pNbf6R08+0KuZIqc0ng+q4EpOstoKmyQNoF1NEIVBOPkMlRVq+6wrQAxZQfsttbRbh
Og13jRVpbN0GnPZNynVZ2kzUZoMjWiNo+A+ghUlyr1Efl0IXsMxcb+95cBH9ZCX11ejxmf4yDoBi
+K2LSPwYm+iUTpxx4+olmVtOxbgZoAdbV+YOXRctHjS1EQ9hB0I8TSZR32BDJ9NogloasdxgDa4Q
ajcJgLC3MpxQBNcIexvFAL3vJfERDcq++8A4ERkMDlWcuY1EJ7jFr/PxS+uNRBdmIgOV5Xaky24/
zER+Sc7494pUEW3Rj1X89QvlIQe3Il7OeMR5R1q8clW77rzTGOHlllKXkc7ldEP+nPCFcXvwOefV
XuWtc0m3alAB5xZVh6kaI/N2/0pQrk4e8n1S+zcy4TkK7RMcqGtsdRBLc/GZvZmZIRO9v2q/+t0K
zYfxY6qtRHaFyp1fB1UV4G1j+Penm1qGyswbiRQxlslGE53x1mwXU03ptdZfPwJwI5Zmh+h7XYCK
0mEDEsd6g1FKaTloKbLCEh3r4o9dHBXjTppmcMztzX2SDmQSB+dSLpIOOxzsY4ufeipy3ZGKDwFU
E61ppT8J4/6soyc0zeWNNLAke5ZJLHPqGMKFu4bGI6i1YgOJfaSvQ2ZXdUoY+MeB/XfMf8+x2ask
nP8R7FJqDY3OwqK25yV3w/bdckgg8TZWpERxN2DNiSE+P07ZP/t0y+ME1RO94pMPHOiJSL91bbV/
yI64Dc18IKUjFRXIXyOTMJKEaYHWGtK8mKIFOetZ4+AzGSuVo45yuOnI8v1UHDkAAjEydTj0Byc6
xBcAUzh4e5L9dY6tEpoKEmNgkCrxwpmk+bPAHZHEc9jV2LYqG96+4vyv//xX4qRVBWaQ0+fUiPZZ
cU2CYx4FMGy9tB/hyKogIcX9wR+IWt6fS/O7W/WVXyuyQea/uu+bLkhwB75VY2K+31qb9NZ1dwxT
ZakYl95V53Vh2pT4H9wxwLGbZgqXUthpdGSzCfABahjdOBOq2YAozh+xFF8YL/v9eQFswD6ZEUuj
s8GOu12f3t6fn0bUchbE137VKR2Y8uvntS+3LUbx83luRemXQnqTGGBlWfvrtwOy57cpvu2fiAHA
fhdTkvA73oDpcXqywzeiA9BO8w+jGZOCME6Zc8gYbPoOWWud5cOfv8VYd1maBY7U2l5b0V57r+EF
lEwXMlBpGkEC9nar3X+kMX2AFeQGOF292y1eTgleOA9HM0NMdcKWRAfUHCsWqI2AvoYnX+Z/hpgs
Xq8okM3LovVY+gooXyJdYjf2DrFlKfdIspi5FmLN1mVnM5aSdMdVcxN5csBSkHKnElPnuuGWDscb
tzOTqDN/3sR7lbJoTyvaekygovd4Dk9SwFaOow9GAvi5tRwVKkYXLUMSq1kGqTJcwva0n3Vi7Rr4
LBvw0iTOgRp0m8OcQt6M8hVNK1wRzhD+CAXipTCwFwtZpMa9AKPoUCykMcRiJaD8rGinK+Df+WUI
G3nCM4gPT3xrPOf45+ttGbjdI+ubXZwDhhEibUE5WwMOmORkhtm5mCftKJ/FkgqFwpVA4kHmi+82
YpTAi9YWKC6JR/xjfmzU/6Nr3YvswzQNa6WAeFAk4DaKpsICOtSMIntzz4qoeVmTr7mLzgMBBpcZ
H4CXra9E3PNk8tFz7oPxD6aZnEfREhSs1meCc65wUeRiRbLFnIJ1Y2bt4IK6bN3me/1lj89Mz+XN
0DrgJN57jaGrV1K4OF/46yjBd3yd9d9XrZJbJYNVJtv1SY1fMWXsmQYjS+qEMzaPL0DmKMwpX52P
9n50313SoxPfcTtsdFcdwj/5xUXAq8TPjLkqIfOt7AGX9k7Bo3l5sButaXS4+5MIi8+tZnggS4b0
mh5d67wfoDXxBw0EG5iecULBGn11olEup1gqQ7/vTyP8iO9FMDOVsSTeaU4ZNo57sd984oPbM8OT
Qh02P79EJ6/J685J3OuW3UraaV7NG72tapqQxXU9Qblh1Uums59vr50IjKB4djHPPQZZYOQ5byHL
MKjcynkYoGOLPPIRJOems/z4+l6U8vv2v7xjrQIGBStST8s87OlqLc3AsnMLC0Frqfhmj6qW4zDM
owtSjilaN0Z2NYRMzMSSdvywF4EkQHwDIcDU6tgYDpTEuuqoPFTDPtltMKpk6hDvVgKcsxg9G1hg
QLjCBoxyGkDhrQ2N2Hl+agcnfxvWoseLtRYVG3JGJ43uZ5utWr2R6r6a4oaXyPSlBeHTZDYGfxXa
reTotNAEiurabM5tInRSVFWpi80dDHFjJKsdT9Sq758WH1a7rbBpWbGYvVTIHXB2JqolpI6LVB3Y
O9lgpeAWmXrE5ZBUnf2o1euKvNSrAgEmJuG+sdyei3z0IzPsBWjKYIQ75XTa0Jr6bQuIV2P+96jV
Mwe/ZN+GVr0E+WqYB7eg9A4ritNBCLQb0mcpVUm8plelFl2783RQslW7xsdPv5GITeJJOk6zr9KS
/lIHIIpSVyjHh7BWtddgPkAreZVojxDbZ0A3J+VditNdxafRL0C6ZXQYRUbZo9iogohskRJ8BF7y
/4oc2MRiMoRxNFvWTwovZya/r4dOkIcw7cTPb7/GemU6f2X9Jualv18KSmi7KwxicqpnGcDlCTvF
dt/RcxUBrNwHH35r3tq/8pigYHJXOd+FOgUZ/gybngKSyTNd8DYcQj8MlSuy9zH9f9RALYRJ4zbP
qguv0sYJX+uZnhDFDTlOzy4tEffvNlsV9eJqgCcpdiROM5JvlZKYdUlFe4fDPo0WyVfg8lzzeHsJ
hJ1DaEalwLiNHo5v8+80oi5jujUr1Y4KMM3SzkzrbGUhyGaJDr6+dn1GFNSlfj+ErK9SohHbVTd2
uSYN/jY+IIYmyFG2N8EOzUMi2Il+x7ZNh7ysD80GOpwun/5wsXj/wQSg4ziezgrLrCixLs5s98jy
oz1Dfizcm6D7Pr2oJl+dlay4vmPm2+6ENOZEuWBLM6VCiIYmlXi/N7EcXZEfkN1oQYxj3Ro8bM5e
7HofdyvdIdQbaqhCV0YR21MdCuy/aOfZakkvUGi16SbesbXifl+4giUJLTD35IBwFDKv6rpvOlp3
weJLR1jbVj1FQBypuPv9/Zy9EDK9fttVOuFp3LdEbQwXtyVNTjN4k3EzgseeNcGK+RpJJqfXkDO0
lBcD3hijbYzOltJFebMqXvtAUVE6p1Q/Psh0jj447C8wu/M4W3thBHNSx7aAjXgGdRIB4TsNgpRn
PxF9McvtaSWv88s5avzEGpv2v8hXIbIFlJ+f+ySqDruy6+CLGGGkatFBNBOxN19/XfU/E4RRPra5
dj8Pjme0tDylLyh0f4d0MNLz5pZgiElS9zoaHBUW6Y98jVihGMGFd9/zsxsqdT4S4b051+/hvepa
jaj9US6Sv4EsL7bZqEcGFpBKZi9FPuBvKtJzhnsbW/MvjhrDP9Kh7hQuhKcIYvh/NDewUCAjY54t
gIj6f4SRVwYvjszd5sFiD4qI4uP5AAKdeWqRVrWipnDB6q4nLV5V77ApFLGrwfhmI2yyKKstbWfv
7e8UR7wiC2gP/LDnWW+LcEkINhAqD7B/J7F18JO6pVscBgvCStiIxYnLkFzS/fJFQ490RLHguEeE
scxVOAPQ2Kb8rmZEq7glFZ4PZ915S/b3onC3iczjMI/t6PJvZCBA4ZLNNpoWlnbvZtxylW9yA7gF
7t9o4Oc8fL3Wpix8I9HsdK0xq058E7jxHVJRHr2WXK3jd+uxxYAXDMBAVOcPWoHxKDDc8kOosXKO
BAQxtZWwCCIgJRgIk42+fjYRsfF8nitS9VaZdF328rxS8Hqg1ykKF1Vhl7NKnYQk/ucsvto1QWCv
dtTrRMy93qzfAqXZJuuqPfMAzQuV2DELMowY2Q4zw4lpX+GEyWfFG8nQe+J0PhgOr5eDCJiPv5rs
lS7GS00xzSvGhYlSdM1Iwua9DEocnjQQyFR6Rp2Ljls9CZU4yqHCfxcTlOLxf5iLZKqbKoso7025
7yJyDnrxANkxu45qvkJC2Vi5twc1NDJ5y6tVly8WHJsgUxod1iDBn52q5iXWFytaCfZbpFfaa95O
jy8b1eOhJx5n+JYuhJf8lsMijM7jSHVYNNBG9xRMhhRUKVwfE+5HplXDfiHeGhcPyMyvfULbbfQz
i0JChlN5+hQMGHxkUo9tOl8mkkP22IsM5cEXc5mTcwmtK9QCy8jtHDn43tLZ+zhWtkRrJflA6HyV
TGT533M6o82mBt/+e2CdloksaIH4CciWA3Tn681ZoHkjwzIHGHbpylxiwwDNdQlHEQoLu3tqGQyu
kx0I4r2N260zUvSOia3rKduh287/8KpJqZ6DOosqgSXPrNzrszGyCqdd+svLYD/1ptcUOHEMFamT
lDcEK2Nn8tM3ExmigP81mSmrjWmtfilvK4Ey7u+lUFHLmnylu+/bzUZtwHt9xanFO0DJo5dOrkKo
SA6AN3UhAkYpnKPcawwBqTa/w2AppIB7vgwmLgcRbGsTjSpUOiR3FcssbZIMUfLMC19eN9c6r9BX
PPBX5r7gonq2j33LaIwE/Eg1gTA5FWHvp7Auc3tL0zvVCWm9UfbVFD6M5gvKHVLFpaHy8VRdeBXZ
PiVk/zmu+87uPqLtj590vEr5ub1yFhvNxcerhfe7G2Lhd0LjFA9i7hCsypSMiH9NCAM29Phqpxh8
hrvWAOcDA1FeuP3S5K4eMH1YRn8dDnOYQx8e4BeGNtt+vIx8e+M3nk1n3q3plLEdOYxLgIRGndHl
rFgxx9YpYGZO+KsC8VdpAhH/cTnPVBP1AnrGrOxxZrLI6sIB1eS/kuAZriXqpqGgUC4Uy3+TwINX
kmeLMGk0Lp/tLryLYEbBn/nsj1NLhRyDR1HSZHydBSJix8qfV+uK72/vtbZAWWvABwV1HGNFQm0a
24ZUrjLYTPBlxwI+/IEAJpwjg8WG43PKwJ5gDmVpnmChotDjB6HKklpgCKphOOrHzLXLR95NNtuA
masYw4e+XxP977eK9gPYAjS/r8vElwB7x0r4eIa+jZ8swJP5tIdEvx8GCIiZACnyNLH9/WDV0IN2
0Yp2oSSkj5nAF8gfaQK/kB7+GdVvQaDQkuGwULP9fX1mmDPcs5hLhXjQmVb4uv6N3EnYYd2N5dGL
07BD6jgQVHo/IwfvAiEPKMZGvshl+LZbQyxk42fRKXeuf316JZlBf3N4DfUumEY9Kv/smE6dKWtj
AYRXIIGtbbMV756yECuVGWFczhvXylmEUU1mSZS37VQmlRYep4/5/ivJmPRGpxLysIK+oXKbs0q2
m0zyZ/QHI+jm1RAyrhycW27ZSkhI3YFFy3Ngzcv6FKaXR1RhsmUow9IYvYATKuPiFRjQWN5cKP0v
VbuJB39hZfctJvLFf8CuAjGBpN1J5aaTMBDLSP+pB5l6mtPb5nn16NiKXtGqWzLFKdkjOoAmikfl
KsyWaWPk5kSSFBoHOqrZISHkN31cziUx8Gc1StFZDtNz4MeNgCgK8cbmRi+nGzbOFfc4XRJ/5O8y
ppymGWnXcb9fTThHdDi2ReVZgHNDxxazrgcBFgJ05PN/iqOKHAcdCT9VKFKQycUMlJaY0uuqQUpH
7mfTShh/JsTVJt/yctdZ2Aj+pu3r4YTVbJtHrPjKzaz81tlxmRRwdsU5VfogyM83z/0NKFDIFyHL
W7wk86MjfsNwiLdHzy7ZT7Ahk1es+Nl/Rvm6rkxN5jrpMd+xP67zlh2hfFYtkqaZCqhJZsOCpLZQ
gh5B9EKdWjMUYbDhJK5ZArcWSI+zqo49EKkcDA/QXWeUIzz/Ap2oAdrjTaVAU3j18kKHIEvjP1VE
Fp8fL/XKkXqKKF6bs6ZJvgubyX85Ot+Shjk4hzvqDxrK1oTiCLQaxcpOZmDZSDtSC6VBT9qBQN7y
83/AdVceezMvbwIJ3G/3ceZy1yppdbzbBZDOIMxLvalq0OId7eDtz8/taGrzuYX+whn2RAgitkj2
v8Cf8sR2uXscC3mj2QUuvvHemjtfJx3dgrKYPAoUG3das08Vr40npvsCx4vx5gYsYmrJuLVBrANu
DihcOVbiju82v9rMrTd65/DGcgmJ5LsXcdybCggPdnJbi7ig0JNDJwgCrnUf4KwSaQ74j1N3O1bU
krGtN51WKNWVk4PdSwWtFTGCu1ik0KnLcjrSwEhJ++2qawWNX4btqDi2ON3R8N8RzTqzgnUzBYuY
hyTNS62AueLQptW/KRidwDRcauDG6JuRyCLtxYkQU5TRjlFOU0R5DjtqO8vqJJJdDIP4cFWGnnSc
vN3KPt3u5av9IiRV1He1q0FNKAkEllDOpHenMYsbzz4O0UYfJSct7bzopJc3TAF2kx1J+IwzJvIo
MYHql3EJVeLfHfmS9ha4V2J1OpglNbXXt9ySjnQ81rWTPvLbXm1R1prmiGBVeRWmiWw8hrm1/9jr
41+x3jaTmYrS/e4Hgbqrr2YXFRDnF6ZoSG9lKQhHomcI3BmX1AyIxN4p9j/d4R4MnE7I2Tr6pnTX
Jd0KjUf6Ga2PGhtK7zL8JNMY91pkWa1RIjzyA3upU1Dr9CG1NpXTD5iBR/oXPW96J3PmqmJH8N8Q
CmzBNUX5KjKUecAiMQijhZjNVxUAGSgrg+R3c4rQjiZqtClS4+kWLI3J5l2D81WtgvK4Km4L0puQ
L1hblsbGqoneUrjcBgfDw5rhbVXEjsP6DX7cFC9WILNt0jnyDBblTQUJB2ZRADlh4rGEz619925O
nCxGCda1KrGNVq2LMgq+iWKjxJ1CfUxv/KLCYQ2cHDqXTT5eOgLTXaw8c6IwwrMJq8cstBp7vnS0
ggkSIrukPgXu4vocHILBQytteMcgS5DiVHlCT7jsfTHNSre9F3NO8qnh6ISuSgcTGTrJ5/ibNw7u
VXWoGTcX/5P0wDZj4Uih3Npvbk4QPwDmvzjiEGY5W0Hm5aTfERLo46UA1ZbQBUyMdTaOjCBYMigW
n8KSYtCWxpipnLxtb1t76zxoCXPp2eUwthmcyh0XDfXSuWCYqDRDXGYYghuN2n8IG/ZfGNS8zOj/
iEDGXGdkPf/SWJELYnoNmzqJQ2nLF6uMQG8GPeQalysZlN/imEx8N5jQPGyPWmSnMKbTYWCGAmfa
I+0g1q2BBeGUmbQEAfKbkjoNnlJsOsyJQ7d1wzaXEMjNbxVhK70lyEnrDUzYP2xFBx7mcNEh8qzX
QWKStAShcLXEefk0qcgOeb9vtwPJ2NJtHuyrUO4DEMZYbb53S5zhMRnLac+XhkECzTltM41y/ANP
9r35a6B5iAwImRuKs8+Hx5mjcpZshGc/JwafxYTgMdzpCcCm2r9+2QL2ET/dP+g33QjmZdvJQbQM
tPRqB//o6m2f4ZjDUahF19nju8o1HHPBgKTuSOHLCQ/ACkQPgVQZ8mplfPzU/ti/X0dHcmbEzTih
aezRXOJtU9YgGD37w+F2b0C7ztcQGnJoidjmyXVdwDXvTOOJpUv0qRGJ+0cSQGyUpzVznrhymSMs
DlqIZ4mWXmFNP9DhosfZhbq/lscz+QQAwZhQBuNnS7I1xuI1vWyC99k1Hd2wdAFwofCuGnEKnxGa
ahkBb7GettCJOpU5lfE9DML3DSRzpJP3F04KPAKAaTfNhDwiRp8+thRvjWv6UMVQDWmn7whL7Y9d
mGxeyyPKccLNEijG3Q2S+HR+LKWv4LFTGfaSm/ipARDbJS3Mce1dVhA329+zBFu4RvfimITtHc/o
Mf8yd3MzUaTK/2GhanxWmamMkgHewaEtowGSVQsuVzHyLY+mJkVDFRmUbXaHDh4r/1s3t9WgbzDM
ie/7QbblL+vSgaE6wGztEibwDgzQUiaJY0uGOEbbhg+LSEIK+utFu9XJI9FVbQsqcX+KrdKH1SO7
LTmjucXE+O/txGWmbrZoA/u360nYF7r1DlXqhNjgcij+TxmLL0RbpEXEqW54s6ynnIDZqBJfkHqd
dqA2tWp7o/0AfPKT0lZai13GKC7VfH8KWj+VUJXYc5RQfU96XaIBkz4tnZFTbVl+8QbVWaheRfFY
eyhhAZV7BeC9NMKAAIMJtL3sbdJeEyvImI/KQTXbbCpcROBWXYpyNuZAflwpPGAemAwEgbHq4XVs
2oBBhOndY7O6petKL5og57LWS/3wqB0fSHlaZWmewNF6hTfb+vkX7FV4+rd6pgV+0TGAfWWjlBXc
q42qJVX/eqc2KyYAvkxCw9wrA9gVs4iO34pBUCQS03nwWC5GE6/S04M6uXmHV2gXfrT6ezEqa0kI
j6JxQVjD5eM0GrQFdKRepGuIq4CIlFPYq3KYQatDcPp6bybbPsN09hUU1WvoZOZTEqGhsOWR3gn7
A1WMyPJDoe/jewfMQGbq1bvz0msZcY7B6gWLNd2yhJoL1bWvKM6SvY2caKterc8SBd3SkK7EkhT+
AVtccyno7hc7Rz/XtcbQX89rFxG7E4SO0UtL7mwZrncKqxVr2MyIQCBE3izpkMQrFmikrjFBOA+t
MSCwNBhoWWjxEF+JBt7KsUlvSVwy63QE7xEeU0dI8qaZVurONY5CHjJYpHkbeeL0JRl7qaAAe/fd
ypCz8jyUOuZKk7CnLBPmN6lOMXTgF8xcajQPw/T4BK9kKJ4RmG0dzN2t8DHz+41creeVjlcdqpVl
Wv7TYG12rTbmCmLKDf+UyJliHiF1mMXquilrtnKOY+XM0XWOQpMZ5X4Ii7wWaNLK+K5sFcwYJAYc
hEEc3OmVMC1z1DPHM0FSkjHD/cEJOSm4gmPI4oGHrGc97AzAfBHzhL0mEom7d1mEXEaKWFTXl7Ry
rhlpbagdwbDXpaL4OKmuI73nVAhlJ/ta+kR7Wv7a820Kgfq0sVBm2z8xd7KgaPVLo3bke1r/eJSV
l87GbV4G1jKr4p/gQJRNXQ89tljXCTlhh/uFZFmaa2aLCg+/lyFC17kkmaV0TSqQNpZUYY0FBd29
5lL01N/xkUJ+/FYM9EaPZ5+noECQKUQeGVVRKMLFzbswvnKkSEcjkgINS3hCGDYWlwV+zMvvexfr
cplVmHVwgP5ITQ0wZAVeAjpOVY/62Ak5FYfSkRm5Fl/OuA+z00yU4rlZbVVTvU2iVxpFDqYVlTcL
av6Aro+HHUC2Nhk78MAhxMnLBmaoztExiThl+/m3Q43LafO4NCGfkgjGpMS6TsQ3q2TctQD+kSCP
MaooX/DIg+EjlZgg0TE2YQdqYM7DqQvVBKticRtIMxaCuIf4hhFjEhPmaYMKgix036zVy3jL5/jD
EYgOTH7bx6GjLsKmds/eSBgfypc/m7FHsfKl5ILUuDGCamc+hI/oc/onzQN+quV38uM2FBBUkR3l
Cfzckdcxjz4zOh9PEQ81LyfWt07VBr6XDRL9GvGj1xGAOYgZ7QbjMaXGjgfOFjvhiUps/Q+7WkBh
BrlYM5LnUN05SJOP3ihKo7S70mlxPDXbahGwtMDC6oFJquuxLPJMp4ybzQgrcoQEbiayMWdhaVKe
L1s3+N8+NB9gxlSqvFcVUKtfLp3qT1hPfqNrtaKExjWkT0FdOKeM3zHoc3uLs9rcMKjWtogSBkup
8NWYhUba5EkIsSRCBFZAM/z9dyUfGRWGumeH1jOqjho1cd34QCRYJMS05RoMmTj632SW3f3do/Sz
6nEpJJy4RY3c0ZkSbRrZpCEkrjWJaurP981lXDRcgJTpXcAgjmMeruCsh98e9Q4qguVvOU/ZUAKk
l91soXG+dcvzvWYGG6hGcESQGMD0L8lAfrEQrLrDyGxrQw22GMdgYNpDjh1MyRkVORqNVf102DRL
UJv3kk2jbb+SUvHDKVReUDb8LFDY148lQ4f+jY249ycymplXF3V6EbsSXPRkRspV2KV+zzt+tuDS
t1Rwyz4ty8ZayWEKHHlvvERhgfQxiFquzzLuaowbk/J5R6iHDd7lMXKvY8a31XnP9sM7Lw3Q+9CC
IRjgFbqCFPYGOwg5ioHX2/B5aXlfohWVCZpJpMLpp6PP+HRYpQ62u5YibstOVn+GvKxtcAdCPr4I
BavfoucMJRwliwdzJHbh73kP6+oscVAfgkNqWcuG75iZKGTiCD25pSXUTAdoOZhlORlGNQgmbUhj
YbzrQVC75eO1tDwilmjFcn02mXXESQzFyZ2R3y1IjIMZyE22sma+zo2V0fg2n2tqOkITyfM2fyNc
oQZsXM1NbiwPeZmu4u8SZ8y3ZndV88ts6KoEKbchcujlgsJwxWgRK+T2x1VaoL2mBLKzlteW8DoZ
w5MREuoZKMlTOreITP0Mrh4bpuF2BOprYaFZAXqcXTACF2SipVfaW6OxE6idBGW7vWv5I8peAeqB
6KzSYgNKsUhH80FIWK3GnWojzqzsVnbngbEKf4y+h0UAecfsUkjyj9EX9D6nywf5ld/GQzci6ne1
K/jwMY7baCUGqgaKWXMsrVfaOet3s1ZTztt+XLz2Z1KlX7Zd5LYoHkjojEXnC7rDXYwrGOmSKTS0
d5B0dE/FUdFyNTIt6RahpAcWdTx68LVZupSXp53uslnKzotGLnji5Iz+2z0SVQPMg6VlF+apXimG
76dxf+CCY4MKgYHKLwY7VUSjrzBuSb1M8w9NO/a61FAReHrni+RY6DIWtPzsy6ATXiWsKGlFzyEu
w5UPuhKW3jfW/3EHMzymBdoixxttqPg+cbx35ADQB7NtI9hXMXqn9pn45AMFBARu57JJqPq1OZ6Y
kbcgyQ+NBChI+hDo9eR1mzIh4ZbaraoFRAoPGEwI8+g8xr4ZGzhF2y/Xoe/W0eaAsJ+DQHec5vqi
6oJmFOmU6+HwIFKwMCQT6NGIjRTB6VCZIfIJQ7m9HECRjP7NdOFcQ/SE4nT4a6CP5tcV9rZbYZaA
PEpK3C/ptub1ZZHA4SGLtu7MbNjEry+PN1r0YXYGU1zWw8kfSsXJHvHZlOJUZCK/w10+pOil4fQg
wBh8jJEwNyEXl/i57JZ0G/z/Sohc7iUI5q5VDETlnqYPxSFu/wJJABnc2iGEHCxe8L3vqxlrZ/KR
iUyNFVJha13hPOKtE4C5CHxUX6RRnlSaBfADrSgKY2VNhoaBScR/Tm1Ic+iqp/0g3wM0YeVk5zEM
H3ieS+mwDsCIGy+76rgM3K83I/cdwAzYSepDjyVn7Rbt+qSdSCeCv2V9d9KYm1JaJdykJ5bW4qQo
n2o2M+aDPgZNzbFrj/KGAvYd8WwSef3DWNChZqqBvp/vLRKJAB24NwQOOriaSG50zSPxYKpaL2dB
1+9DNWopLIHM/d8ZAkRCUXpfqou7SXc6Sj83VhL/0zyEEiyow0FvwGuLxn+qrsWlW9nGDQo6sC/Y
Cuxb+yWUaTAHVXu+dmHYvE7L/Ja65S5dxfn/Tct8ey2LL96hGIuaA8aoYlkoi4xXfr4KKjBt2eFV
YXqpwwo2tj6EYEVCEBWxO+W8fS8BMfOgdDk0M1LaMZ86LmhMZiIKb7MhNReaR2pdoS9mYwcjQwgy
2nZmH9L0itF3DCI6oc0V8xHj1V6cgLTK/1cGpXSBCOX7+AQ9VNSQPpO7PUio81lrVm1UTeP1WEVQ
b0yuwv3zChSk9Jdws5GO8B4K4JaowW1wWRU6cAvw9fGP8THkwSzqeyt6bLHmiCoCUrCdcbEqBh3b
0RYzjV2ZyiuZl81OC5zzl98Ql8beMAh1lfM/LgcvophavEeT9f9C6LbOASaM8gU9cQiMJzwYnkX9
4WxKaaKR3XRm8kijYfm6qqdz1l8g8er7RDYAYAlPle5hlBS0NYO7xcFPPXMpqagoFOW49IUx0SL0
9Z41IYR1nIOyVWKg3VHcCJsK7eLXASHk9+AtXekS5a23dhg8HWV7wL3IQ2yk3srXPSIgDDpaGWAH
6T/BPCQvrRXX7Q+nG+JUVEGTpUAIujHfyr3KP7bpm5ZhqAs7Uwa+FK3WcG/3f5mtM1p4PmsR9Lvv
deQemYAOuMGx53VoFJOKxu5pFs/AK4ouItQLPkm8ru0IgcLiI4zEaaz62llGR3BdTYF5BVWeD9AM
9+J+3K6NBIVxfIffGB4R/Zd2tdZ3wzzxKzGOXbxhmLXIQJ3yyrid/hsagLOcgWbUDJPqXEfCKrRZ
kBThRtMq0tXlNu+u/A2n94jqMoX+KEKi9A3WErEOOA4nhJPp4KV6srXxtGNN6Q/a3ofANW2dtQG+
SsdQFPWapFeRakojd9oUikawp+swdBbOiWvPXkxyLMzzgRAVe2Wl31vAiEWDfzIsJoMqR8IOKKvx
KV8k5JBxPIUrpuSDvMAkspiseNfUJkwbAODJSVUJDQkIJ04BerJ/dVxpzwlbQ7a8dkLBaWw0Fpbx
zH5gYOUGcHoJRehl+kuLeGxz7rS3L2cnYd75SymkW/JVeDG+LPy3JzisS1KIUfqMEkmp5Tj6R+2T
PTMAw2ZKMeCS93xKjyYz1NXvpH6CpgEtNGabFd54Xr/M/nG0P2fepXAD00M87IRSNPvxqcp0/cLp
yYcE59tn5pyqx7ad8sy8ennxlaw0HHxB2wiRWt4Ggh0Zkb6N1iI6xwm7QN6v2uhT5hi5K+ywRBQ+
Y9WSWnNBfGDNCZu7yS+miw9abuA1I9n4uFLt+BYs3xnylXjeKNKZsDq+/l4CnCND038Uga9KTiB3
ZuIsTLii1iqt94c54uccuLfb+iDidzcCI3AWccpJ91SdoDj+XxJ/WP5ApBWA6TcNUS+8EuaXe/VA
GZofGUMwcuEleyn1KxU+AavC/WNUi57xTM/uqyvFi61vduNsN4V9Tk2in4v0C0C3agV+bQcdnBHU
S2hEC8VBGOeTTMSI7chi44r/mMm+MkUonElMG2PLgy/2P2IDOkehAhq0pSD9XwQ110xlO1E7WP8O
dDqAoEc/R+DtIlUv/hpgCQ13W149H8c24XFAijNAz73bVaxqCXwQOPwB1X+wFQby9v7sKdaIY5P4
x4eY9jaaK4hoqUx6phSBbr4RoFi8q54rBV1PRifRzCA2K1cTVhn7VAdG5xYqXawCrsDr1GEGo5eq
rtFmHVZ9dlQGoc2QYByFRLhZwV86u7xYnAYTyUsdBuFKblVreWGEloGenXDkhcagsGhm/KsVh6gz
eiWgdjIkQGm0AZySChIjDb3KyX3rhnHrkzOSJKkK/cL7XynEMACNpUywBpllDXsC1iGSav2IivG5
8yIdBSGuzvCf4BR1P5dim02jDmI6k3LIFcNGI0DPLvzODoQOK/vYdMPQxS4gNDt6Uztl1Hqah7aV
kIbojNDvaUO8AdQOExo40sJaJEyy7BiwfNqlurpqIgdyMvgydrifYfiDRLakhI+rp9+XoPXcxTEF
r7ErpuWYcOG1a5T+Y4wESgk4j+a4BAIGapg69xj7GdC8Ge3kaRfBfcvwoMGK8IikrHesfiicgxUL
hFgfwCNhPBn+64n0HXk/mGNZxfJ7JpUrXj4KWdeRdPDC4q9Ay+sWi6xFBVWrttRJ3EjE4cVGcmqR
lPrO9VaALjOc6IHBkz+bHglOjNueLVDzYlHEydGYsCIafN6EuoK18oA9ouoS7r/LXGXc8fMI0KrK
/CqmgNJK41Vaxk/ojAunFbGEcj8DeJ2pWKFP3vyHaD2f3A6hBt4B3tkmOV3T0S4lOruG/Oy5HFxe
laCbYoXtSi4RbBln3QfQZDF1iWhQrclWHgjgPAZo933MjcE1yJ9lbOG1O7jG5o+ctoFy62KLaJ8k
0BFCUVIUktbfOELj6kOHljoOfike04/gaMNyrIMRl+aacmtr4oeJOwxDdcjDIkwcY0mojqqxJhHO
oCA7E+5lsVyW4hLByJhR8YmpkqVuFTsQuDJ/rwnEpIq2mRUC3P7jWUVj957qafG0kHH3oh8QA6BQ
3Ap8t28qimPBXdgLVYi5e0LT3DbPX86zVIUiYQs2mMIgRNc5Oti230eP+Wy/50/q+We2WSq7KtL0
olBVnB11PgOn0ONm3dVnvhUqPQHJlcXsAz3IwnoMOe07uFH9iP72tsEyuEITznjHVvHgUM2bBxXm
xrMUb88MBTYSou2PZHZrZ6VuKIlhtJpHPtjc8SZypmVazMziLGJhR9GhDjrh+BQ5F7OTqzV3hD/Q
ghal6CKPYv3vqu9BDYDuSgQtqNxMDTsTU7oLxhnV7O28RSfYAL0OfZ9+Xt8V/ZwT8oMqasPZxhvj
kPSDb5aUqw1db7VAozJWUGuZoH3XjWHfe6yW2gKcVv61yOqG4JtvPRwQTQDBCXzVBNChgQHOORMx
q6zXQ7dgW2AJtqmanxn3ROCDB0K3pogvHWhAAYel2ZJwY8zX/kJt2y2fHg0WnWGSXswE/v2qDPdH
2dfat2rYDwn92CuSV/vsw3w88qTxPNNueMIxOY6ynJqBuazN/xgUVBWnHufRo4pAUUFKsYU9qIrZ
FW14q2j5P9mVEJxott/RDyG+BkBy/LvvsBl9hLNWOngzXQ6CsoHlHZa01HAK5Kb5Kuw1nobmLRPB
hy5aBVn32WHeasIobI0sbwgxcZ5u14DQL6EFKQQSu3HM1mMaMopIbxdwrL2aIDRSIP0SmGzElRie
TV6s7OVnBrKTvcQRaLSV8+lKaMMfQOjLrKecQfpHzqGayYQdAoXMxhC0I55i28/YxeGjSFJZKrHB
+2uTYFlYHzS5mysDlQH9xrJNWQsVDOV0CUQKNJeYo03FTM3iqITQ3lYsCbO54Lm2KIWGRrKZzOVz
bBSlVO3vT17/BnxKI69gBT8VVpVZFrNaA9+chxv0Ty6n4VYGv+D6GW2k3rvCa0fPvwczxXWob6Cm
mijTkBELjuERrGxD39AuNSS7i0CR8GjgckzIGViRKTemg4dUwaaiI1Ptgz5mNLzI/9rzrarCpLWv
E9YmR360iZLzAvcH9UFcVhJRM9i1P+yXHR/clfVSYlHyKNOhBeGD0BLqRsEAVGgjx4Lffic8ZzST
UItnh6wjKVfMXt0b0QwZdqzR8HxDFd2fqytz/rbYL6tDX8pdoN9GlIWtkkrEz//wynIj3YqawOpm
c+eDGXfyE9rKEPLa1VHqaMS3zx0DQksEoul66bUJjoJvOVSbxCbsLquu4708hOX1HgN1SRjKiPe7
2fiy1ybUZ5kA43YOEO4aYQ2rPjGCi40pwLHKnYtxMqHKsrXyBLvrymh40RScP3NUByAK/xrxBHHC
0VRvaz/9bSRmFlai2KBIsGkrO0O/V+/RDvPrKyzT9N8O+KUvq7XjQbcOMXfQeWZdHi4/KxbHopXd
wqMSpt8lOnETrLrfj3IAYYsGyn8KdOwJ0/Rx+7zAeNRoXtO9a7/8mCGhrlPwkM0PaD0xgZxwRtUi
OlOs4skZxC5Ggp8y3I57nTYi1STbmsTIfJZhkY+L2+AGxSlA+yumFBSaSJBywWUJmjNc6sRHUFkV
ASANoEyKtFZi0TtC/YBK0i1ibSAoaH9xmcEgixlftpS7RMWquFiuTa4ecR/5ZC9mEKxU3TSXQ/ck
4cZe4S7TW5Z+1Ym7mtwjLXVyaKdP9W2k1P7HJcMItVW+y/kwbwMYrUyK+ereZbtp+uKu1XFwIQ3X
r1oiHuhjD/63RooyJSiLfSk27tD9HYDYI+NTsPEQuLZ52ZPOctlVuOl8w2hyKet7IPLWHJI4zA/N
BsLTmcwbLNbz6WZwHV6t+a/ugdTorJafDdYSmYTIz/NPNL9Rub/+gXu+FuDrLl+tS+5pcwOMbzYk
zMr2/5w1ALP8OwGHozDSW0WKRi2llWG2fUlE9nRSw4rub2zoWspXk/lRGCuPdd7mEO9sWXdlCrkp
QLm+/xvUmTXdLcIX4PcVtuD1kAd8CLwrfnypKstVF8xapS5W8vtx5LXQDhusl6ldqOS0oh0Uzfnc
NZRGHWLU8k1xgqCkrFz6UM6Kfx09Oh7Nc/wvmq+73Mb3HAzylY4vH8gJjfjxoCBdU7qml3okptdk
+eWp+H3gOKtoTL1T8oy+DPFItgvX2FnYGobaj6d9eJVCc2062mevaHqmiF3H49wl4Mk5r+wO3pSp
EoiVfnLsgvhCbwlMOmYCficVX6dDRGA9iS8XkNhT9URSVJaUbyIUs0u+mLzmKlcCII9uhw9zWblF
Cheu+8Z0Cxl4H1WVPBeBrenZ2pwYaoENn4i8c8z3i/GljpNx5qqC/H3O8hejMM6zs2wOOh59P/XZ
uKHpgDBcvmUi/NuOf/GkylgTnNEFnMCBH3D/Eq3CBqrmLwHetOfkQiekY6gj8RKC5X/9JlX+C4Mn
qC2RgkGtz7agGVhiwe8fMIQprQzxLPyQBT9YHVqMOJpLlBW5giuIbwU5PU7JSNiFOS5G2Jy66H1p
s+buTGYmO4eps/VHatSw0gL8bx84vY5g55YHVXW/C38/iq6jyYNNTUgFPfkcGlwffHQtcn9afz8z
B79vfi/WCbyikg3bcJfK0ncprqsw7diKjWY9wLLI8nPGBddw2R399mENB4FCwF8I6F6cPfq3Dv5G
zADUQZBlViV36Y9ZViTgt16EEWBFbtI2YdSePwVlbso0htvulh16Ed4vkM/rjVrKfeq9SryZpc3p
tXdisdmwwGZdNfkm9kLXAmp5STxquMfk/tYFHrLhRKC6Jas3tLAldndontxvPtlu4gMAYs1SgJ6V
qsUyMtaPq18ZYvYLKGkHUlAxnJUTfWBjuydK8tMgV+J5jsscB0hQmc97HAn7Vl8vEEkRVXUrlu/2
w3i4eT7ze9T62ggKjDLupXZ9ei9C38NwX/pbt5Fg2PR9CqPnMdGg+gYrVMThMpeZNmAYWh/KMh9o
C9cvAad6Mae0OL/h0804tF1nssj/Tqu/GzHbjyJLaAg4jptFrgZg8GHItpmv27c5vqcOdn+An5Wj
KXdPJUdk/vTt18IuRjOeNP1XIBmjHKOEnjBlBCwNY35pUbD/tNQC1K1WW2v4bIWDXZRlLdbKwHf3
FCQRb/RhWj9qO+QJV/wptlrWRBUerY5hqmUfyupiyQtmymy28MdgD7aYouloquJzHySBlCRshUsk
gxAS9tj2KyhR33LKMbWJhxg3GYosDX1F3zjuTIeoietKyeU000C4K6P3roQp5RKrFm+uGltvgzgU
/n9rsqVD0x7lW5yWfrgUYbaHvcTbzgmbIC9lS2hUYqGLy6n8UOHU77C3w5r9eTw1nMiriYT6zzdF
8+us05ZbyQOBUxmoRzjSrMHwoeuXlETfBURt9mJ4k8Msh+VXHBLdrssqaMPL3JoNHB1tm8xjCh1R
lFCzIRoBybt+GEdt+O6yqdscQDe48gA0ZhL4StncG8gfQ2dmvogJLFO1kLclVj+vqYXkUuLo+xLE
NKF7KOFevzDKvoZ93RgcEWUEFdcQzLFcG5+suTXEidgIIryta5baSZBoBQsA6aQq4oE5a4qN/bBY
LjVRb2Txc0kWAA5nfm8fNfKOHpw2az60vsr/s7jwRnyZuR1HusLauE72KiN16BjcO9+eeS7l5d+a
ZtHSQUcxHh5ejVnJUnpwz93fyy55CNR8Ky8fLREu+LrofSnuZgp2iEHwrmkVjSR6q+ghyPXmhX8k
nabgEa9TmrqZS3zaVJfKcE0UlRer+nRvwGeq8Fm7AUFXkUQqoykM7FhUpdJDeeedoEEveACv9til
W2GhGvHgU2W/0KeaBGP5pmABXnk+zeMmS6kQANgx3yzRvPFMrd90PU0dDz+e9HIfvXZil07luP6z
dUdPluQg1cEPkVhNyzRFE07EosFhMi23Ua/HrYHiKoZSea0ePTz7fDn42hrklmwXU6buGi8HXEni
CvbG59+MqkkJ8lMICJFGBC6VYkMaYYUUCSq1iNh4wvvtTXp44XXuE15eyL9mATCeI3swSZ/JGy1p
tm+BNbHSmKIIUyjuroMq8lmF7Bf6c5WRkM7RYh1P33Yqin5sqpPQVSUoHo5h5wmHnkjT1kt+aNOq
GG7PiaeF1S/813ZxVHLrIIIBSSS4SmhnMYB4OoQCtk+7+buNZMDXMyHBtnjVBwg8AwYo/D+AJZ8X
krFacjIA0WfPTpzN91jHtIuxHbHY0X9UNX7I9hUcufD+WpP6LADf7wTM+ytM9mljuspTB4Ugoa8P
Wgfjt2SQjK+Nk9REF7/rjPYeqiLWr9pTJK/mj34h667LcXz2kV7/ydp6ViiErY/afVQWgGiP198w
0SQOAgcCTrVY06Ef0PGa9fhpsnVDu7Yz2/hfcg6zDBQieMevj3llSSWg7kJE1p2IJKS3a1mapokR
HQ4tAks7b8ApcAk0x9SKuiRu6NDHMHrqqCni0h0QdCWN2Zgx7Wk6tzZ5DsitZ58AR1T3X9rp8aZY
TulQB98apD6A6ggI8j/hC9KeBbjMhTOlIMvdw3Snt2wNN63EBL5mQT0ppQjjyVJjx7o7CLs9V5IH
9pMapMQBjMF6rOM4A66reu56SHi6xXLYBlJqdCGrnlqUBXL8gh6IFn17PWhleOzmVmHFqT0yFtNu
EP5BKaCB6mbFV7fLKAuac/gXlGddmo1G8jbnIWUKBNZBP8nQncDQaWHcPvVicJ6u66hY09AutBg1
rJByG/AhwI/AHtU53LZooFhfXG1u0P7g2jkxXexcoedTKOfkZb+10ot/SQJPU9LRhJU8/cjxNms+
WEj9eRlsCrpew/9URGK3cKTDxWom0J60cgux+Gv03EpFhoX3jB4xWy9/844dYF6XdS13QZsl3341
CQus+K3jp1nM5LLi8Yp8VGVqe4B36/5Djq37xW+SiczRp8wtlnniIgDRuXcw/DoQhIS68C05hwlD
aDXoqaxwPJnWOu5KV/szszGEep9Nuk/TkIAJpK4bn7sgU2IdvDRq7sG0x8jGiQHbDNqQImmFp3ql
0BbKupniAFzG56/nMeCKSf8YWI+2ZP4yUdvM48D3Uy3jgzj3OQQThDQE7aDglN1Alv+MvyKGiUek
gwdTuOpB6pjOzm8ktmq2eaMB5FeOszwJ8T9+Mq6QdUVUxfspkPon7iM8oF6ySp75haJvEq6dYerp
7+af4vUMlVJTtf0Pzo0jwD82LvQ6+0pbGSrIK2JqaCE80r/XgmmiJVsNdfMyLstS9tmdrFFBosIi
1blTO8eLCiHWrEdK+A/jkhulq1fU59QbrjR8PPaWeO84yAl4QRAHvurIMb5wAjfdqCpT0KPTl9in
E6RnzlK/2OxaKZP+5N/fiTnDuZ8U4SEJ6aObXbX5JdrgEpuJJt26JJyPzndP9cTc6fC9uzsLBRYr
WqZCtgi6hOZTvj/S+1AJvioJA7IunM/nKdMvGmw7jO5uTodorQUBwE8w5t33/6VfIFny1CEcALQC
ZduP2boFtHnP94eqsAivEuAcVvETVvWP+vCFXndYo96kJ1eel2dt7zy6LXS90w+wxGacOckie8Yu
vJ/WTkfHLtY5ufU2aNFACqdKfq/WcY9qaX9f2mnr2+qWcRWvkZ6ckx1qNaMAfSCYvV5uCqfTI/6/
XsXZAuV3t9dFkNlDCBDEfCmo7MgvRfup+goAxDdRUEj/Gdc+QCV3U4HuDoPZTgOCeF+fQ653BvS8
7E+XfvKBGwziJy0/iSscryfl1oN5jcFySuLID9yp3IthEknho4pa/8X95jtqK0IRqhIlAIVEx1k3
Dou/bocGoNqJCT/a1ySD+BVDG2/LUnXlSZU/pypQnT7doboS/Xg+kVr+oktW/iqP30aGehrD9zTH
XhK3EAsPk+GmCbCge1TvNy3v71v2Lmni0+44phlbatewL/nLmGrtIZF/oWoCLxtDOA5lclRjKbvK
DPHGX0bx4ciueX+D07APz1ujg2Ybu4Ed1i7JBi0qDCgNDPfDlc6f0JIn7rlIk0lrw7OO133/XBXC
3+7+bNzx3xss01fHU4d2mxmgVJtFpt94e1rdrNs8Q032jooFNtcpgfaPGJRXJPZYVdqmnHOrVCCV
Ksa5yhIsqn2QIAxOESx6Zx+SbinqzFwFoN2Jkmfo3GTaByuKXri0VJ608v/JRD5PKZ/7mpZosKR8
s9Xm34qXnqJ9YmX8tTw8LVvRs0jxVz4h8EgYiL+jlXQavAcNPkmqzgV43vSeyVDFK8CHeIVnHf5x
5Ncl4NL20Lr9GS8y14oRnABCEFO5PKUqgWrFpX4xEZV0bCOdlku4Ff4/dDONIeeHZtum95e7Zo7U
O5OT2tLYKd7iU/6asopIYXRlFcSxuBdctPmuRYALGDpLdQRzR2ZKQBQ7n+tGHMWMHeg5JIWHyLVT
f6pjpRJeI4rUgJe4vEvSU3hxz4FAPTUD/Pmxvo8ixeKKmuQt9FgNN7r1Ncskqv3nKalM9t8lZoC4
QbJHw46CNBP9rkB9aO2J7z7Hf5ZsQUO6R2pTl7BLhtLZ9IMew/yx0iA6/CpJoPrBpF4xd2z9qoA3
rueIzIQ6ehJSZwCatFcSVQ/oU6tTFOWq4U5vLBE/h9HXYx6rY5Nd3bsJpvetNnA+rum1SDxGE/yR
PwfJb2e+i0SWhhC23tnbcWXyAJ9zV9qQ9gDo5kfOh3KOBaULASrv2fEDKEUvrIfolfZQWPKXS2qM
RDNS8soZbP9CeKJMehSnYfB7sHo078UOsSAWppUDDJDiM7QINtE6xGAbvoTaclXFdo7WCW9nugnh
O1PZ/GHa0q9SF0yQHcm/11t2hbjdA2xJ0aiOwnqV+uLaPEgOLNkCQH7Ud+FoSkMovUhlIGQ9sQ7e
78qMUIqHAT+mA3wqeetPBTgt613WtaR0mWolvU+soPE5jxKdIUZ2TZmIkm8aKzVQV0iVKxWWV6dn
g5MICAWvoynGf7dbF1GI/bnsHTGlpFBGfwr0zuKLRNTEKb/52txKwXFUTqmaYKQjpdylIcGJY3IT
xLV44/rR2z2eaXqFWzYat4ZSzUWepjZjedQ4N4+GUsYvsAy50ssyef8Q7nzd2Y2SYWT2x3vFe1Mw
hq+i7RcjNo+ribboVvHOPlgBDWT68wNqmwbAPQKAN5SVAWcGSe0SmnM/OIRxhRPXtRc0IuXvjeo/
FtQJRIYNumx3VVNylLYfu73RnGm6SgnKCZVdTbMMnz/HhoP3fFy+Q5x9JetaSlkxSDFGTxpmFZaN
jHtWfxLvoiE2VQvjlXqnUymLa18dnoAMPKQ8VI6zfXDIWMTZTostYAmQtm9RFqq1XlSoJY6Os8kQ
MUVOOLeImMr/7SmygtQ2CuR8mWpesk90pSxN/s0WjbIOihCzExbA03hm6fp18IycOFduo80sX9WH
GW0JoY5KtUaSVlFufSrAkhCzYtgnC7mZBpAZsA/VWWeyyh4m+ETos9MBmsFJ/HczN/GGFFJUKphb
GxWtYgCyp3EqE4Dgcr8LNmzPlK76JYj7hRBdW6t5Ghmj1hjniawYgR5QA51ZfdAvjEGlPHljw709
Bzp3PklYZnXaNCT/EV/Dt9fGwpeG2CKg46QoFoNjxGi+9YoTIFFKsdQjLOsPL0juU7TyV9wyVEBu
fjDNF1u+P6kLQ356YDnIr7DMyDeFh6SyfjmWJwHuHpad+5G//q9SEHceO0GSUE4rKsHlf2k95Jnd
+Jsm4u0gKre7T6keSNFgoxHvpgrBQj6RCi6crkRsEKDsPi7WeOBaLho7xSl0cA56Ls1lDcys0XRv
aa400jtbLO31Yg7ekBE+hAxlWM/n0B6GgwzRTpAMTF0bxh8MuU3K0CqeMGdeMmlMlr1cIJYyczR4
wWP9gpn20QdfRzyTS0zUaR2+btMYspyV5ggUDNPhms9Xt1UGKp+vN/u/N8mhLzw5Q6BV2yAoM2ZZ
4oX3KB/X0R0n1QriovqpspUY2+J/sg+6ZdP2HQFxAlOkBZ3Xn7L8FeqzuKYes5a+V29FIkLONt9U
C8Dslf2a1ALzY8fvGQlGqPFPnJINAI4od96AlrYzu66piwwyV4lfvvH+ee9p7yl22EnMgCggNHu5
vSFhfYvb5lyuYtVpXY336GScAyo0U/YIVrOQQ3AkP/zQoL83dCP/NFjIsvenyqDoIPaRBOgzsgef
YLFS2JjGoT5lNTbBbRfmdulnl15gVcRFxpvJSZeQ+lrC5SRDYl/RBi/F6XacLWZAT6hItQkh7dyi
Q/jQoA2Rsgz+yjedgDrdqrbDUS/X1gynp0UGm30bbM0+axVKxiqmGJIyTu/y2EwnuqWFxBJ/IDeH
mlA4IqC+tXLm6lX9D3XGhiw7PpTRjVMhYomD4/SsWgdkdZbXWGeqe7BU58fByYf4JSEqYwyiOLaZ
fDLsrAuGfItmwvOGj9gad5V3YZbZ9gobdtnAV+Jit6un2JizujGKay0hMGf0DWRc0xe9TG5XHLBX
Jj8BwYrBT6kaxZcKXAsuKxDffyVCb6+05rr/ak8zRz3eBGPnD6Z6AtUpoO7crC1YXxu4a8hBhsbm
EE+bazvtxl/njO+4Q9L4uZbmfrJTIH9N+R/Eg/xRfq0Ja1donGhSg6s8gudMGpTVcoLnxPnrsOHy
VwCr78zRqcgQSWoSsE0MjhLmzZGbbwwk7fbMmRFf2XiwHeUpOOmsbU6orL1LIBd/6Mr7GOZboTFN
DnyqiHyjFZP2SGWTsIGuzH3Fa3rB04pIsnYNkFbRTTQ9NUVfGNauS3EsVWOUgsv9I+1AGnXUqxBU
Vz4oWuqxyOR2NAwm99ldm98scrQqm2DCqLRMm7wHkKUylHjR8WAV0iRPkOGeXneMEcXHkH9fZNPY
10cDuWQmvAeUEPhQQ40uMsWO54PgDIZa/rKmFjBPKc91p125U3Jaz7AtZV2bED7luelGqVWKTz9G
JTAa/nnPxdnN9fTx5yJ+oAhMOHZktB2Sq1F+sBCpPrjwnbXg177ng9lZD7JURqklxiKqOMdHVzLX
9U7o4BNUAKW7I2Zf331vId3tTUEKoLuz5eyIvPVbbwlieyeg/9gxTmypBXYsrWE9p8BRXfL4+h3C
g+SOGOkq6ZDW2nbPate5/bs1eiDTegWEH5PgyzFWvCtDiLdnHWaNayKLxMwVcya2dwJ6jxPEYIVM
uheixVF3BrxL6ikZGE6V9A5JA5J+6AJ7qBngwqRbuQJfbUv0dJfqgqFoVjCINEoveD4xfmEy8MTV
ycR1UtGPDdBm17FI4AermYh7Tl5odegVTdx7z0s43RxOfkNGKfw/yLRbJWIseBLateHaJY/LSXHJ
+cYOGGoq33TUsUWL+WDN5FRThJUtbxlPxozXrSHeABEULBC9G1AXTUkunwBRmAnPMoq8ygJaw5fz
SRj9Si516xmI3kqqQZtiGg/0t0pOdk7wBAsYcFXz/94tx392KBJQiTnZTg3FlZwuZw4q4XmZxfag
AJxZ0AnIweyYJy8kQsO6oHNdv5CI9AEGb6d2JfTFHe0ia/Mrtii9UjaqF5ncugW7l1jF1ZYksFma
GxHBHFkObGJOMIgRSxpKlm6FadIzPy4+rbQFd+U0niL+vkn1h4WTnYjnnyGgRFGSlv4FkQkAlh96
zvvLOlETIDFXoEHPNlzKFggMITTdvYqqSL0V2prXzLMBRDcJA6KYSYOXHsP78E6MfaXXqCrl6rTG
iO/mSIBoJJ2JHHAdn34MxLz5XdnsNzYU4rbqN7q4+cmK114epz37twL6lCSxQ3YfgTRwLjzfaU5q
sEMQ123XZWfyCidg8tbyFyEgQ8djttXNV+GB/Yg5kUgpAuWMDU10xN/V4dJJRp5ii9dxL2B11uhY
p0ZgFxceI4n9ThqPjaXOaBQF2Iy+ymphQTi5YWPzsr1zSY1vy81PCuCaJY8Zll0PL2C82Q8qLAHZ
cT0Pb6wXNqcr+Iec/nuIUu8HfoQNqbXUEWOyMfTgQWMuRUZ2nVvGCVa7ZFxQ2wmNK5H34O8UM6i5
D99oj9FOQX2+qeRL4bUo2H+5ZWsQ8PVjwkLSGtoRH+p1josB5QdfihFx71eb13CgYV7BrEms0XHn
Px6zZgHcnVOPswTpSTljSpUQjVr8Pm6e3QR55h0dtudP/xOh37m/QtQ4OivjklbT8vDDtMM9lsp+
FfKDXxKo8Gwyz3LBD2FZw2xmPYeOe/q2TPQcHgHTG5hEBhdipuKMTXb1ZuEHgL8xWWI4qzKeeoPR
g1/v9ScP2mKPuF1jLE3i7ljqg1mV7aLPkXEL+oua209tQJPdaqGbn8qJHq+k0sGudeugf33RPV0z
5SAyDBIfyImwsberELPunOjhPXupPeFypLK/DWxUkV7lgYows9KAnYQa4AsDgi9wKAW+TxR7FBhg
nZ+owrpNexUJ7OXX/trBI1T7cRqXAYdw/dO94PY/UfW6Hr+1lx8PLA0rO5sZTpjDuAfnL6wmmlqw
O0t6cIZuFV/Pcrd20+KanHwSpJYZfj9U8DmUudEJlBp0Ivj5YyEYLk0oHWjNLEiddWdZgPiWAkfo
2thSb0vxpFBvQEFD7IGUYFveQjoWNJDDqJQ7WH7TQGkEIXjIoqH6Au0e3M6Mu/X86ymnGK5a40lP
SxAPszaHLTeOH/Y51OjlguT1o48CbFxrzYVnkdoJbZ5/q/nvdL/AD4qUyrvLgGHH/rdiJlUISnz+
K3fPLZk+gHekE41N/MHScgc/z74jhvz/fUflVJ4MlBdW+iGs8Ob/kdF16nKIZtZ4lSk/RSDkMv4K
d0HJi4oP3ku+rxv95Ravac/zG/ldN2fUdhXBjNUPfi/k92kLbV5vTnTgiloHapPD954/sAg5BfgT
vCSpVOCAC//FkkHLTs2t9nl+WcHrNDAc7U0jcMpTPaMST4mkMYmZwk0bGWQ2p7mt697F8FhIVhOq
nLiKUtIsR7g6SV244jD4iidHt7wyYoKvK7HUGU+oJXWCBrkV7DsFZad5JT0e8jh7UaRBivC9klHD
u+y6TwpmAm9snSI++R8PXIfcskY0sIGwocyPIu0NntNj6ZcoEhCngx7c9eDYH//PXaebYLK5JTYH
IetCK7QumBfvGUsSIe8ctwIVhAYSkfMzNoj1fGP0ma9/qesXZHR35y+6NjT+ATmPciNZPxXiaeCx
/cVIavGanV5o0zvGqY87nLxsfd0x99sniEtj/9WDXkLRnRs9CZ6i8WsjaaAhBZHJX/o4/Hdz3whM
7+NiiJSpIPMc+SrsESaRB6QQRzjmJyNr2AFAP0hjo7GHIb+AwLezoLpOYJrkdk9DSBbCGHiLrcTp
o/vQA0IjXQ8NLVqnjQhfTcLMpaZXiT1YAOoisXv0itbGQvTcqkm68oeel8Ckaog+ojktnBL0XOyI
ptU6Dth+FAKUB7O6ik7FkHLYuhVFsiGcIErThI4w8A9atXadX02M7u0m1IdM6xXv93VjHA4er7uc
opOPM32V0fXlFqusYSSbX2y5By1eKX30nSZhAua3o5kJtuvQPtIhvc3Jvg5JLfS5NdkR5y1kB2Wu
qaMQxd1PxPeG/CJObFIR4duBP2L7pb100dqLIAYv/N6intuE6bgSE0S+EgcLVuqz7XS++TvXsSAV
iqsPfMRRp9l2RALuuAwlDqZAX63i1J9LJSg1+vFE+m9LELafVagV2Npgd2NOEDio3z5JuYVoY1J4
u8zKv+xlpEPWYlk/KTQqqJqKy4kSspl3f+SdNGek+17+dhQDA9HI+nDfuGKOXFoVpBhtZVni+xcE
JvnJKADqbZtWTwBM/eBdKey4s7+ZTWm63KYqoAY3eveL0idPTDoK5rZL06j905veg4fWs6SDbXLa
8dtvr+FDO/FO8JpoCJX8IwcDuBcVa0CmBrQK5hpDJWjxMGEUwLgpyMdLRxE8X+4HhNzugcldIjKU
Mk5DfoHWlJDpRGxt3UlJwP8NrZMwWIEj5bLRC5p4u4D/fMAStxYYDzs+fPU9Tl2XuvrcanvuhJ/f
r/QiH43VOUCA0dI5+YqM3kUjwJoFHi24SrzmmG6gyuoQFoHhedoV62xAj8L1xURJ+Thd9vW6I1Fw
R3nB7Dg5TWUWXHij0GBqAzxYGi8cAc1NnhCzIEzNh+4nvEqWKtts+b8YvRmlrog7zGQ4UFQ+pd/9
AJOL+zWfBh/8cfggxEGfB/BckAWnoPgFqaIv90plg/3OBWPlbHJxypGXMMTppKH+VJPj0S//Ax81
pH/OzMTns68Rpckk+Wp2aoeMuMJRmpiqEpWaPQBIjt4EUf1IhGmzze9RbDLST9h+RQVecU9Flfyg
WlV3PIoCmv4jQx5BMZoHSf1pA22Hkspv7noR1z21SSPXZbcnQJInsjvr3WDZBnxbD6pvq2FRJhvy
cd4Ee5tBRRB7kuJKoJk7zWFoJaY8ujT2YQc/VntDSu7fplNW83sPkFd2a3+KmVI8yeJ2wdip894Q
/KHQoGgyK0oRk0uedA6vbChPHrXxPruj1Zy/ElWdmieejVvB6ZoMDjgfltuWZ0iIcOMN3DWntJNH
a52HlN8ZqB5JI5A/7ARL8wCGBRaKUFe+CktHL2i1m4wi9CL3Zus0RrNKjoCeOQJEhZUFwomP72+B
4IZBguGabkCPP2C8AQ/M1N6XHAyMi1NB/r1BstkFKjg+TLxdUbyztHNxCsy5OBHpcGAhW9aERFyu
XNjEQxm471p5rkPnEh0OsLP9KdjBmWJQoaIW/u+/hTQfRJseWF4WDvIfB+uw91EKm5Ys0NyvL8kY
Dyb5N2+vJw3Dtj3RqWKGtW62j+kEP9iR7CwIBMX5zMumteunQ6BYwvC9+PqJYBYS2jiDwTrcQZWu
eK0O0YO8xYitF5pzhB92b3thD8Jz9mPvLvfHgWOQn9IdX8ZifkazRfodFmQ87HE4Pusalj8ZQAM5
xcsNZRuWg3UHbrUb1uiUfzsuxhsv1c3DpMbFUKM7gXIIOUMktR0PTGLm2k7cU2qOScHxK4b8DCc1
rSSosdEN/kK47/mV3iUetew96iCKjJbALG1UGHoVgrUtWcicM8T7bT7H6ZEtD8jB6hK5a0Nj73gm
YlQEN7QP2kc76FDQTXYsNK2KtLNWgAjw+E3nJ0/+PRrUwQHtvNx478lZFuRwQb7TkK8bNkVe7Gp0
u38iZdLFO8Wufk9zU7x6ykwnYayIc40pLMEtpfHMIgJ9qHYgRheWMOfEO99kxHmM6dvZkv09O+Qs
Q+vodXLZ9PLLJxfKcxEnU7LRZieYMnSS3L0P5Zt/IQBZWnLE6wqeaxemUbWUD4Rac0fz2ZoPakwY
RVSHj/phMPh8zCHxazksGeREEhg/A+dnnCAMZYZxFYvCrU/h0skOKneIol4F5m9efkChlhUlqun/
AKYjtMVUPJ52jM9oW0UrDLz6McLaZH1Ou2t4VAtgxWH0OPheEhQg3NNLuaoxNI0xRqgSxWIrGiaA
QFbRLf46+QsUENxSt9xXMB7orP9VJJ5nwp+LYTvKo4gJoaQPhRldQiWXztC4OfHWGx32YFJePyYS
fEOiLcqCTShBVYNtFMREntP2J5cvaZMDJl+VuKjJ13TIdRrv+cDUXCEJJIRpz5jw0udXDdXfKxxi
LAMPMWu7O1aBVmTGkmt1N4COo65bzgpjcE40tVx1osLoPRG0XBBZTJjdBODphKyNvvgpSpf6SSpE
7YNaxsCa9LnvMFFdK1N4cobbtUsE2eibRK5HWQS/B2EX/vnxWZHTxbkgzvQ/VXpIT+Z8aVEEFIK8
EurjN8ONY8jQFcls8EPddZalviK3srbMqTApO1sN187M0amO08eVFJnBvXUdRsDWqWFpwyPWIOqE
P+Qj7jVO7Gk5jhR61rpeTc3pXybzeRvAwrpsAHqz/aaryPBH0kXNk7rKYjVSKo5qIo2w1bEPLEkv
bwcuYRFLYMv2jCBMxnAdqlE0QPmrS9jpVmxON9o2vaPxbMPsygCDChQbp6Q1ZshN4KfvMve3R4l3
3/M9eoeRfF//AneOA73y05VVJOyhSW0+skPciHYCxiueFJnyR4WdhLSL8zlalYh6+yht/eXNe5zi
5ZEfycRuA3aqx78C7XzGNH+1APKQU2/jnZ0EYsBkDLoVDehMIRYuyzXLZZyne8flm+TbvCxZal97
+8Bg0jZOL8QvTiWt3dHu/A4FULvmyFhgYMqoekaQsgYK2bwPiMTgcSiAk4US7DfQ7hw6nclIPtP8
ip51FFsCiIuIbKvUTecMkEkKSSsbu7XNhyVFLJDf7ebBxQ19KhlhC8OidmSTPb7at1cc2DKwqnk4
+Wyrem4nMjvG8dwuosl7jKB21lYI+nOPnZNRJe6ZgsTDBRh31AT9ZDkTCFTF+4Be9xkWb0WsYBHa
bjpRZqGmSVyQN6rqUn6uwLbDy84WuXjM15k4PzkfbTgyhFSz4pxSs9L49ZErBa+yo2TYKYM+IIfK
NoybxkBO17WY19JsEwDvoX3122oJo7QxAhvIugXFmgu+IedPHXTuxKunLrVw+lUUf4NvbuuJahcD
yFJNKWS/VDCWJeneEwbgMbqGocZagZ5U/gh1p/EbTEpaVQoVO0YODWpUGjVhk2uSmhKKb8CmZPZE
XVpo5ZLXNvXzGEbh3UwKtthdlHhZ3uhnZKfQ5lA0dwAXVWoHj6RLPKGzdA1Y0bMZp0esyKLXcO5h
WlMgIdju7+M0n44as3aNvld8hdrlNZB2hllYuXYMiNyBTK2dZZYz1iukGu/LWkfPKi4Sa30UL1br
dXGvFZ4vAFUgGbZCFAaKW7XhtiWaaecpcAeEvJMgQsnAWzeg9IvVKpAru5wI6L0CaGsoWWSrKcPo
B7F1BLyCWPLoOIcOanSjQX+HDH1dxsITgBjP8eakiN+2cxT/3KAQo4qbJt7z6XhyfpNcs7ioqfqJ
ZPU0jz+tuwIKTLmdG61bPJOENDuafI1o/W0HiEs7v6KkzIsaLY5yXX+oP+xyC68UMQ2iKcmVHm5l
bYbsu+CvUOZUCHGaxX/FLt3ZvafyjuxzrTWcaUHKF1cwcUxIvRV899lR/9BWnhZhjuIUBLG+sMLk
GCoZMpCJoRcEm4wQQQlFD+bZOnFtsrJTJIHREuTB2ynvkxabqLxWb7Y/JWV7bcDiCVSJ+gzvLQoq
f9ZJOJVredoPXA8LCS66LQoBt5LtSl5KDG2ijfzkdtcoRhFdxPJTUXy3NOW/sQXF5OLDnNei3HBD
8yAXkUu72We+j9ep/iyANn+Dx6tCTndTbeU7HCmQEmRPVMq+QqDoaTcJJsuCSpkHVYwGFa/VRB2y
iMOichOmxMI0TiHpi+FaKj7EvUCxOkw7KBm1Tk3SyL8Sf7gsLTyUF7hKwYH9ubXjgPRrM0j8r48S
3X+BBb1Y6uzzGA5lRY3RlTp8rBiIRDAzX5PkbkDnwzSS/wtiJqCNwLhVXu68HmdUcD7kvrfaXA1z
M82T/SzS1/Xz7C4bTiagDLMkOpHqeR1xfQeCscmLDEhm/y/S0RxdXh9cQjHmNlsTkwRxeYsIyEFn
nPA4OwfQM6r/TDUj6Gh41M/Q96NItYLPaKzcMbccTxBlJ6s7cAEwOV2jNZ8y5Pqx107Kaoon1yk3
etypNGjuCFexnoWNhf1THfPYs3hEHRmME4D1Xqb6sT6qlR4+uFBSpDlwdC2azfbZp0JXzIwgns5b
21f6VFrCoC6/WkJecLU7AYkOMcDT6HNmXO69RjwoTTFbDEtFRp0Hkl/fuNcLH/6dT8KS7Jp/TLYk
Pgshb+xnRL3XZoVl9IvI8BHX7RfbtBqK/qaSuHGOAozX/sG7K5hElMYkKIZWIwOz3S1Iofu0N3Uk
DgZJDxBuAv0PFiDaXjWrL8kdPzRvc/yjIPXZCsqiBpZDItKgTmaui7gnhhQwyJrv40ZRumsBHYyk
1fe8A/xa7ES945f9VyqgKKSwWb74eakwY1nYIhzeyxRHF4PmE75H9V+nG9kfII/6M9VaXN7w6sD5
tHcSavwBH4Hzws5djrqex9KYpO5QVK4F2AfOiFX4VvLussneeil5Ppd01bfOYtwSQYiw+xJB9QMr
yxBOyebaJdMr9OVnb07z0LhZQc1vZLA1NEIbxjjbne0icO/fWGEsCDtm6EowjepRCPmF86d8BQ9q
wZXA+S4ko6QDURFp6+oRvmzk5wdSGNRqDBhJew4Ct1D4a4ibZcQvMSuv+M/lyYIWo6exCBKgDFPI
9cOI2z+/8g99iKlO41INcUXWUhKW27XgMfpQWV7t6mXhUtAzF89aXcfDJm0eVtxzbIAmBxb8U+g2
mKo8uu9iaTS/n06YsBAr42adNpeRMyEyvuogpl0tCfiXHqgjuc+EKeXSG+wRgPCrBUqBPduVuFS4
cMMAGokDMhCor2ge02NtZZLzXUhY7grT0CdavhfiPSLr6aX/e8EaaZ0yBZt7TZP1OekE87U6PrT+
GnVpSuBmtQ7cqvOFB9uVbVfj4uXOwUK/6RQ4i1wLRu7aoNXkIfBzXUkcfb6J0n7RpXpHAnsDVOEH
J3qvXUyPA4X5pLbX2/mhb0bE+yqQc+SiEe5AM+w4t8UvNBxbbo/PMGHX96E3t+VsPpKBLnRb4zWm
/GrGQHfHTXjy/5HzmBowwFcnAc+NnCwJccwbBBUqG8BEil+nn78VSGLXWV3TH+xwAl1gbiLl4IfM
wK7Wjy24OXumfvXf1RUMDmgtdUjPS9R5XHCiinWAT+d0gz1NESrLq4EVW0PbXw4djmxl8S8YRafL
OVs6UTGP0eBlpU5Zq8K7cXBvG6Y0TRkHYlKJkuu07ozF66c2S5UlLCCftC9DWg9xmDDM7TeCIMO4
MNCPM0Z08anroYee3PN+YZ7e3gERbHHtpTpAC5/J9Z+BON5vkfOes7KZXQA/UEcdAordgMOHBAlh
WCJRFB8c6qyhK0W4LtuqJ4291fGUB+YLIG883e1MZb0ujDSgx1wBHov12GCg9039fUZJ1q5awF/I
IhApSN+imMZCQ+qvzdIVEEVXxAdEOBHQYkmjCfkyTGASolkhphf1ubAGJZ9ATfD/4xATPDM3ei9a
3JJkXFdRvX04Sh37KUfOw8RugmEwXC+np2aAnakq77hkiMZqYB0EB8v8NLYDbgziJfbd9Vl9x21m
+/YOL1atuJcWNBn2p6zrkk8jN6tHxMiqcVK3im/25/QD4T77iOM15DenaN7TI0EDgk8XqAghLbFm
x169uE1Cqp8snb2oak7lW/5+5XvDoXPsNWrqsxsi6E34xrdLF/BR/1d9od8CenyNLmJV/1XoBEO1
u6sUAeaYfFYfdBhzW2UtlQgwAMdjs87zAadGrG/22MPf0I8R1EGxu8cW795uXV4IDEBTmybm+BWx
rYsvLoZVLenE36rEV7f1XG4Esbwm+DR0i2bqTsnKZe6tH57jvnA4DZ9HqkInwxWOv4h4bjj4mTtR
eGBB23x04hHnmQlen2JiYxXg1ZVeAcoAKTjaOq1YG6UwOyxTTfKSqYTi80dNYwIntPydbPSrNG/K
Vjfo1wGovZVYqO+TyRocYFM+dFWrGGq0bU5XZL2Aovv1C2qoMDr1lGpX96Y432aObZePu+dhSPA4
HwoFOM4J/24bTxq6JB6Gv3fwzVCEWPbzEqWZhYA6whCjPIDkgkRtwkj7Rt4CTJqEO/eX9w0seU0Z
+ai5jy3+6tW4Q9fgEMu0CzwN5NEdUjNgYpKQDLxpZB1/ZxTWQI2PkvDCVu0k+W+UZD4vWeSUePvs
51TTYUujtVdd+JTTqdm12A6MkjdQHaHLR6+Sne5lVdWtPDfPr1bs77rIx1KEYHzb5D9IeeVge589
aaLgjFyP+MUyp7AebIMMqmesqtNq9b8ormvixgiUCzDhEIKAhW+wntM44PK+Mecl4BaAp1Scviyu
/WiaL371FSzZ3qhUkETEHUx45Wc67H3tilz8OMQlWhDFpWZBKawHT5sbjpoZwDXPpJMzh3sG2HUC
NfrSbYg8pHcTwiuf61YHMcizm3ohzMGzB3qk4YejReDtwHhKCESdCUJJu28Zs1/ElmErGk72Jxhg
8lB3VbnR4n2P1D4mMu5ar4BERdJ08TsbPj2XC/prG5zDIDJwLm7w6a4Y/U4LwUfCscFMfO1vcL36
BJXA2Td/5FW+L8S6jhimLUs76s1rpNoMSxfrWBOXGl5ci/yQjeo9VUGwmyhfEE0+v6qMnE8rNGtS
lCxyYYSxt1Ahm8W7sReTkYpdI40WY/cxun196fUJjCV2hgjK4v2ejugNB9/sz5gsh9SAhNUcsPnO
HTgacRvm1N/EoGMwetuS0/gf0NG5T4AAXkNitz83pewoTAxldHGnWNXj3ZX7PWJOyKYbIvKzzFl7
nOCqRF5HWyw2ZxT7f0zKF5eILwe0bJEv7Y1N8aZiZd7zNdlK0wQBPzoNRETGEkIMTpoNcNTo8JyG
WBaZ5dxQROXWco7KPdlvkkkPKh5DwBHCcvTyzhb4EF1PaNF+R93OUaC4f5SmVDVPZ85ucmKw20+c
ArXw86H5o++weJchCbOMc1YgCgECKTTNUhXwx/O+uJzKqMUYoHEb9qiCy2q1O75vEdVP9FXeY5ip
i8cYJpzV2/DukgbTE82xlnSrBjcPDZgXKNTGkOOt+5wrSHoO5Kng90kiqVn0f2xdL4NcHOY0NcBO
DnmaNqZPTK5PdEh0yV6H9tBa+ia/9/pdO36q8HJhSaAvw+fzmmU9I2IRw4EL06jFyht/Hksdxr4d
tLFK430LxUkHDAUA8/AVxc4ETJmGlLsMxtADujpUF5utYLmW1lYVDoXXKv/tlE2SIy6bSG7LmuDA
txMlRExN+fGKQi9la1KMgALaIqwoEQV0RT0bUipJk+OWpiHoZ4Nwxnb6RTdzJk+7cbBAVs9f6pwG
bFf7jgwL0ZL1EI9V2Cy0kaQszN66PLVnLgvCOM63MCko4BFdIA/8ZARxg30pyqfHQGNq0v7BLnV2
9A+/sqN2dKV7OUkt7w/i4BiEx7EFSMV5+qN8NT9Kjlqc+tdJXdtE3h65tpIXl6LR05aHWXpKfJgF
NJ5mTUcRnEjcImesg0+V5ERNJ/1vOcN/txt4VFLfsI2F0eZk3BLUHazLg//9sXZpih6wcdEkN0OM
ntmQNMKMWieYrY2Gfl6F/wjsJuKzkxFOROKhSbE2E0aByh5ngWpwgXmF0ouKIkQDkypkaS5662Tg
ixaOThGvcytLoF9hO8vlp9AYSayeX3e6uMVYmNPU5PkrrSJhL3Biq4RVorT41nPv+Cwho/HsiHD+
RSLXNNy9ozILjsgEhM7oANuqQU5ufi3KMIO6OvdAT36V6rPhL03/nJ/AtG/0lxlCR3DVWDLgA6tU
zR+5zYaxB1XmRVLttpPaduG6Ri0wF+ACWsRocBlosiwoK9veHix2+7TtkXiT6vNIM/Wc+yoYgsRq
vi6Hdc4Hzo4aaGb+nBkW41yoWnGesLSGRDGM3fDs+HpN2eCgbUjipK9Zc6uSizxS3rSkorT8X6+j
iVoSxEEiyi5pzFXpKukTK2uPJHVfzbr9LQAtB6VWBnh176zmGlFCBvOojhqzmY6lmcmqL4kdyIqk
CftDgsXrWRjKbEDLT5IsFRfOGYH1PgnQ7DU6yM1gW8vZT0zex/oM5u0jp2PL/aK5T4BfcWNfNpW2
HQw7TRtOx3HTfTGGLZkj5vgyGbVkFN24i5sEuuthuSNwkUz0D4Kyv/o7ON5Eek0wdoMnzOj+Nmi0
mL5Uq1YrkmuVHHPsKGkLBbrEIXr4w4nozxdq/D4T4CBs8y+xhCevQJX5r7j4szMDXgapMs+2tJ/M
LnMiUrHegTNTO0tFo6hI5D7Pv4AF1+YvpqyzsZ/Kh5F+UE5+bKmTwErasncFoNabA0q+p3+oPAWe
29HCFw0K5cyoa54EvssoOusrjfhX+elU0qhAQZWLrOHuzlPvZvpfwGjfZNUUds0+MEt5MQDbOdA0
kQx+wEzXyewX8wUFRmDn+i3Z4tEBI20MXwwzCRrsu+HKRjcUURQYQur/Um+VWPcPiPbDfxJ1Tdye
TjZODF5ZRO2u+c6sNXy5Z4ZQG1T+WDIga8bl5aTf0NUFlXlIgXP/7jm0oApPNNXk5a5XteTU9OCJ
alm919E9o7H+hNiDMBmDioqjaVC31U+9Qitwj1DyMIBC4G41FYXou1VqBwhMiiYF9VSq+8JOcRPG
eZpIq8Fn2+Ytc28RuYYexbubfOKiBe5+sv0xqlfJej6cQhL/ksD4mOOJ19JLE/7zk5ZWHfdZrIIh
jPXybaFQp3SWxzKP1E5vrTWwJqLadt/D6NCUA6uJkUMnw0nldx8/eYvZj2R6QICF/Om9s777M1yX
mc2Q4v+YgHKKtoK5wi+55iZjkDqNAkYK9NAVOhBRaqxoLoJWDuMcHCvpFN1D++bGCzaBzr/6xajQ
hfVIbb50uxGLg+TIPK8bVCQkjqueAt66V5REiWT5u5YuNm64Lw4rJICfwWS5YudKO4xOrplQi2sA
ScLNpDUEbe7CYuDg1PNd6L308KiBROajpQgHuEHPL+0Oigqpk/Gmk1aF1fqVR6Sbbf0kckrKifa/
nPOVzjJRtETofKO08v5MN7XyKe0BwYwFIIhAzhmSKc6PcUaRTIzFJRel42fjSLgit1vGIrQE8BNY
HcMRpxoU2rpUKbSy3T1pb79Eis1/WG0tVpUdWxQXOKxfSMXseCwF8Y6K8Z7W3ZoCRpOnDGg7J+Ck
Sur02Unb2nZb40SQAs0/MCbeusodfn879xkOrOeSfqTvuBUh9Pf93gi8EF10oRtIcj0kfNJw3hYE
rlo0so8thG2TaViaUqelH1O/IbjLUdtCDeNlFlStKM1r23S3IGUjhGX/FhEXhlKgD5ZquNwnDYrV
9J3OHDiD5obSUcnrzIMzWN+WCktKpNHmpbD9ZmPb7kzo75u9RRdyXYhp70nLDSgHenVHPYjlUHh6
9e/mn640CaAD6++PpJRhjbSLFQIV6aodjc6GZNR4tYq4pbypGThwKx24DoiRiAbxEy6+e5w3dlHX
r/Uh0OPDJ8AmR9SlJ7SWqqsatGb0XZa5tOW++ojgjipJsWNFx40mhdHAZbEpyuWoVh490R/Ur9rD
3rO2dcQPeeglGX3Y5NrrBZNWiYmIMueFLDt0M2lLW2E38QaPX56YDDyz570uP6xr9xRF2befee+0
Pgk5NmMmtolIRCuZwx0gSXD2yyzZtieFgBRdkeHsK9EgB/VqsBBo9Hcgf2JX1+7N+kX0oaWI3uVq
gfbSgc8BixvSpAd+++3dA6yPd26ZUaYKWaasg85o0xHQywOhcw1IERvkddsjRW6el+6eR0w6juLc
jCunmJhaGoUrXtIt/WYab9WUwtYlxVL7Vq97EiwZX3Et0Uf42q8z+X55brL7D8cmfantbICEgeIW
WBD/Dbg/zu3/bZEuHOgRX2bWoIEP4wAsgEeXKE+RjYxHX9EaZRRqMQZ9hZ7uS7Q1XIFq0Tc41NJz
x2BTlkJkN1cb5mJFp28QseoE2G54XBDPCUV4O2P7bLyfy/0q8ykB2PubbNugSXEunJKilZZpAhK+
R29E7x9yXwgADXI4Vlx1eSeoze18T+YhASzDBbmCD+v4EHIYpSz/tm8bCjxX5QPWc/bqk0PBd9ou
b1jR+AaZ1dfxJi7UQn84k9PaeZ6eU3yjbGfTFufZzLoy0pXMkfbgAqecP35szCtyMwBCpwx7bORY
lL8sOBg5uo/c4SgkOt97aXsMClqxdsKv2Wx5jNga6zuiG/MLD1M48rmFXifQNwG+3UtOlv4lxtOJ
u4++JDgCMPzUlfZj/t3EZGJkMVdSPQA1SnE+gLQ5GHueR4yGwtXQJfAz4/0nttZCYPvwOasCAhs7
BacI4NGfxmDjuYiS+e+wUJZe6h//7ZSwWApXrS5uuckc1UhjNml8Ovog8pEETbOKjt3IjZy2m+Tx
BH9/K+5DkhPKvGq5oFrtt1Q4Jk3GMQt9JVP1dXbFwikXTQ2PkHJq28xWTifNNJtGlSVoPC02InHs
QanuYxqR9ZF+Lc3+btS9rKDqkfNYxEWcoF2NvADaPwg65jYHFFEKyh7d+4vA6jVaAmUxPwvo8K0k
JNJTM22Ofgw9Xw3N7kXsqmQ2V+Pz9NgpwvUth1xms7OwB8av6Nj1R0klgKNGkNPi1td/fmCOG31g
n5osN6SCA1CO+79AtBlWCeEKl5Kz0C7HrGG7Z6GMP7S8HzB6hSFmzkczN6cD0TWiomMmlN2AkI9l
Jgx+Yna8ZmDxC2SGtrBDDDqAN3swMlEeY11u8IzlL6DK4od60wuHJFuSGrk4YWhqT0+1+ruEpvsk
LcpJzlYuEXT0Rjhh03BXffI9MbV/eaDKkNFFByHuPhp4xy2XDvdiAPF567JOx1JyIySUdWYg4Cdz
E8jfrsNocOguOcxeAkcG5frKQinNMJDNq3mkZViywJUaNM+PEd/1k47N7RFVbKKflznvasZ+ZVeq
bXeIqpm7e5p/uF9b4Nx0yBB9rm0DCrZTLuvi1p1seTyTOoO/COZ8bspc8W+xw2DcfWr8ex0r/96K
atifHnEf2piCqZHunHcCE3iBaG/bCZHkficPn0XtB96kK+hfg0o4xxennSEVZXVC/I9SakFLK2Na
KO64Wak5Q7VTp5mY4MD25XGMpiKoBv4Meyv+vQPuCNee6pVomz5ALPi8mEMcdYOSf1nFV8i1e3a6
RVu9ZB9DRIGkSpKNRBsuxsE6M6bYcQCysXerzNJWJAn5BVMkG7Me6iiAXWdP6zgpN5J2tHPU990G
sY32AgCCOeBq2ipjoc/3To08SIPem++dqK4C8S6An13WG+uVd/xpkxkdRS89OFAFljnsq5mTfVaX
1uq67Qk778kvgontBxYi1VX4PUKR/yKVngjBs+FcOyi8nCYEfyvDaQj1Utp1T8DaFin/Me2zmhf8
gyvrtmRjike/gvzAkjqhT15QHh6ybEO8MmcRRhUYgoHZ4CMteb7snqA0alMuCllLBRgwuTvgCOvi
GUF4b08AbecZn2r5+la6kUsNWy8PXF8vwNP7F4EeqotGjMrP4T4K5pR4ZCsNPaA/80ey2vjhqVvy
E2P5+M9ml55ng7mzW7wqvpxp6717BzqD6p4DQwUQI85BjnmqWhGOsMSCVgYreocthX0BkKtXZrAD
bVwOCZe42NRwGtn8uFS7vlk7OmjVu7uXmhLIQ1Ep7PfThcQD6sfmYugSHp5jZvmyUdhl1YdRSiJb
NFgeUJvaaJ0HBltLtanj6pKa7AQSi10SpZ+EOo7qD407YkYtyYYp+GC3803pDBbJHh9O8QuEeitU
geC4FnFubsDsr9J4hCv7VEoucUfZtG3+EuPxxa/YwuHcZciCHZInHeU/OY72E0Y44r94XfPnVZ88
95ZAiN5vnU7Cc9VpAGNtivXNWdit6DVOXRBpNvfxcGh1EIFB+hhA+y2wlKYskvfah5jxRsgLSNWN
roUov+TS1Kvdk/n+iMhaZUaoCypMi5I4cd+lLv3UsXdNJ4Cv4D0Wbcppug3KGsmreFpPr7S0wy1S
H05YcjF0a0irlSe1CF2deZqoR6s8FrP1XvSFknFh30fuGw4uLmNm7+IdFROsM87sbNCTX+jQHSS+
kucKRnnBmeYqCzWESU6OwGlGZ3BMUC8eT1Dz/3AzICMvpT79Yedxty3bIsj87IeCpCOqPGAfzSJO
68yWek6Njv7BCvJjBLGTviCDYR00E055jADBqnsJhN1/v/WiPuJuwcwOqeMrgP9qLgMTSzqYhpu4
hTAinmY3fsDhif9582ivGs7D/tfFjFX/C/SWly8pqqhTvOow4dqUZJNuZvgkJUmJRVRyngvAFXO5
eC0k32mDjT0BWa2oJTFvu3VsmooieaI1JILGSjPv4WmnHJiaKl+7qIb7OwKXNZva0qtIdvzW7FUF
dP2pvRX+6Wbe0mowJfald6liqC5+eB1fG/RB/32zs0qCZJ+WOEbZlSGdSRiKzUyuk/Qa/X9pDitg
h8+9QmKevqez70yV7UWUAfrNOFLOvU9goxGoOC+ZWD9DORVElSK9INfJR2MaZjsS7wlKahzA1bgM
EhXr4jmhKglpLesPlElvx9Gnr/OsXELgpStUnNHNs8I6vMNJ6WzcNDXAD6CmmueUDpgYUn2dndns
7N01AeKjRNhOAqZh6ReyslmBCWkQljfqn1Z1U/wrQ1b+1FG2zydNaPmCt5PVcLnHXDCC5x1q+CXe
MdFCQb66vbsg+uVLoZe8gXgbLISbxpW4ted1FIDOw0isKuhIshcTcUPv1df9bei0EfVnFBzFfRSh
LhJCfN7NHcNIdwIzreLOzeqZUgMy6Ij5Q7pJWAMCAEwQsHfPgq21QO02gqm7WCy4VluYbUvRrf2V
YUd2vNVNK5J3tq1O+Oj+f3ArY6SbenbCB/XZrsrTrUBvgyCElyVVT7rS23GrxQ/CSYcoZstY5v6X
L0rTOX+kpG9AucAojdhienm+G8UR4vo3brjULiqP7Ncf65RQ2g1WZd0wa+gU39/zxap8lSBFPoOp
z5EIqkfx6oUM4+2hWF+CNcfTGsRGalSQgjOqJzoH+od5vFwYDB8yoRMYuC6VY18Wz873Xa6xOsnM
mr7TgRRyMfwyBd3mJ0bMwjCOsnCG1tKBdvIJL+ED7+lLk+K8r6mG7/S1X69eTgvZEgWzHoDUR1ED
6/+3njqACpE+dpKOdrlN9HcjMU3JMigjtxwQcVSP6XqJhVhGiZTC2ODiZuDRPZAqbfNU37DzqNXL
FmwCgX44vhR6f9VUWyGU2SI71kOTeqfFQyzNdW/sQQVS3JtU5M10Tmtbp4xn8ZQKKjgkW7MexlXg
3Amv2Noxl4Ol10jiP9Rafp36G7YgyMuTmt9dcJZjvhkHMvtOTKBCYagFQ/BT/3Sseb7+YScVr4zG
1a4EzaqLB1fUxljiTEfUQRay5xsIfhSdOhdDRg//9aIeAd/3H151hHc76PGmS8p8y7DKJCSyRpes
ePQ1xMt28UWo/V5ieDCozhdJQx7rIz9UWUQBoBZ71/38xE6CfRSheyTCG1Bx+oqVMe6zy0d4oeDq
Zr4NUr5seZV9jN//NPps5x7zMBj6Nu5+Z6U3+9T6Z9PVdQC01IZrb5M/njkI5aDB7Py0yKsi6FDK
BgQdWMM/18AkDizjaGweCA7sp/fYitji1KyHCAII2LcFskYUZAakWy5cTxDsF14lVakeYTRapEJC
NhEGBbCryjTo2+dabq30sIpJSlE+mG745rM1ANbEXljZaGf7kabFoczZDHjaabKkTBMSpwThVxee
WtLYB3IA7lkEaHYsCRQei0bU6FH8oxvbvjRJ4AjkU2FxLZKkuhgV0bt5+DInxidHEsvpNygNoj0L
Tm2DN7lya1u6UKryboIIZMj8f3VBM9XnyI+93aFxshavJtH704KirJyAnfRtGSB3C2xtaVaFSHbw
FQdoDdGBZeX57awPA3Ezu125BLA1modyHwFcp37EB+FyU2d/0BoM2JOZUOAvkKTYfoRbkqf2Ma2u
gS95hZxAvr/F+895KSZXEzl6J04u9KjE2ulqCUjjj8xCpyy4jKMRjZNTFtAlFoCVReM0EKAzBCQp
/4PrLP94CDJnB7374j263GcVFiiDF55qn8tOmc+J+Pl+60OfMMc2aLrZiQp7ZrEYeid2gBRAxGAE
ChakiYBKTsP3EtospXRIOJNsWDNlj2oT3GeKqT83fuZTjDjIFl1HMUD8O6lzRbaLzNZpg+N4FXpd
BhFyVmU/kjdUTRMQa5OkTGEcMlp1p1B/okp1govWAL5tK52DyrCabU+5sjPCQsnD81JuNZ8rLB1E
/1ZRSBowdRH7UvW6MT/Cl3stW7FaNlQVKd8Zthqo/F13U8DnUr1ddLtPN17OG+ye1/1lFZm/i+1W
8h16yoig+EH9lQPhjZx/jWuZLsU6nT+4Ies0DfyAkLW0imeY9ha0qoL9F4MwhWzKakE5nNq42l/F
Ej09I2tjMNeNOvRzqCQ9pDM1QcCNJXsrx1R7OyCiRVcktpoI2EX1cSetXe5roMDMnYf5xDBYT09r
XhxjEDJy5aluFzOPxncgdxg6Jm3qgRSnOu/+7sUs5wojUK9Ca48UZYYrMjq7f0K9MwauuLAItuvp
euE6lTy8Kj4r2GcfqjyFKe3MIw9fyNYYNBkAd+xGykTsJpCxjmJzTmyeJEMUnooG4/457xYm5vwc
ls+GX0i5d62RoDQbJ/RRVYj84oRMFT624hw18cTKdPYe8abqAstixIPAGHP8lmFVdq/TWQV9KgLe
iHTmMg+BZbJ6BuFGQfLR0V1CHVFlnitjmin0MA4KRYPuxVjVFR+oiT1ci/l1KhY7s8iJzRb1GW+q
v63r+8PNJP5cC8AQDCQuZbovMwS6/pi1XF+7f6WG8hFk8L2PmD7qbBTeWw9u7oT1BA4wMsvp2gSA
XsvxOUZSwxaJLi1qVxmt+DZvmzhmYrvuJt8w7UCztjw54j3YG3/Ty3TT7yBdJTFgR39iWKMTeFU3
fBoFtmdcw5sOA1nbF4E5Jp1KA+I/GqoOyPk8Sq2slJeWohUO+A/GL/I95oSkarERoKs5GXfqnL3Y
aoEXjIMsVqZZ9Kt2Lh2hOuBGy+d7UUr998YivQ8JTTrWyL+enjaRET5fERbFjd812Gn9mxP+lC9v
ETuIRk4w/ttq3iKN4i6LZ+cdzcRWUCYc3cmgWGy4RzI6xOspoV8wo8yp4dXHHdeqgBcyAYS5yapJ
todyxv5cpQEX2p9prNBCPtW0HAgZAnsMohT5qEjcc7hHcDhFuk/VGgcWfqcM6790eGJWcEXlhTPE
jTOE8txkrOQ9IIOeW3foJuqwpDMc1lo9dimMA6wvWlDdD6KR7+YpiqHXr9KrAdmgMYFlCNsuCkT0
A7utY3lqjl0/NNl5SEMKTG6lQ3AZu06S3VVqd1k28j7ySkZ99Lqsh2LuE+WziahzOCZol5wOnb9i
3BJvrd7jM65NfkNB8Zxt6ZtbOOm+yV1BMCW3aX8tdo9TUE4Rg1JwkLXPdgIKviny6B75EsliD4wU
o/dkKro9BhDKc5pEZDwDmQEH6F+Enij+77Xi3tS9cN0H0wXsROP0CtgzSuvd8+tj6klQ66wGyb3i
j3C+fixAmRlfKoFMggKF8ipW1qsObyLdkhbonnxdbteGLVFBgaSRAMeIOfLxcVWaBflDslBxMktB
YbiHTCcZz0nCJWXrLu8Xo9eiL7oiuhJllOtS+dPkQuK5qG8xuoT21orCu+kp9BNfA0IjugRSE4s7
LQoJ78Uj8V1twrW8bxz+G+UajE3HrpzD4mA+iLarZP/pfmAqFdkPvDnSzEL03XFKuKFxSc/9n7W9
Oy+K2cd9I2XyViG1RndGA7/GNuTDxSfvSGpz7bXo8lP1KRDtl8dc27D8wpTZjl+/4O+PiDTnpos1
2m6JtbtwETjco47sSzznekFzIUt+g4uCWPoRoOeAx/k0GgqGQ9o74zgKcagnOqTSgrkScE2SZ7H5
k8dbVZIRH8ivfGbstCw1Ljgy9/PPO/3Bb5M9X7R0/pGmH9QNzqlGabxZn8tzeoloW9WWSAryclTN
5rEcarRvjm5iNOC5K2dla7QuPxBG3VWsxz9TMT03/Ewu6UpPhXFHWCwMgryPmbawrK4nIh38ReJJ
om+Osih/exXNNn+Xhq6nYrhZXBNm0XS3zbJ0zx2imT1Z+8Hlh3ebg4OioHRP20YwUC4BeOGZNtqd
0NDadCAMi73MYiYxQ6FKQAUqudTFL6Ljjv6+AgH5ofq8bYJkIqzmqeLYFXUqDsdjFVPnIYloU0Hg
dpc5wQHQ9sAakivODIsDUm9JHxjI8uJmT0RveCZoVwH+QehTSDzpRSTw13mvDOR0FC2UjqdtZ/2j
oyhmf6lKL4vu6ruYN/LnGMV/2Cmw+4l+ug94/M1e6UowXgow17aKIFoXoadF0m5ziKIe/ohxnxeb
TBmAREtSUdJJWsTIjwO3jSsysee1OctXYmwHiQqUdMxOaYdmAp86udlMTJpGayd1MZIoakg2sEMs
eiovqD3TYs0lKOv8J9mTrHVgssjNOvA9pQ0F/KqosIwMsrewS1UDRjTEuVP5ik+ksQbVunAs/8aD
i+dnAr1pUeKUV4bvRi9v6cX/zb+swCxDZaTFkHBAT5Yg8vkzOgnhqX6vL3YLxDxs5uxgxZWimlWd
BSmPic3meODG1Vn3mLU2JkKIj6pTqNBBu6SnR35udhQJ9yIcZBZBHbKwdh2/8+d5fJPePbMPe56g
zjvzYJHfFCDU7dEymXNAmsg1RvadXvz9j+hTxpac7XRgSBhrHnVJ5EU95deJMhD6VpY+xC+Lqgpv
c1FtS57LI2nAwS4zx6XiU6b/pIxEntE5FXpEOSMB/xkZJesLqtbDfY5x2cWfjUl2uYf84cjYpGPD
vsUKIE7Gc/oHHqrhh/CjjZgVN54r1q3QitjeEfBf9RSM+qRt25GO0Dg4MiidJ4CFCxqEEEkfHiFY
E6TW/TmD6IIamE4TTfw6oc7U1/kTFHQydMoEzR3VjnbrZO7oF/3SPftCXz4kDYk3NYusfO6Cjjmi
uCP40jBfrNITpzMEZrFiUTNg2fBhnuot9/xi7MD3KRnxe7dajY0Q79m5NvcmRRlqvwcWhQtMA7Mx
Yh18bU0DvTQCVRkvDwLWTOjMC0zI2asiENjAtPQA+UqAe2bLPugELBJe2HTlF+2uBqNbgHc0VCUw
8MQo7NorbDJYh+4Zl6+8pJDsWp9CcxnT2EAonc+EFjwQ6mBqg2xRtrM/a4iUM8Mt3SO6qks7arTP
QkMH8xrIzHz8bLvF5q6RBfQAK9o8zf4UkXmAPU3OKwImnhkqoOwLy31qEQCeMeU96wrSTe8sKIcz
53oRhy2/bSUDPRaKqbOr6/WDJYfwpBynFUgru8riKucbHYky60LtFT7VuMHDhhdWrozESAj6GdO3
CbZ4TgaoVdJIj165dkhM1Il8WCoXsvP5Q0aNo5sWKCbFvMkfXrmyGg2lhOrJpHxpx9ngyba+W1SB
YbfBpOFPSM1NcGgSWxfRqkicx61C8Uq6uWGKDQ7BzN3RTJbK6iq99eqggJ2kdDcgqB1RdoHs/1ko
su6gRVeM9tsBeBvZS9x7ddipaD9mQfiuCrv00PgjPyLfMr7fEwExZjz3LLL+0WzBWiAqrD1RHQ3E
3gAIK8VfQgXofwlJXx3W6T4NRbLxdMai8KUdVWUcuOX5O61K8f1F53Vc+fLZLF1em+vfB8JXRpxV
6CkbZYJnqFnSwQvIe9GbJ8F+2Trl3lPc1YogR3GsHg4Ms0+/qjGEv5vCEeNXbZr77xPZ3dFNZZPQ
o6i1GRu/nhjTLGHuLLN+nQAVVgeISaz6P5QHflIETxKrO5JDWosoCFwFY5f2R9a7fSvc7sVq71RW
FRh3F9g/BNAA8xRr19E7taW1OZEP/ODzmsb5aik7rfzTd+89RYcEJqph4eWgMYanUEm8KujHEaUA
dOvFXBvGghwnuc9z/LUwXtk/N2ysKvzaR2nvgaWcKtypCOuYfnFqsKohnPz/nBTe5kMdppvFnMxa
J0Z4TVULyiB2DOejz1XJvqJDC3ZylnwyJ0cWUW2k4zgPbh3vLvNV2k6/rKqCricC41LglR+FLKps
/R95DYcWsYl+EcX2r+k4nyawR0AFqNbqsB/yNs4Uqgq2EV8Jtc2ZFJOc/35+HFxgER8cZmvS+wcN
/Wus1+iNIU+4IIxOrV2MiUxgzOZwfHKpGMqA3zWImfKPsPb4LI9r+IanYXPjHJ1ksTdwOY9ZSArO
/MwsGEo3Z6SNlWwT5R3TxIBwbmsL6X7yn3aZHFsx06OVbX/pqiGJRET3bw3CG6w7bnhmPe4//i82
WWfqMcWC8BhoRxce1O5IgR88jugoa/sUxExSx20nzNROsv4Xi51J+4MPTPSDaNq7Hk/DBg74Ckfl
0e8WPPBUGAmFrehWQ3+GljIiJwKEYyzxT4nifJBl/u8AmO7osY/V3TUxW1mztdR9e39gqNFBSWTW
chrMBEB7QwcBePQN0NM1N6KiHWwLQ36bRdaDbux/7PcBdgvdSV3sHkWFCoeOOgGzWhJo4OEX+FH0
Rh75sKBr4c5CgUajiEfZrTr09MtieK+vIntcIMgaQzTB1bDdhJrYUwGMynKTtk4h/EHh7/QaHJcp
OcH4noQEZ6Ui8PwGYgVeQ3BbzHNNrda8ayJe3FojTFf0MAJIZU6GpqdIi2Zv3799gzp60oBK0cJi
Nuc0a6MyDgxpIdVR5VKat4r8P9KSiikY1BsAED9ysiB1uVZHpYz2nbRMNs/N7KDnicmjVK/SGhK2
X7EtGtYhZNWvWPDaQNETOSQsnrX/xtM5bEh5yfcPvDrWOhJ70JteomgAUs0DFmG3aii353ZJhIZk
cnHoXJtukid/p0JvBnyVRiUWW6k7vMowabzO9XHUaQTviMLaBnC+/sGU4uyK5VlQjy3JTF7qlEoG
kTTkCqKVQAEYkEuMbXYSFb6/yNZn7Sk8Jul4l4FgXY/zsnu9srNpQ8epvmsKTi6JUmRhAqQ4Efh0
ZllM6rOUvX58Xnj0csCih9jj5jIg2VCK5e0YCJPC8nJFG/AYMDGqSh7eKCEEiqlhunaUFtbnua5K
vQ+ifhh4yF+wypwaNgQJMk7jAMAkYWsvhaqEud9bIRoqlxv4CG1peRgVTyGmLTzJ6vxtsHqC6Z5v
D7NDSbWnKGlgKkuqC+byUDGRWoVYF6fbMuFJFMHcS7eUmxWmTIwTsmmhjbbIhdE1LXLAlxPzp/He
JvOP+pwUs1Dl4X8wqnfTyB6Og5ZM0GORX+N/szDHyRE79nZoD4bicwD6jHp6Du8EJK6cKLm4c6ld
rvMBr/VOH05LAYkWdfhcOmB3FGfNfJYHORnSg8tbolY5idjpRjPMUUliSHPHXNqpKDWdn8i4rkzP
1+drsZdu+/ad1KlzuFRAthZmOMDnvBI8myuPFNVWLkcVaJYFNEu1UWv/ds8DRvOVRFIIThnAbifd
vPPRUnD+Fs1ZZ2VmLknSYsCgTuTyPMvcvXgN2Q9Zm4rYIo2c8OtMwkKOXZnrjzJaPbxqqztX0T6+
0y1u4CPhvyxtrZgMJbnKDjIkvCS+XZuh4CqTy2jAqF0rIVSCRbOeYzWyRSKmg7LUwa5d50hvdpSv
1j+UH1k/XeTYF7X+vP8xeic5B1EyIuB0Uc9x0jmOcJGPrUAjxKFuJUrthQXhJCw+Gwaa3qMwWPC4
O1cJoxO7PY+FlJ1H/5Rkfvs0YmUVfuzmnYkU/oJU2+7+qCvqwuK429nspLxaw723kPGCEmfFMMRQ
jF5QpiAuzNekdk9FPfVOmrzhi5oIvJlPgpyRKvGodLhO7Qgx2aHhZdXB+c//77KFKOz09ouwePyZ
EIOIFTUtg3a47D2JyVPbhNLr23UxmOpC42LTjk+8Hvlj+bq/TFIG0MF0kTGa3osqpGx0Wk+7ciTK
PJci3MKO19Nv+FlbEPiAuiqvgZG40fYcwSetY/PUvbvGs8I53lkELWSkEK4eDkqkQ/xS5tHvHJFa
oGGxnnqNcgWxkhi+dOO52VmdL51ikh+Yj+7M5MOoDvVRRF8hHbcPuXGjBEKtirQbEojOe9PY9h21
VdZ4/mvSqfye8LkfRTxBUEtCcOhNQmH+n6BjJJXuSoMLfAo4lDQxrdBEvYxkc22Nm0KBmq5dHGqm
L7gI3gZa8YUZaTOuTej15R5B/RE7V5dNKF6Tf89wFY4kwzGCboHBG02brzv62hXj3Py6veLTdMDG
O3waqVPIy3OQnXJIwe16MLyl/W3XhbFb/MMVwOjn5ym88w+lAElZn5DqhlwNnb+bhf5z6cif9TgD
y5cH6KbHamkNzgocpkp8S9+ZrUls6caZW4EWM+ZW4qglXnKM+QoQdOpFRXWeoQ3DkOKkTeP9mYf3
T//LkcOgLmO0GYsVoNFglor1VpySombT/FTpMK9Wz2WX4q44RclTzwfSIlTI0OL9zL1L9idDhE3s
agLrofHjfK65KIKXVFzRoi+0EtdSVvJBjZ97QtiYN07Z/CPo7wG2veM8YrGKT6XPURbJsfcZmmNO
SCCNAbYSoCBEisgpKf7VigB2iddLXCMKGWBvJqbWCN+NiGM5HXJMESGMtdMgObxR1e8reO+LL+gK
DmvjpZuRZ4tSn7dSCmHKA81EVPDSprCSMI0N9/qe3mAR4kWB4giKkOr66EKxNXuUq9dKD1scR9bS
iLxY/zP9i97niXXnEe9PRijhnWt8ccP8Fkf2M8mvJY+wquQsUGykjGlC6box4VXImw77FSEVKd5U
pvVjt87mIVG68Bi8HmSjbT3WgCa06ppZDNMNUM9K0TZXfumJsSO6XEpXN/Zrzm5fm2rkuLH0yRQH
ibtB5sevqG4yrkso8Pw7etmEVeD/8qdju0XsM5S2Oz4gcu4rTDSiqj3kLJjxykwPMIjy156xgmn4
ssnVssRKVyuxkY+ZG5Hc9XS85JGNqBx/XUtxZWDs9U/ZSxeWR94/FYxBiLXFjhD781WsZ06Jgjqo
EutnrJ87PKL9ZCjIA828LtVi7D/h5E0pH676hmwq1VQHPqbZQb/rLbRatuRqptMHJjj/Pvd74Ivh
y7/ul/KB7SOSwmzFHRqHzfgt/oL7G9ZYt7VpREZ2g+iD3n/MreniTbeZ/YFeLDR19GnBRnz0xSF2
4HyHRNa0IA3V/zRrzPMfnr7DFhNkAEghrmxzidyLFo46Hm+tTUV9bnyiX/NAvJTLzfLa8Fgj2LQx
T7xxXQw43ah6qU32wi0E1sPQc6QZx73vlgAXBrV7iyf/n7zjjRrUSxD57msO9SwDsdLRWnRA5HHF
DbT+hqBM0Rv1PWRO+nO+PsBW9PwNKMWH9NMTQ8oQAwGtkanzcX7zHustxby9ZAp5XxWAPYTGpv69
OokVeNUKVRXwQgQs20Zhz6agm7Q6NDYkt2KzeputRkyOh64I9sUHyxbl3O+OL2xz2e0N0sg3t+C+
tJr3g7XOlZ0pxDAxb6UBf7wJB6aOyL7hpBSlZurhqonlH4bwjj+ad62Q+CmRSmyeb32pQCTqhCL3
2eIpwwVN7CMH89egng9U+IOEXSDwEGAACXV5WwKjT91Z1/aywkqmi0SJDNBVLT0vWfOVDxMFJMXs
xcEQOQshrjhRP9fNYGvXjUo31mfIhKJVFNi1QQ8IJNP/y2gBvXfWUfLeu85ZucmHgZ0pI37A9V+m
iJXZLOvHJKxAfI4nNbPTR72v95UFmJEXtXBNc1fdNvHsiNj9tpmQKPLTbPXYNiGLTwHcXk2rqq+L
h1G+iwLQ86YOky1nmARMwZQLzqC4341/+hVyGkfpp67mzd9H3+k6AcD67NaSXrlyLpDRfvGEDHrz
8k/iMwlkKmZJAe3Znx0LU8Lq3SH3Ltqe+RJeQ+FljocuQBPs3EQ6U4aEOJicQi9FDULGI/ppxICz
tk8SgQghnd6HvqOlZx7Gt18fCsBuluKCtw7ZS6PY9JlxYDZlB6XmM2E7qZSoXsa6WUSd8dcr1SiK
E9FWCqXRnD4+VUZkYzJ7MuQ3igs01B3OfR8Y66wt8JWb3/YimOodRZlR7IoRq+GFbZc6lvMscW0f
3uyih9WA2XVqbV0ocVbpW0wiwSFAow4sMaUcob3xKx7WuVydQFXkywHXMOttE2yAiXU2aixZdBrD
cmW4zNVgYCvADpMkARux9OTRuycclockGCitxgZtyCmrD0Ardv32qE36kRMX4rCQEmKaytgH6d5v
GQOO8LJWUINcTBmHmQjXl0s2ePKcwZZw9ULPX4vEKpONj7SkZSY6c/Y9+MHhHAsS9XrzGFtFx3D8
MVhBNN6/q5/fKLR29jmM88RwlCiOFNe6/RF+oi7y1tNVufu/xZjAPtLLWce8SJMeK+s09VbIpJZM
Fa78pnyOrOByqwx7PcNlt+VCL/FDxLzB0j+CjBKzBbe4yrWSPieAcnD2O4VzCP6XqmfG4LhEp+TI
/ONHUTgWzIM9ykFn7lOJzYtqdOSOOTe/jP63sSmBIaQw1cszSmVI5Z4uqpBc5jH9wLqz50t/eeIM
btrTai4yscVsT98IW1ktVrcTZtwjmQ46sqJKaCYuFSr6Cstf7G2xsPTEldhunhMoERs56jn/Aj9h
bL7+EyFkQ2LaljWp68a7I41UMUNIdOltsIv18bs36CknTfmvewtfw9BNTfoNaNFJRWCRf0WMPKES
lU/o6d0HW/CRWcNAEz1YnapU2/udot++3PyY6AkFf6DcyGRkO0newpdaeTN4E+ogwSDW9pyEdk+a
DeiJPZSSZhTdobMy5mO9yKgc8cB47TC/biCPu47N0lANN0Vzr80AP3DkH5CqQInsOr1Eq2giC2I3
8ZusYi/H5nuxQModOG6DjimWzSu8WGnGAXb6Nlaovq5jzABr2WmZo/poHDQsfQPfHmhV64WdeeLM
hLyjBTPf0nUVTT4FIjHbJVwT5tbHw5KSWdRV0hJfJ7991jiKNYrUkm0pwtm/qcfL/5mOETCLhXDM
76YbBRsvUF/7MRQHhAUdXUdfot67NjVTaHRIxSAM8NoecTrmA5J5ThPQ2jppo3dksGC1m7gyyQmY
/XAc39U1jegp31Re2TI/Yi5lwTuGEpDqQ/Dy9VExRi34WRRfV/VMjrLF5uWvLm7cBve5VPX93WlA
tRv+9RR2Z+PBY4oGvNl9KJ+ox4KlC0M+Vot2GoYoPfOvmIPBoLa0L+DQjChpwP22CjsYPLSpXy6H
+njG10Ddx/6ywxnq0EN+hkDvjdqK8gHg8OFKbk1MEPsH62IIUnAWU7W6uColWOi4KfOG3uCyf90A
dU75bRin6qh2SDuJoBUSZ2nBlTdy80YeuF32sw+t8iserABk5TKNDmtODiQ6QbyOgX5a19n/wtfX
66yNV51kZN9tBOHLRrZXaduWJmqbtVitQdF65D/wI4cVysxtXUccumM/dm+F1Or2Pgt7p53youdo
V1ZDIgmYtsikf03M/hkKhjHk/9UnnzAvS2d33emHdlgn2EO0RSQZq9W3W4btPWbdN0FFT+v9QWby
YC4Ywf4Ju7LEbqlS5xo17jVzCf/4pCTzL+ReQhPZ0fBXv+Wm63SG2n+jJHSNK/8UbR09d/EY7ckv
FPBu26zi7ftiXWScwt3HAauLd05FYLa/mS+egaWAdOHoIQjtAryYK2HImKaVfRniVI3VvsLYx0Ug
nzhpP34sV+pLpNm3PFfb9Ro1DiqtHvcpIH9vPnjZ1Z1AaZUB0NEYcUhrkkagJRF4kTMGC/S/M6i5
iYweQkeFMK+WCAK0lnG4x9wknDRKl8DaBNV6Web+LElqdT03uKuRp0lY2Luho1S4SakbWZ8w2BYJ
2qwwzfVZy3wRoRf1FKLIYxm+zzqX+p6CSKmVGon4mA1u8XdTLrU37HY1b6MOa65mm2dj8CNSzZI4
cbU8cjhT2QeL1y4YaBXJ7WQoXSfs+xomm1KrJ9yOG565xCIXi6Ly+/P6IQqyWFzVD58GQVbn76vx
Id/AB591rjtnwmaEpk0aalZzmHbJAkePaoOZLYou1aSchcnIWhLNyDQOQ7mlnXnCrEZcaDICBS/S
hvH2P4N4rr0ihSk1WC+3v8hTYMp7NIxGYD1kpWoEoB+NqNcVY8JS6EnmHIdI8XniB9AxAKb8uY+4
HeHs+RUEDkwAV8mVCJ02i4H0YEpVscbF6UtJhThYfOI5ACEGFQjN+kmTebU3se+DIpWQJzL2z7kb
uXfHvP0/mlK+2AmK3SGYIzkx4UPGR76yOsGbmL1cL3yijyXM5m/KnamuwhaQh16rn183+ufeOmm6
MtGmXmW+g4EGCcQ38tkGx45rmGiemTnX8Evz+1AHc4dcY0Blzheao+rG2UpdtVL4UeKSMAseAkVT
T10eli4Lfy/TFhQT9Owj+BR7FSgkCSI3kYXaFJ/rbFZDycZXmeUXxhrUJEUMcVrjXIXHk72PzoN3
doCT8X3nLBg2W3/w6EQBVx15pAYpnITQV/Oo/KVCtM6GhxCy4M5up4g7I8PD66kDKdQq81Zb2WAr
yPeFxR3pvREEpqTrxYciTLXSF1IELvogzJ15EJauLFHvlJXLkBBgyj8zpcetyYKI9xYhpKVwyLrw
uN0p9Xbz6CN3UkJyEbDvFcq80Zfztnv0qvdIesKpa4hdf9Ef/qJ46Ss1eJLJiCu2XvPxSfiJ7FcB
ceUdgsmnU0Zrhm0S8f06gZftFOusqIqb/yKUfgFdJqBAXCiMkfYJ4yBBwQwl96UXtBItuQhcNYla
X+U37XwxeBxYYkNVDyMfgccuOHUO3AVlKkFHl8ukRE+pvDFKRRlgknqxcxHKJkd70Nhz9H0XmhKM
5836PXssy5cHpOq24Dr6C0bTUAehL9QbOo9Q/HqAqOvBa3MWQDSBp+jTKplSjFHE3OTVEUo3l9JB
BIsyv2BdYbpWMncya5sTpd+AqCvkC6gy79xDYWYqBsUSzFo2kt6q58xnYiXc6Cha7Lv6zlqziXVu
i4FqkVWj7Oda0AYCnCa57ntSfVfcr0KZbZ23FsvGCu//BWiRPBzBlFwft6ECNMii0OxNdfeRz7P+
1IRnQ/Z6g02m7uxhh9UxcU2yMeopvzG4yUCRviviA2i/4CHQ4lV25iDtKf97nI7+R0MItDektoth
qffpsTED8Or6zEgnorXf8CmHdcQMrCCl0HmK4jqaXJXbL2ACWEF4LHGaoobMhaKbob67BrEJ/uW7
Pfen7oepwmFZtC4SUSDzU3aoLeptgoqnEgrlb0fAb1PD2R51/QUwLiNeaIVQIpcSMycVF6xHIF8M
yHkCfE+1dJafxmDPLlahwVV3QsV43p1zPY4gaMQZn/iTvgKhOXCCE9NpUjtBtvwfKVEDuFDeDeET
H3/ZdpofPH4vW/Tjs5PbMkrYlUzD9bjAEYhRfuapZLQEpfCRFd0C/UJ71LM5OXYVd5YM26ibVukl
l8mYf+w8HodU++k1Dx2vcs3aRKWHZIcLF1B3OBynDL9eWPwzO5vF9fqG5iGkSMKZhflx0d1fmcG6
qRaTrza2Jf3pp3H3/1iUkRJg6l72KHpS1ZKN7q4J9s0WxMu9G/qqZZ8+8z9sMfJ9P25CkUsVXeLp
DfaWG9Ww3id6RMbT72RVwdJ2Z7Zn57jvM2z9bzlolCnCRP4XKcPeD0a75BkhM2SJC0SfgqxdXcvj
uOgveSGu+ufKkx1Jtiu/KRczdwF77utVXLSuthPYCilnPj51PUEuOINT0TjfMEwOdksZKLWWUg+5
Yk4dgKh9CVaoGHAdRVDJdPeJdGnGvBqh8dUgR0pS96yNKr15mvElU83tycQ+14ydvRLX0VfICUVL
p5ZPVOK+EUYr7iRsNG/8DP5hmyetpHLboPDXKu3TanREQLfjkVmdTE7RVxEkxeQzyarIOSL+/uck
98J0Wf4KMBNuYHVSU5BffQwtNovPArxe4Ax2ItFNMzknXchELJQfU5jKy7wX1K8J7YNWw1MpDbQP
5dhMqIgGxkOWViIJTB5zHy6EwtCg1HEt4FMYCapRLO34lblRASOm7rsdV3+GB7/uZuIe7mKv9RLj
AE5vLZzRNH1gsW9BPnKNlE6f6zSunju7qBMX6YqazAMC27PAhRC35i6g8oDJAa0mtUAqprR7sbnP
cIGJYdrbFYXxDViMpb+418dRm6W6pUNpO6MvDBp3yZ+sgRmN/gpECwsR1Ewa1N82qRl0F0F5BZX4
XdnttBAp2gNKjWUAAAsufznO/wKkx7TtwXdVDHsvB+oY51pjnGWEKEhZuFQDBZdgUeSFC/tRONHm
YjW63pIZJbY7AV6asLaDkK2xEqXbafX0T+nByWA1+SaiqaadGyjoXho3t7o6nQUpd4IiTrK2ZGir
8cc6FYgIfVOoVTirtKA0lSFrDcNOCDHMUxyLmwgg4OWsiUwd20UIzZWbZNBeFXtx6GAO4yIa6F6k
peOODlyJcgoXXkp9G6hefdm9ApRiUgDrgEy3pVS0zCl7uxbyYHBulEUTFHX3XM9j0K1+xoFCUm5F
j6LtaXisnUt2iAW6jwqPWzmK8Mzg1YOw1ADszT47dQknFwNLDPXOzvk+X3vyOmhR/QEWFbHvnBBn
CybwAXlS7BVKD0GygGO8hDUr11KvcqNyR9c90eKokiMvSPewGlXkV65hODsdKCxPHSS8TlOsQ28N
7Qw94mIo4MKt99ooser7+KiDi7ctkr45QelY8ai+FkYINMgJV/kbZlms+4LnBX27geWzh3dzE0ME
FFA1+IKLLizaG4xTjDqHsHax0b28zsDvWsz7ineLxExNQCrETKDR1aMP5VxLETFTAAudnT+cB5/L
nlE2f/GNbS/Nj5TN8qvDBDeBybEhNDTkUMSKijBVE9n0h3jF0qiKuQoin1U2kUakpg/lJFuFvJ95
xWAuYGR0nRFZ2fVNwMW/V/M1+Hny/y2G/6v+vQ0CQ+a/vRUW4Jc4wtyaGPfViV40WX0CuR/vpFLG
rB9bZOw76Pcbh0vgJ4ECRXzbRtwPYJSwuIMtOMB6KRwXcG/XDou811T4XtV1khY4Y6CMGkw34a0y
xlYZG8nfG5ltpHQbYJAAfhOzu5wjsiDE6/BDERjTuCL9lQABt4aRWCfntZS10Hu3PLaeoeQZp87w
krFCJ6F6Q+DZ8sJuw7VbSmK7rj5CyNfQDoG1baR1TEz79paBUOqX12P0R/QN83UoDYSrg2Ycpg4n
SdR8ZDkYIag46EU7oIaKceLx4021NK+Fycea2M+3Tt+h4bLgyc62azDg5BFHHsAVjWL0sUl+s7Bj
XXskqzSrnwvH29mYczezaR+6fqSAKt6tHO8KXotvWzNC09nVFYzkJ7L+wor5pzyhOx9NKF1afYoR
9Mbj7e1dqr7UjOBYbcMIXATTBGL55gjOgCO+74ycQGtGMkUQjBzBZ30Da9AxZzBURh/tYI81NFAy
kpoQAo1ZAQ7GQA7kSnOV3OUfOG4lJvWcEERaUOm3K5kyuaIyDAL1XrCHHBBr7zEMvrIWJdTizmM0
JVIBJGVdhJmORs2t8z4ernD5FWumcFPl3HSxa6E/9AmB6vbubTytQLIWZDgWBaNrmI5dekofAPvh
UBNMQWhzhkYfpBdf4/PNuZVAn04Sr4Xnz4mmuKSNP/ieD/TnjP5q9/fx4re0q1OzTUZujms8Vouv
ILHGvQTcAagaSjAv7H5qlJjw1x+73v3eh1r/M9Irvt7buo+f6bAPF+FyIRiEa7VJnAEzk3+pYLK+
vuwvKOYfAbFhyJGyJjYNvPQ6Hu4EKOEUTLR4F4pSiUT6M+GP1ESYLsCzk8xFCm0OXM7V8MHhSatw
FsmanQGVtYVz1DPCcOjf+zYe3pHiOe+z50RxLKqPL39832hZESc2vzngGpayG2qFrLIcKUACaMVt
JLVNyzTLq3V360rknUVCn7ToIdWM2ylCAW+3jJUR4tnzR4fwu0m9Xw25q11V9U3gV0KiGWWDXWSK
+YeohQ7JKyM13bS9O8DDvDil2z6hCuA1JSJ6S8DMT4XcIkvcgv+tYaq8SLYDOcU8JvbY3hdStaZw
yIeZ7yNfq1XlGUwfHWkubbkrnGb8aPAYiFD+3sUQpyZcwrzYxQgXjCxXMbkTEOIiMzTa38/6Lu5v
nDDdElnYWFmXF14Qzmqm+VfX71qBV+Bk3goke8WDJ7A5bsA5chstP4M3oehJCKnzFF19lFehAScu
zYa6G04pwliNDA8m+ZBLjC784DphqXgxe6yaS8Zhmy48v44bcCHc0fWn/meqzzv0YAof1Y62oMz7
A1q7u81Suc/VbSXynI+iWH4DAaJIeqquRCCm03+aq9epLCW8TnEi0nT0nwYrKA7W6CtPjadsHnIv
xAdwlRRC3GyGa/nAsFUX8mDJ2mDbYVApbGj/+dHJOspsXSwiw5gsO3t38nwyAuuf5krj2V8ViyHw
0OL2NogrLbBFqTdLMBBW3EvduhasG4gsMj06eKQamwrQMT7+FmHHW/eTB+ry9bQmn2zGhtBvNhky
2DVMbM1xP8E0OF6GzrzPhmNEbxHhfjZ18IzjuCyqZmV+1m1kiS8bZ9exxwwYNISvyB/q920EtR11
XcHY6gZTuRrnwpXpnd6aEKOcZK5N2Y0kXsZRo5SoH8GSHWsN7DGEpKGPZV1ZKyAB6oOpxI0fNxwN
h8sj9hOYxzhf2ccBXs0f23SDXZtbZBHtVsJsH5M8eOnCXSWW1L/lcxzzvncX7ZWy58elPnaKfbIF
okP6AiGMOOA6NW0VG2lORd4qwQtjKRP+MLoershcH96TJ97c9TAxGV1zjENexTZtZGSEm310P5jr
IHJ1nh8nuSn5j7QjRaI82HkAqUp20W2Cum+1krtPPKXJygFnDt1F6cYZHGtytTxo1bvfaanQBn84
EQ2elxH7rQfF2LolXorVtPyGnDcrDzCevw61VBEbL52aufuwcHLGgEoyIbITtBFFZSfKYK5uTF5a
UlJVkn5s5178MpuDot6oMZLzFlbU3teqKOopFDlLxmfVNxlc0ISy5efGDlZRRaBdlxmsmUKE0mYI
xj479pf1DH/tOlzGcrlCqGqt8H+DHwNyU1okW/r5kqgn9jv+w4qCuHXCP1cPap7tDIL+cKYrTTUH
95qKwWaV2dFsvm+NQ0LxnjHCrfasWd80druSoved419VEXQ7GAP/NOhJatInsJuMTgndOQAevfsA
tr+jdXjT1EAYqe6M/dE4/tbR7DZi305FLY59D9TPeXMuFJ31vNMYOlV3l475Otnkia/PNLzTo7iX
ThFWFlzjBNPTEZq6bEKqo4azyv8GI92M282gFQq+kgH26qun1Q9f4z+qlVPmrgh4lRW/+V4hZv1E
zdknBauQ/GL4tMirOTxN9SfxI6ylcW2yvXQYZJEjEwheT9NzDsjishT2aPXNfA+A+g+8Yf3JYAXO
FY0gwD3FhRt05i/1vY+iRhNmp+Jzq3lhslUKN/SmNBnUwHlOXauHRlCt69UXa01YqFu0JO/P3lLV
/SK8FtQonYAmpUNMmAdDas7cR5qTYCR66BFbWQgOOxX3n4I4izt0ypAgra+IE+M00w+2WlXISG4o
G8IU2NQAAAtd6eS55WA/ROHk9u05RWhKhC21xKcp66FK1lq/zI+61/eKfhBGvpcKpPpnGBcrjwbC
jnKmZgm14+0AFUYRuXm6Mg7aiQFUlaQ/fdei187tT8JMLKZmpDIn7hEkR5VhL5yftCwy0TFJkGTc
1bWMWzAVNNcnykzK2kamvaFeGi1Qw3AW1YhJlsxA6TvFw17OG0YLxgBF/+9SPHh8ZMbcIWFL2i7y
Qt8/pqU3jp1TkwSRsMgxeYn+0B3zrTTR2dJNdLYz7JlhCjQhvBnknVGHkmp7ZTgTSLuxlV43Ctgx
Fz5n2NUEz83fE686mb4yFLXK3wojG9QnnszihIfhKQWXBfi4tA1wSlumIeU9NUcrS5YliwaX1Tod
deTiJysrHLfiia3sdem3eXyGq/a//WCCF09x810GWFsxjJNti8qPhW7awJCgonp3CLdoxOi8UU1u
rHyaAYYkiv8tevyzVb15eSa8By0hsPpiQWvW6jZk5RPrwR25Xxfq/3EyFWNaCuAx1lHVVnMGyL+D
up8kZUWVLD7nGBnnl2Vbsx2pJs96ezCm9hsXdDr8+KBG0trbUft0ro33W4LvVf7kNQZdaaQCZL/b
sBKHX+cZIESwm4u+lawmNmi1QYhpcVmIDfCFiVRhvT4h6OdJ+g3X8ivbxqZqf46jmVDdtez65Bv9
ki5CEt5FaWHCet7ysFdWXn9K8wt1Y2aeyNEj08BftVR2SmAmtQWgEgWuz46PLoy0Sj316Ukiub61
c571CklY81ekmYnTUNLJO2F/KTjL/ACSALH7A+/aprGq6UDpynNrbgRIeiI+yavCCD+yMXOFPBfj
aUv7zm/YucJzKXtNoZYWHT6GdPZ4PxSZNg5x9qhlxBSZgE2PVpf6seVNqKdfZF0XEPAu5Xz3ZqWT
1jQhq/Kpz32Mc91TdBIHBBw1dvTA0PJosgF8CDmpEAhsigttWbJKNIF53qAKPoBJueFWdv7W5TuK
C5cnBlESHR4UPBcSu/YZUDdYBW1dmyDoQ36h1BoYkYbuzOUep1AK4DFu5314lvWLLSvV5nXRvraE
ZfRns85H4elB4LtdaA6Kd+ZKH4c9cdtnw/W+IiF+e+DyMVkJmsczBmvr3IMVD7+i1Y5w9dIJ8BEA
5Lz5dbeWKtSBUq1fD8f0asYLZKC5b5Q8bmI7z5n/FD+WVMCgiAKJDxKVdCSFoIadVy8qKKIJ4FfA
+KliOtGtzfO6LC6ZrkFeHJ+A8nMls+Xo4tZacDubJ+Fo7b42klwADqr3dJYPDe0v+jkxlMx23gex
jXYdFS0sM2n8iyaF7xBj42MvIEoKkQEFqnDdnUQM8iZ/lbBKO2Fr8geYHSvMAgxWZ6SUV3qHAI7x
Z8VjICBXizTe+J2yaUKWkMVV14ssrlx0F4oyo5U3DLe98bbYSUC9Gk7hn6e8hX4mm7S2Qq9eATa1
hwgF6Bc+dHDgeHHDyv4yZUVlJyiPC21sD4637KFSTPo9/vp0l27BP7LjwHsfsg08amNu0LpJXn41
Pl45zLYK7qs2ju1Nur4nTqrqck26u1Z5u/GgFf3vw4tmtWY34duSp+L8FO3ZtzblcndfME/ZjiRZ
dFHahBxyBwA3349hsbWGoajmzr73OnjdnpK0CDvjVHvgWlzWVwoFVbJ18R8R0peB1D30eRExr9EL
DFqHe5l3RKlCMLL+Y1gNGIwDHWsjBLLRoENHI/D1RpR2Bj01BO8cKn6PS3qIH7k/iMvVWvgeIqWd
qhQFBdU/LATQUL0nb2XtC+AI2UfLLltktL9eeUJ+FMaTt4yD3qwAZa0J00YF4/9nsoKKho6H7zqU
SS8rkg/23/KIXWjJVdvvjmFt4ey+OA/SVWpwMU8mGlmsNxHozo5g2gvDgY25U3cg7ePP1Ko5w2am
HERV+4e4cOCxlW4Y4XZtVOdFjdBtsh/N+zVLnvHoSeg270eNSJ9Aq1Sfg0cR7khHYUwHTor4Xzzq
3S4Bn79fC/nHssVthYYgZtEmCJzQfcOpLMptp/uLfpJENjnlWnHB95fskOuScx/E1JQlu45mi3b7
/6l4qzzconrWcO9ShPrxfhb4iATGaT0ID1Td8QJPDe6+/lM5tbF4njOSx4kdg+8L0Lztier9ZD7A
xRrNiKV5kwUZjH/jYrrUIS0Hlh7SeYaWs4/BjGC3Q5t6nvX9V9Gw8YX0LU7Zwpq22fkFc0emVKln
DdFRiK6qPesHL76sLqsJYxhPTPtRwthfUq5KPXL+dUGaxqKI8aeemTN8DQqUMYmJtYsSMJk5v3Mf
dFDOwHW3+mZJamJ/IjEWIx3h2S6kIRKvABUT+buaFjCY4S8/nQaTAPI08aMQj4zGQBvbX/jLeu5j
v3909GzK0btI7AxHujG3/XUXnS2sPRd2PLxuLhff3C1f8IlgS5MMjc1IIhSQiVoLp5rSa9Pevwe3
jDZo/yOwq8mngZPisAn8G9wxhJ3sQoHWi1YSlxnGOxnCG4y6rGuC8SoTIyQmkMsFUkdurUft0uvY
bXnWsSjDcdANwX4lc5LxhrCuvlCfp0y9cJngYDbPNslyBTccndiW55wbUoeaGlqProbUNjP/jn5y
ffcYA/T0Ot/UbZFM11IeuWgeZQj5UupcRUEuycArwgkEEU7GOTXUpcfhn9nRon//Jnn+ZTBRaFxV
Ixhr3kTgUK5qbqyHZC3vISDvgx5yoXVAWnTIDSk24Bfl8YWWxTHj51W2WOBZjOktEG7vMPpWyqLu
7sw/RRl/jAWHxp21KBq69a7DPPUgSEP1Y+ANU8sY00h2f9TVl42aG1Xhd9BrH3/30lNEUROhXln1
LajYy2S6t/6WqF4cWlGHVluwfYX2h+ZyZfIv2IWlpgvXGBiLncX5jeO/iFuIGa4+7Xa4URTKdVsx
sk/gXzBT4j12H2Ym5L+Lue3ryWl6VUmIGENdKyPxT2bpOD3ZqiAkUB238vHTIMV217NpOCtJ4dc3
BXu46mDGTGXtqHj9N+qXIlNeaXxRMIOezQJA3wO9ge00uv2jxTsOSnoDBFDK7YGFM3J9ux1HvJ1C
t+xKe8qkOsLwJNWw2YZPdUFj6M3MCrwOjyeiV/hmOiqJmzzkT9YEDOXccQ1o57vMyn6b1Hc8RCD0
qoqmK3UpNTSp5dwQjBDGSt7Y99BtG4Ymp4+V9Mgbd4BvNHpC7p3f+K6fh/dc2Zas2Cn7+wGIAFnH
veOzv9Z1lRNzNrVb46JpTcGzWdj91M4F5SCsPwNUTYxtu/pROjyMIPT/lyGJL+eMgPuPWStGMr4r
PBHSUlNVHd7kvHNyLyed8J2FnxejxsPAUgnrn0OshG6hxMVngPBTXlTrHGt2itAe5ry9uzUMzwm1
YRmdNdRAKpGCIOU/3Vfo7uApRZyyBLB7XZ+NbandjX57Doy135EgHIN8x/czfumzIHUCuL9tw7GG
2pEjRSC445MBcgT1O6Lo3Lz/JntR/uzeef1JuamMSBBX5VU/K8rk2OKAis1C5lfOwTWdCw5/bxcg
8iDCEmv20iQvJ0xhFXkSHORgrWYJVJO6NSMHm9H5Q6DoWQUo3hAlCjVXokiyamowAd3ROH13pGv2
KlxDmgJcBD5ZqUcYyl1RF8obola6CUGQ4qNlcelTe5hPg7jLLAM36SWutr1m6Ej6cd1nKwyC/j8k
IxwskMDVtCcRnZezd4vHTRykDx8cLyf2x9zwk4lPslq3FIp1AI7PCzYfS9BnDNJcOUHmt2kyN6vB
P1AoxgNszhcofvdo0KxXiE+wOtkC/GRS6WnZPoP+g2ZBnBRwdw4P3ySr5F6Rl/AjJd97wT3U6i9t
fD+nopG/ONkliw9b01zeIv2hsAQQXhxQV4UDyIWYfkM070iHRIik161mt5hCCYSnVoxqY74Z9w3W
OtsO0EQoL9Swadh+mUO2UatFOlYUjPbQPk+dmxNvxTX1Pr120v0XBNtE6QhaUKsD2WTDrvb3iZ2d
eH0C3ZZTZOCLKMinu+5MOrMuxtxsxT1FdnpZe/aa2Jqe5yE8y0KM1+FyewVMQzXMHkzBEYz/BJvy
Rl2Kde1IQqT0fksWKZbm5aVPhFa9BPwi5Aegi6Gb+O4U6WSc0j9twIxU1zZTeAlEnDmesrIfgQ5N
iqfxSmPelX7zjG6a3342jsraCcrOa7WxgxKARoS/AP2i13fObj2TyLwjnk1Wi09TnkyBsk64bs/8
VVovy2Pj+2asyPco8gbALPN/r3F3MF1zXC1zdQIkIY5r7Y0BcZ2vZwnUggPwW6TqMqoIukJ+LXkP
jAoVrCtzcOyHSS2AE8tCEHb+gzwWJqetQohxa8gmYTj2tXZU3qCmsZpz033n9yW70TbUp5P4C77a
yNCFWlBexZwsEsCKJqA23B+ujySMYNqDZ9woGbBDMyKr3FBaXjIXyHgSW6pJH73D7RoVGdxW0upu
BMCGN+2zghsQ11NpbUc/9IoKtucpIFqIbyZxDMTB6aVLzFEfcMykAAuZMzN3j7fmxhLNtOaC/f9M
DfknZYb2L1PoX9U0wntP3JB2fKUiWYzdWaNLGVw7+rDsfXa88unRJHXbx4fH/4F4UODIIRRZnYwu
ta5sd00mpi9sSUcw2c1E5kAOb4RrHfP+ldMvYSNNfMGLg0jP53IdUZyFSCBKIxTuw6jmLwUlluCH
MaZYVyIYnJxXNgAtT5iNvbGdaUOXb2FvGE0AJPOPTJjBN2YhYBGs8vBGuGO3avTMjpMcNpkwh148
8mWjRgrxMyn43v8R7HJZbBmUXHk1iZP2AaGp4Mn2Ots4dKzy2ymvEuVqwlirp+Sl++K1wMGNVyn+
PePsShZ/92faYs8h4BVhpOP/mhhTPI2e9gla2h+rSrKbVh9yN7/fmVyC71WVwI8OeZ3zN4bZYq0h
zuOZUqr8exNtgwe8TFVKnoJAszrdYKi9Lwy8w3Ft+DJVQupIMkInZPo0261kn51qbGSI1mJT04BM
cm6sXK7Na900lJmPApaA580LTUcibqm/Pq69iMhnV+BCAAQDRyuMJH2jUAnp/yFyqURlJewgWHb1
d3wkff9Gm+BfsJdxSw+S8ee+nQxPANXpJ2gNK3/ALUeb+bODHGFofBFGk1dGOYy7znOn6SvDc7TO
uEqXIEXJNXUEiGPBRCMSCkBzD87rVP+3X+gmeNiFBKyWVkJHFsPfLB21AAtubAUnQ8gwKERE03WH
jSxUGDpdEY8zRefxKNw8f3J02Iv9TRYzzXg3cCK4dfcoImdy0eWD3A62dBKugCjgbplsr787SFps
bF+2RDVegF7LyVJepqH/KyRQ/oPKMAj7ER13zp8W3yu2G/Kr1rd936a/w0qEUVaJ2Oipxv31B/7E
w+pDmTIL8kjDYOU4/4GwpkiP7YwqtvVKtYdXH+gFVnKsAWmEM0MMkzihKfIK29ZsRU2TAQ/n2Wg8
vzka08tpC65i1FgAigjWNSe8NQFYoTglDR/IVizOzjY3d5aap+ZziAS6kz2hUFdBc0I/IqOss1zv
niv1OOgZglD2BUoB9VzOFtzVyz37Ct4p7RI8qc0I73l+aHL6HyT+vf0eLCxUDLyxlXgZtiJZmXOo
C8ktpQ2rWwwBx1j/toNAG0w5TWfBJCVfMMYaAVGkz1PXoAnwF06yweDelO+09UGI9Y9rTC6nY9Gx
yu1xoOdgOnK6Gy/y+bwZuYnjQLPkONcD5xpb9CeNo2oMTM0jO0Si0b01JFKIMgSD/Eg+0lSRmOxU
bjDHDEXuav83d6KEfMaEALKmjknSFSIHyvDnzMdgdIr8zZ41OmSILfiLP62AIJBlpu0VwSIkaOpy
2c7LBjIw3XOEHuWlo5RyVpDI7w3WjAzy9bGavyxOXxLFJyvf/LbiNsfwbyLIlfH2QIGhFcvVVTdp
op+l2+vFiAuelTP41Yz0uFQprAHF1kullQIlXxEHNPtzxlI/7WlhR9ICminmpAtCtSy6fYzqKT9c
iD+OGXbxHvfx5l+Yc2M2zFlB1gUavLx/jb8eduwQHZYorMJS+d4/eAr0zoXuSDcqzY+E379RJQ0e
5EkB7gZnBPbpbiAs9wQL3l8ep4GeD3xfEQTb1Z96vu1iM84TaFWH3Z2trcah+eyI7cC0ZVcZFItp
o9nwuK2bPSCwf/gu3DT8bWO6mt0CZ+pbZPoE5SABp5ApyktzPiQUBtXmvfg192+hhEr5bjHu+rny
acpWc6ZiQnCjqdutP9wTk6+EhMLvb+SOinpHFi4rZXG23jF2QjwhWKkarLsjYE7IX87IMQGGVPqf
reeVp4o03FJjzJiu4yVDieBjY3EHaU7NhTMmtRPQ5TDl9YLASuE7qYylfdV7kROXlS5Xin97bvsP
i9FV25QQluivostmouNNqJIytjBBl+HpUaKtRPfyJg6AlEnQAJ3IVP11E6riCcbFMilYUOs0BSOJ
xkd90h86kP7zlbl4ISvc64ezEy4gOGQ7Jv7omn9rrIzFPsYBxtXF5bNNRftHupaB9aDEL7+YEzX9
89Kv1qn6+kBAGW+Spa4YHX1FxjXgP1f6hWZs9jNkukWS5AAkX9GYOArfiKJRFznZuOwgat5gXFix
fP0EI+8msSx/DcE4ocNjbaQbv6a2yz/23YxQBNof4Mf1FUz9IO+fMuVMy1CqLIyjojEuQ+bUQLNi
2TZfZqgaDpfVxOL0d3VPA0LiFCmTEaXNpH2W1gPwP+Tgx4aSFHH++HnuIoFaDdzXGq4xwq0kODUR
yTmBgAvGhtL2IcwiQRLaky44zFLlFA1hQamA0Xu73FTClec3OMCzt+198+rlb2whswM1WDqkvCxR
a+9S7IXOjN09a6WegFFiXQI0QIWBrQuVxabtL5GKWdtksPhH/Vs1BNQEBYDCft+0TkRbFn2wmnnW
ZUHwR6cl0gZnI/cbZOMls5FgFktHeql6/OeVIdQlTTpiARXxUgwqPtWlWC82FVA+0MU5Hhy3MsMq
DsQeGvWn37tYSEswT+EbD4+ZXqbPbC/0r2iA5mVbdEyW9MZB2QVl3emWix7AmuHH+LAm22w2hg4s
lOwkJYURrmW2D2H2TMaS1+9aaib74rBs+AM7B3/qoLSphNximQrSkoeJ7TxboHOi8B3EjkiDDtYL
a2dfHoXpdHnxehrXLpxAVK8bc+aW1ChNkqaKl9HBKlELqg0Udi9uNDJlDxuG6LuImeZX5MM78YId
XGo66nlGTuYEhAGA8pwtZB9qKW594imJ7ioEEJxvQI23gYiPR6MrLAJkp/u4ApRxUYKQ6nXExe2e
GEMQ7JJ0/FTe56LWcKOTLGgxklN/nwJepcNCLUQIw0rEki9o9km7czdu5yN61z3dWyII9Cqr2bll
zpF+DFNfW0ciDu1sCI0W8tMXCPc1fV2cXhY6o3SSFHLu6ERMRSIe/2fSvZCBqAW7eETxOB7nWYa5
8gBCtxJsKQh0fUjScU7XU/zgs4Ul/CxOsqyGwPj3Kzo52V3qFkG84jvQnQ5IOe8tc4wOv6eZ4RtS
rH4j1muHEBWNtF3RlcJb5BSriNv8p8yIOrx0gtspQHvwhsrKssPZZAHjt/9eoPIBjfQlDv5P4qS+
db7hApwCLYp+a1gLEUw/afNVKadmlH6owTfRDt624rrkzX0lvQlKYyqJel7uNEH3fEMrskPp1p/8
Q+PZz0paY4dMNHBA1FyTbV82eD0/GMwREA6FJCvRKmfXrzEFOb/tacPAGaeTOyAzVzAigpnWkefL
PVDA8pQ7Cu2jT9E0CzbBE2rHrJYKS69GSYCdUnLIBihFsutEClE+soOFAbM6V/mdCxA0oFISoFuf
jQCZOnsyfiEa6VCpI6sqmOI6eFRkZLwVln9+TYKk+JniiUQsIkD/ZrW0BvSnewd5KTgX6XEOY/yJ
uLqvZa6MDoDZCo5Qey8XkhMJH9N/w7ijN+Esy1FOVNzUxI3ZtshitON/MizCt8A8oVfKEgW+xc5X
La52b5+RFWzqwTE2nm6TeQLltLrdHpYeqt2kztBsO1/Ry1DL9fncYrtnUzzyVJROq5L6zWDEvAKE
taSs8dL23UoYF+npv+x7seFjlg0knuLvGzuzNw3bQ4HSpT9DGh7c0NmPdDqhAeLBWoqIX9kteEQF
EGXGniaGwm85nRBsOUU1WqU7VHJ05WTlKzJcCQsbvNM3mGMsmOsKxp89ehpDkaceLXIkjmF/NwMz
08bJT2oM8Jxyr2oxJQdntyJLcRN2N4OOGDdnWxsALO/2ZLBGlQNHPS0r0SWRCoEu73IbVWKFFTBj
X+DoZjjLoKAEcIn9vlMVOvwohG6QjnUfuq4w0Doj3IzmSXlwDTpPNXwsxJsCQrAd26RZ5AJRvnTb
RyAw4XJb4wxgP/00+dQpX0sbQEQMsHGklmqQZgBrtCZMp7fhbVgmwsB1EwuTQOYgXw9jDCXrnBMU
Y0wokktqrXC5qUxHOWkJSg6lrEdPJSH6skH8FuEIzQjeWWgKLAgvvXpuVBnm56f2RwverUtfu9Ir
/OlAu0RsKxu1OVUK1UBpU5UELCEqQyYbFntDkA45BaP7zJEQ+svjWXtWOQhb61Kp8pw1c1i+orrT
G7vQm9AmcoJnntW7W7oNPTFpFF5Xrj5gR3YcBQWzpd9ErrUW+4rd/ZmPGV8+GWnZy8PjedS+RxHg
TsyXWJpYuAAEbeRSQOTR8jp3CyQRn9k0901WWK6/LQa3bgs8f7xisGt0AUKd6n2w6oF5D5spoOuh
eRcBwXsU7eVDkjdnYjlZtg56QcU6AdLK/x18akH77/SkMmR8BTGWxzsnha4AjqbZhUNvyeWW0zqQ
z7BA1msKZ8yL2MsKi5i/bUFeC3qvDttYCTAtIiYLs3FyA0rISK0XOwLnBIF10UcBWDViAUaXEqG7
p6WHHaXVqt6cmtXCqylduww2R386i2ydd0uZi2r9+oWtCZtKfW1Q9FKnQAs4IRQNLeGNyBZHPO1A
sDcEfQ1K/o1fVrI5UE8+QhQ0wXOnA5Am0nNK8VuwLBOIfh2advFkrxX7nTdsHNOSIKclgUAPhUXH
6qlM+SDj1sLC1/aWWdGOQ2rARzvbDC+Wa/U2cxKOWZML3/wiQ+SXvXCe5jPVlxBRCXFMKy8bAyEL
2uK/F+21gBxPByxKWVmSLz8HpwsIBfyLk5+kWCW6rMS+JCmU54gixG6k+tQu4ryxMHHF5yinQxym
q2zddx1BFhcyaXt0jgv+bIOpi3anarKnMKEFRkNr6Nh8deXZKOuapxUUwsT2Wx+HGvjSYNYsHQXm
SjThEMbamciCcXa9eNfjrZQDRb8TpaWEY9HgGxVXiIwxGqGF4YhqLm9kOp7gJsHq9Yq1hyM7X7YY
nfvlgXUhHT4aW6b9RSRINdAHOZkvCnt1JG3moSx1/abijlLJzQHKhbdX+2aFof5Gpqayj6062Pq3
zW2igAZkclCavmRVj6TUfTzW3k2YlgtMYvCPXeDJT5rud/wIoH5q5oYp0ctgCwDsaorpHdkVF2o/
s1ODfViNr7pa62/KH16iFRJxWMU3LyraLTIUaEKUMVe7SfVsf9VwtCef0AcewTRRsEUomCEO1EbP
SVDPqW356TlsLD1fhWkPo4EYB1wI6oebZ/8HSu4pItQEvq6SRFZogbd1CAI/0giWmXPh8FkEVYo1
J2xrAjdPhbEeSvqaRkTRvSneIdhhup9Mj7myzJT9Z1jFgyTaHkEr9pPK+9FuX4nCFW5cgDnQyemt
S6Z18OscrcjP9SW82bHyPDLWl4JU1PcitMVWtbJhSNifN+9FAME7rGvQDhAhVQEm9IGkW4UmhYuW
RZK6usdImX2U2ohqg1+ps7klIubI1hRddrXpyEhJZlH91Kj/jFJCTEs7N+0V/dwmfNRpfgGFBY4S
vgA4pU0U8HLyXhjFDeFP3aNVmW+4aTnNCwJro3V5tP0J63kYw9N46DfwsmS37pghunTZpj8vWcxv
jVFupvSzzcGGR5bUnBO1Wy6kpR9aTwGFvTnT2QtyiaY1m4R9CWTl1DOojQTgFbxGxbYnK2HCydQP
bzBd04IfHRJw+qNucNukga3BtryhrXuhQ93BsueD2J13wLXm4uBvV7d+LzQh0M8l/Byf1mBoXgfG
3NaOaMylYK19fkGWm/HGzMQZc0pVlLlVmHnB2nP/FMPxR94C6MBtUfOPre4mmHz0KGtE6P3uJBdC
IcebHFlXS2Py3X8IjOxh5tcYOt4ekDE6ULjZsBXjEISTMIYgWLyFW4uTkeG1xDRQmdOQnDojOZJ+
Q9obIhXfsmo11n7YxZjSBTxP/5StYqWvp8yPb6szrjHVi3JJgVMTJU5hnyzoJyDUCVlSHSc7L249
jqbIbZniEGF7asOJElJg8mA8mhq2cZDBLggCx+MVnAieHwQYUPsVH+oJbCBj4gsDk3dAGu+DqtFj
Ux2koZf97WS3Q/RI82A7hjy+z7axUmLtPcgj5RC399AEaHp7otEtZflypTMovNmmx2dpbzU/wzfR
o5601nb4p1FTVNDnZ/6xInTKCMnehwtOsAcS6qNApb4SVuhJUH0um19yMSiztRxrR6qcDInVvK8w
k8/Eg0XPxMGlYLkZwCOHaz1Iu2S2UWCVBdBwzFp9os1rH61B2CT2VnlGa8jgGQJriQ5j3QRoORNP
UzDc6MsrtNX5ZDGXzfCg7mD5wIX/OjM7daCen9RGlWMTPjiGqEE14fGeYzI8cUC+EWU7WGdINLRB
w3ioBv/uQpFrTTn7mHn8BkRnyI78FE3v/OeHhEJHkyb4yyeHWEIKpxDSgBYVujkJ6u8i3TBdlsZG
/73dYuney9NUKMovm7R4B4KjMAS0fYTg9Br8851zz5lc+5UmL5K7B+N1YCcSd42/9IYKAfPaeucz
QDlA2ZY3sqNAmo2NdF4o0qmTFyawNv5unUK7Oj7D5PajcN2CP4wQyOU/aAhpqbpnPHQLWBZcfG6S
ofth/1qrFBn3FCEqJB6XYWsSD1KO9GGjRm2JjfCfD7zTccdlpTfTX6FCJdOBudnV4tWLi8G+EVKG
1X+JxCOYGpK90dzaZp3vyweXys5DRNMMa0olVMwlL6t+eG2tIDRk1J8U5eYr9d3EjHqcoY00FhDS
doNY1kwt8dUy1D1HNBr1vzD1nXZcKyUKuWd22xj/ncCRs4oPHEbAtaVz+PLoK0vHvdV1qoyrYJM7
5Fz6STyj5HINe7MOxYRS3LI3bNwS9/IToovRzA4q+1Si9WdncvacwOWHBEu52tTFwr7UG2BJNnjC
k4MFxURIC4h7225kb7j9Oc6Dc2BcRCoS2+oxOEeRBgBgLsCBaWeZxR5xEvf3iOT8CaVLuBeXdjUY
MV5YEqcorvdv4WRCJpvmc23mkhbI9LRnidDVhN2Hp6vK4Kj8Qrdy5o67jti3IxbPqN3ahfRRiSEL
FOoWxNmINY34NP0a9YUyONrq65gVnbm0u16rhQPmiZcn4ZpAzD83EsLTRXY+wZY4o/LysDnzCqsV
ddZdo4snQ/Rx4p98QZ4iS+hwYxDeM70FVY8SQE7hEvQvV/YNa42IhF8t3FXSLCDvvBr3nI9x1eTD
+0P9gjwIgV8a700wW9DhSObqWohbIJIhVbB4MatgHa2RgMyO0QsKB+LsJywC9YJ66LFyN5uwh0K6
KAYABhskm4A8+z7vWzvUA/l4ZBNyCQJNbfROENnK3KvyGNLKaViOf7YglbAiIfi+0pw3F/dbNLv+
PGTCpEZ17WSkIBrLYrXUUul8EK3W8Y3yqx85MQgNT8PztWvFUJ4Ko4qA24PzlBXfiwmsQ+FoKIAF
d4i7O2YFeIK8lsC+d5LXVlVsjaYkeO/mGE9S9/YyaZh9toSfW4HHe16tWDa/iGFvSG425pcw5e4D
2WP3LddXgzf9JhRmBOXS50Ys1ABiMvAo+o+OUJP4eCfa8BUMHCGfdZGBn0wZ+zMC602RHZpA2Uqz
KzzYcgeP6McD9F5fMCLBT8l28q5aYDtWwgBhsU76Fq+tQ6y0jnobRI63qGauI08sl2QSv4zcvTDZ
WlSwkPYg+G+mouPMs3l7CWinJ/tCjJiZJBS4KMB1rLGz22cKNIksQ26Zgi4K3d6f8FSgvMP9AKXv
WINP6J+IMnHMNNx8ZkRBrJeYMxM6R+fSwVScNCtUoaLX81W/TOiLaLu3rYsskhSheH+hEqsCNpiE
46cpVTBZEuIPRN2nHkV13fXpuNPr1QoRsjRkHkC3seP4JwDxw2/P9+RXQx4RloVisugcPs1+ANLY
S7jXAzhazTuoTApJqbOAfSfC3YhlpyfG1OWuEJsJwt/gqs9KMW57Bg6KxkT1OYWJGqbCgdAzIGcP
aVcbOW4lsb+0vrl6YUh+G6qh+WZLTIAM9nkUS66514HUNcffE8bsJI8jljyL8HDTXzXEhO62kx8k
3+bXnUkNWjFvCa08whQh2d1iz2PvoFCgvO6diMpanY8DMybFKJPMjOnniIP2yoBMtHiDwpTyXnPR
bmUljvf6pcv2QZNAqS5AG46h9HLFbZKnamt8UaurOGwDnZH8Y4jgAKyqPG9ZrKwsheiGA70ZJ9Kb
anHHAmEIW96HK4RTPDj34ZuOx7nRJhpQp0VMQ7mf7i5BExwGNioOXsfZ1UKpHXiv7GFjV4QdePey
qbA0Uitr8v8vYH8CV887zWDiR0EQrdTWeZDrrWteqjrrtysc8aRMeewUeYjselDVvwIG1jve/ETP
diVgivAAaqghVIn2CW77NQCa7QRi1IFKxe+f2VhBt+mfU5E8MlgHnz+UP+oPRrb5ANOb2FxBImj8
7CgpZGgbhnD11+6qNZQ2cS/2w19JinGifS1IXoUhEPC0Fpx0lLuhMs8Tf9pLylBBTQnHdaZr4E4N
usKF6HqKDiLePiN1qYf4KHB/FfQAc8xYQMPp8s3ixbh6Gm9jnOyuhhiCkl6isiG53mUoKo/H8tqY
aJibCqT8mnK17Rr7KrNzKx2/BlrX9P3AC2Y0k5lAK3w3i4pL+hLvxrK8Lz1EONAssqw3rym/Ixph
e6bXldb2aeVLh66N86IYNtFT581wJNYirvnH43yBISVdshJuNX1nqq2BJolCnyjPO3MIn00DJCz9
mg/wJXMkgEY79ABwV9s6xGMXJXqkrRNCFCc+zP8VHk1IZS3AXpl/3TFQNypew6kys4x2UDpW6D0/
wfug3lgXCES3qnRDA4NjcLllSIvoE8OrdaWfezUi0LKwql5sU2+eeA8DWhtZX4nCNbBqZOOsZcs4
NU04mr6lPgIPBlIorcKJn5tFqDK+EeezKfcBHIn7J627dOBSSLa2mHCYY31WlAi+FkJdFSAqLMOJ
9XBgwLxhfy5FgboHVXGxylZnbWxuSVVGPd1xNU7rRqEHG2NuLmbVYwjjXm7h20LxeiKfnvJgYvBB
RqiurZqhLqVZ7VF2VjTaNqGP2GOKa6dNTY5oQGojCSiNeKUAlzYq+JBK61d+H9BDzM5e0yuQ/4UT
pmlLXBX8RrLkCcZ2clnFSDM4PXoMmI+23v8QMdiqQuHa3WBszsY/AG1vk46cOq+GNn3Daphi08sg
Mx41Rw6AZ+pQDzyl5WE2OLN68RXzpkA00OQ4Wn3t4m+GqQX6JoRDXJyFdh81bvLiN59OXSSlXDv6
x3b/pnfVJpjE2+ovvYWxmvuGpxCWeKg4DL9gVlz7dpq84oMZZIkG8UOiYdEatS+gP/VizOOMBWV0
gat7YA2cYaxDHu4JgyI9iCN0qKlhed3wprJSJfOjo75YXsh9cfs0pDFR+zi48A841mSt3UE1pCwc
mhYhhKQCOhqcFb2AyjEEPUr6fL6MjZ+sOlctwLdaBHoorm0Q5NfGp8LYaWsJqmDiXtjkPAxhrCTV
6sfVEIE/h9NS3HQGlat9JQmGuEaUlDLSPLhoghYp0N5SeesN7a7Vn+RoiAow2sfHaPsB9BjHiGLj
VDV/GaFaGxpJsO2tLOYQki7XWt2gPyH7mvW7os50oiNEK3HRVEDbaGxbDZWOiC3SWTDs4BCDRTVs
pZzPzQcnhRsRv4/G0ngPx63+ZScYOKAxbYKS/S18bvm35RCRCDJsMq+H1utKUKDSdC34GCDkcJ1u
iikKucSQVtZZmSsskuY1rPJM5E1NTjEwZFErJURVLWt41/8GNoURpL93sW86jtPbC+7B47o+fmi4
h4T2ji9TEVqYIlVMgmJMqHu1VlXNeQft902EOIh9hp2dhWE3Y1CFTLuWFEDVz8bMBFNXp9civbra
sahzEwk/RRqqTDWTGGEPB1h+WFOMssicKIdIDMI8kOFiNJoY+0cST/jnB9tkaZ19nigXBsMnvbEe
saBYox236BBVlC2YA1/3Bh3rbGUd74fbiFqxMToeQANP2jfEdRXEOZIvefVKCQsg+9YvCTGFN0nH
C0TzdbFZghjXZ08pSR5D+S3J7a8ZdgPuKjH/h+FBnLy4itjJmNomJSya+FIGRP/fzGzW6iDZLKxd
ESwzCRB9hpEKzr72srG3r9pZgIpBFP/q9U+h3+RBQi3BEfyr/3K+KLHlYiSyCtq5r/FeinpGqesX
IeqsOWTo5om68FcntSiezLuaw5ksAv3GFPT6UhFAi4Wnvo9m+TO+HZSs/4vZ1Fixb0yjQ+Ylsuim
HMXWerSrxTZel1K2MQIrzWmYf7Uem8rGvNwkskQ6OqCiNBOSe6TeaKHIR185Or4NeFLJmDInvHIX
99Y3onwTkWZtPdps9MlnNIgzBbVE2JzgafgkmdQtVF+Bh4uinQkNJ4sSqmQPRvEgooimuXD6jdkM
sfD3t4rvRdkHxkQh2Vw7K+6vqzq1K6UTQq44BCn1fgvHo26UGiGEVg2ozypPbPrtGO3jzkQtoBA/
CyBL3k+LOcF6659k5kGVKdYHuq2fd15AgkL8l4Up07XKAiLG7DtIVshPXZ4MIvuoPn++ht1hhGjl
gLy6M7dA/F+phhUU89uKqpjAV6eIUImChpr8JtiUlKa9sY3isCp7LHOwSvihSrHKo9vZgalCvJAM
G5MUU5ZEkQEgDUMwXbnWtrFFSn5NS0umwODDXVEyDksCc1xOZbWmD+uy3U9z1kfa25E6fwsvIaue
RHjtpTjZ1WvMJUH6EAZhAqEH/mSuL1HikotKrhsH39OMMCnnvYJ8WOUOkiHAiJ6O/1CQZYAz3weD
kaZinvrevEUXgzmaZX7kpvIuuz3wmFFE4/ucHQmDnc3YZiaHhw9AW2amJtgbwlFurs2hUZEK6Vsm
r3f0dxL7Orsw+A0B6qGuBtGvevKpUWPqxMe22JG32r+RljjiXPImtvWYAbmwHa1pQAldGxho008G
diDBuetVAHLSHgt20J1wSYqKlNaa5Fsu0U4u8ZDK/Y34srZ7bTZGh0+MHHtajYpWV4dcwk+0mICy
Sd7qeUKvhaUd+huaofga2q/gaTev7ZdtAArszLfVeEvC/A2TI4Tr+5n/isde6H2ckqvFhJt+jeEW
sBxN05juEQ9KiiF/NVWnZ9H/UoeI3QpnXtvSaXX5UGxkAeQlKkBI7r/6Ie/yUDqYNuVYy6HLQLIa
0qqXejQE4cdM+ma6tAwI0OHwXQ+WFuYSfdnGh9dSstmjoiWYwAADSuJnIKHe57b+tTz/1eG9MdWU
+hl4p6/Fv2rN3FUUvEqUpR9RD1UQtmaLOuqqcLt5F4nFrzyzAHEisTbRnc8+OeC2NnV428RoxwM/
qEudNa6Z3u3qv4RxT1JN+1hR56Heg8NRjgJ/9wZNf2aFLy+lf4Zp2NGWs5KaBc8hDLjvfKSVMHEo
TdKQslQFcESNbXPgojLCs07itDW0TYbC9rhXk6yzbR52b5a7cACX1uA68k+xM4p52V3UIIPBXbsh
3x+ghjhnOgiEu5BPmtHwS/nJlVr82MJa0TwLf/5HhxA+unyRR9ixSB8TBEhOaN24trzPY5sI66Ob
ACCQ22WS39cPlkXAFkTmJXcLiLOk01wQAs/WcFCN0MlydslTmAtq/iK0XHhCM1Pyrx6KTT5GHW/V
CuxwKIf1AZQ7kQNfMYwyEvI5uGK/qjlGsn9ox46kieQwnz3ASBR1xf4MWCNQ/6wrBe2gX01O5DKZ
U6v2pxEEsNDi2GCMVvgrk0TxFASHx65aF6It5tpwkH6dVLrLRkXI5FmvnfPwmkefQCSowjbeLrzt
XE+DjGSBaCqygXxK653vTzpuDYjhFNtgWUtdghBbmmTPcpuEeJtwAIonI46AHV0yApqt/tWMpgTi
miuCjs/bQb03D8bmISWFdjwpBq249NvctTdBshmJvL+u6srTjxmHG8ehCRGybZ590I0UyxcoVIC6
NqHliPCZnCoaNL7c9K0a+bj0265S9XXhUlb7K9ycvqBcmsoJUZYs2wGvrIPq7uG+qEhaRAI+gmTx
8iQh9LU4uvGOhVp+MlP6Uh+Coguy44VTKSmV4KZRU3tOGgb29KSDeFSgJ+ZzFk4aSY596ITfP1Nr
Zz4U0KKfDnUGf7XMn72xyvPY/VFZ997ALs+RHrWoAY/WD5Gh5q6bx/iZtvVCpZpUPg7enavm2OAT
TCB6dDiLDROr7BP+K2rdKTrARJkLg38xQuvU4iIpmsiyZjHgshoMYCDo6RmdY8hD01eGVS04vZ5P
zvI2SGXopdYSbIQGR08Tu8fdCc+4Q82Ok/ZA66+od3U1w1OpB7rORM1D5IaTIViWZqnPOp/xDT4j
Y4zx0/ajmgTFiaQbha0TZd4fMDuUnICV/wmPuSJBUlKhmDsiDfp1w5DtpFkbdnO+JZONceQNNWtw
lfIJ8C2+4jRNRWZSHq4yWtRdAKxFxrSkRGjI34/cniEV2HYksFJsBpxvwWYfIQrx39QmsEmtev8M
SJvNcUS01sdpeOk2wBu64VohuXOnrnIsUM/G7l1i7/pNexQHCch1FqTooTESmu07qvWGF58LdPA2
wJCJUljRvu0M2MBiO+H17wB9cpCQ39sT5B3UjHlMAFJbwp7I90KMK7uviCZZN6ECHC/bYrQUpZT+
WBgjQzO5AArfF7NIWa8xZLHlAwKuCNr5bKrosbQXjVn1/yfEpQaZEkxITopWID5Bn3GmfgiYCyeu
Z0Mg2UYqLIxz05XGvq1EqLSrkzNgF2IZecJTNh6dg6yI2SEUMp65L994gNY+Hw4u2lB9q+oxFT/u
M7lxralJTVudRDDNs98zfIgh5sRZVN/LmXGgeW2nS9Mit2Lz7dAbZ/8JyIxBgOoBksy2YN45LuYV
yXr97nF90sl4ZU/69GHe7UsI1PNJnarVwYxWPK4SxRQ7+NwOTqDkkZj9z1aBanbOPGHpgom/o1I6
3xirgutJZaYnaPDOu7E8ZMYZBGR1HRz76zegf33Wnxiq6DaSiJ2apH7H3TjXRbiZdZvUmfmVZRUn
bSssvZ6RDQ3XC0tC1VkxjSt9qBHyLxUpoRFNwfhcRQIo5ZUfeT3nlQQlp79M0wkPzoOi5xhIaR+6
lVDVnyPPyjDVmCYgEvJk1sB8s5j3Uc5oym51xZ6PdBxx6yl93z6i5/3dk67Gs1ELQRb7Piltuihi
Qj0gp1obIychNr0osUGdJztWw15Pg6fVxQtDZ3CNFqFWYhiSIcV3umFTgP33z9jdVfmxm7JvHoaU
cFdkg3PmISYMQdSfh17rr4g/xBGZDiPcOmR7hNG63LCCGw9N/gx+DMwtg87hdBljmIJuoeEm2uL4
NIzg5rlHD5YSpDx4dc0oK71K1IqC+Y8Nk9rtyeel4atlE5Al+bag3gjH1mRa9h3LAFcMGad2jCj+
xh++mfDb7h8jffn49/Z+Ls73nC9QQFA5BfuDiCRBe7LkSxDfhQKSgOH4ta3RPylMZ0XNP1e1UM8P
K2d/CyvK8LRJclGqqd1xxIDUtkp7jP9DMo2hmDneXvb5Nskk3CZNLJ1f/sODoRBwEyztFJhPGqAk
dr4NRToKdpwpnP2VOVAX2JcQVQPLOWgC790HD4BRPF63GNt6LySUOEx57m7T16xSYfBf+gP1A4ba
dtVPz6V4YDFu0bvSKTnY+AvOsbMF1JzXnELTWrK8qcyyeZFVQc/BQ+vm4XnKdvDk+MDEmGJk559g
wo9sPr3+TO4MymYWr9XDEwC5axHzjIIaz+Bz0CauisovUhwlbPY5C4HoG5ui/suJ9EnyFix3OP+x
y2ogN1fME5WOowaYz1ZL2vow6zP3BpDxKQxvebeO/C/39fcqwCBJUbztpuYhojAYQ2+2G5Aje9vH
IB2YfdoLPu6caDOEnFz40F/WstKtXEtDaTbN4PQQCi8OIKFkoN4aREV4v2r/zwLnI1U4iP+GJuA7
FQAZu6N6C73HgqHME+X62U2mz/Vvz4fLOIB51qEf3MJRnfw+Msyh82+hoPcsKiZUGGsBluCDjleU
l5aRK65xaTtMhTL9WSCMPylESTYg8nTALL6Ireijb474F9K9Mmd+XT34zKxmrH9vG3VK4F8PHrBo
G3fwivPOV7fl0hstxSHZkXEscpFP+BVpPVg6DKbN3LI3Ypa4nXtg5jrnTvwzBXGQjy5J7hpAS1ch
Ughj4b4YqdGBWHQoZQsIdi4BecV0KSuwV2gDjtlmEs4ZTQvUgdNzV5Gqkosb9in2YbtLDuiEkt2f
6TtL80pwy25bNjfdrqiwYiVLpytQTqJIhBzsPHU5yr6/7ixbNOkFec/PD/WiHTZMNNi10O23Gd/D
K2d4ncrMDHh48KcxKevCz7vKJBLBEBa7lz0MMCrLz/6yWl3C6Rx/BLhLJ2cqUjJH7MWugWR6MJoQ
eMB4XpB1ohs8I42mO8Gm9eGP7Nz+AtiLy5EtC7fiwIBr//OfbXLnUhuK+5xgPd3NbO7RFA9GTHP6
BUpZqa1tPSu0P2MOgo0lUzBsJpaM69WMOuua/OxujSTrud8SB0kMWN4+HnS9sTK5OtmnTpkcwvY5
xuy1WB6me9kCZOcbGnyc2aGY5jo0GizmQxF3ElQ0YnYCQ11hV923G3bSAyHp1fG48wPG1ot3YxYw
6sD6SG7Dr0jcY8zQv9XTUCiZ8zAlNDr4Av9Y24yUMBMwdWOOh5izou0wv5X4CyI9S0BnpT2PRgZF
QmivERQ8BSGU/gAzfaTMm6kI0qbMziuQ82qUeDQu10j3DwZ2YYNAFAfy52m4AKYLc16vkYZX0Hie
kwUwCBwVLk+kvdVybHCIFRJbmqg8czDUlLeU0fTul6vzl6seYtwct4oF1M0vkAoufJGBSFoaHZ4P
ql6RS52lIVX5C3DNUsXzKOvejmHVs2z3K7cYjcael596TMyEJy6FWaBDPIEJBnFbZ5VU6ul4Q4f7
erU53c6pfJQv+wGQHbqNbGJl5cHvXP1TW+VhSKUOEoZiKDPcPcAkYFoaWIDmMcbP3DqLU6eGA5Y/
qGUbjAbSuYd9MPt1dZ9mUK3p6MTRbyidZeIPChqr9vNa47zPtL8TLswJJ9bxBbbXFgXULgNPIoui
JI5NR11b7okkA2rvXESBi8W2VI37TrUxCrVc6drZvan4CFWV2AYIUhkaPsHpuN/ZjlGO97ahJgND
UImRRN/QcemizZGNlmp+fPOVaTJIzUjuIlZ8eq3S0zcrPr4duCQabxZiQ/G1C1rhzxJWFTW6rgpr
qm8wOcUBzKOTgEEQ7//irUM+UZ8dbmCi90CxQSzBcXZ+y+3kb++OT3AyM4+EyuVEmjnBksOfcALw
Y18HZ++HIjk36nRjc7P5ZivpU4vRDGZjJYi4FwjrdQmZGGK/iJN13cn5Hz+KnaaK21chyX0cMMh8
dpY3CXCVW1pTy4x00JPdfydm+oJQRAwEQsNHJXS90CvRrZa4lpAl+ctLzQDLWB5fBH++Zaihvqwk
zwEyEUL7ZhZQttkXtkGvXVfv0069xUnZbTteMRrWeJXooc5QuprwuymSnLVR4I7SbX3QcgsGev6K
uWMuTS021Uh0Q1wznXKeDKap0uuiHM/Hsy1RvBFhm162Tchmcz5GMugTqOGXAv6Lz2sW/kpxmxbA
459btmOzx///vSSFY2IcRqYnXk6Ao8v9nqGMeThCjm/LzYwJK8EjjSIBZ+n4Pj63jNpsTXk4mskK
1epRuPdS5PRS6FpmMR4DBs+quErAvs5PR9cNFFT1ZDXiS6L6WwjEsPm40hRHzVmEaJmTM+LDCbW9
O88NENxXXg9mAe69AoO76PVuyQjRQ73Pg3JiV8LuJoTMvIouv79eUYNvZXAbL9Vf1+YQT2lizqN4
b5I9NtNRUNIC4wrx27O8DhRrTXLrjlCTeMVyWPy+mIXm11EVMHmAGTftV8fZ6hvfyYaq3z10GQhA
AOcSfe8yYtc8Dp14yamtHCmAFRPcuf6fHiUqk0o+ai1r+iZnwCBWBv7EJENjReWnfNGqrLIU8upx
rFNjgCTyzhzUietMSmKyZ2LEqcTHZ13mWS3puxp7a5XFk2RUxTyLEPamQuRLbzKUp53bD+4YJDl2
JqA8hu7KxqGqPmfu2DtPZ36B5roMXLj1F8rwUV+eS+Qm6YdQ+iT0HZYXC45i0s8wgOw6ycU6FWnD
z+J1IcfZKThzLB34wJsW5v9OQqywbSNmA2ynvyiblSzAcS4vH9RdznMt6FZu2ULPhdqBX9qZ8dwH
i0LnnxNgeJi4Lf2ZnSoaoi2opgQiBBPzMT+OmBenFraht1cYkyo0AoEebVFDiodSXSq3qepIaOkC
lFE+x1+gLkVdP0ZD/Vg8nkWbWl0NfBYFKL/T+3YkgEOs8LMeGtlux1+zbY3sLTX96HqotHM7+ebl
SXAKqWPldM8jVJ1merLGAepfXpbw2ZPJfYfezCpZQEqDBmSTJDD59nca1Oxo3iMR2CxuwzOT3Xiq
vG5Mm6JtdUWtauh0E/SHFdeuKgdmoX+5xh9tDvGXiSy7G/Qag+mh3FvIAXHqyIka9+OP8Ewyj7AW
H/QYli+yG9OF8ZQdCiun+Ddr+WLjxDKMN6A7MSyDjIwF4JWv7CvfReQ/QDBoORCazOUGYjolUoyj
QJaTEChPOdXPAm9QpnFJbc7ZI5vwUUGlgTMU6bmNfKSxoZcBTrmz8GzY5GyHPwO6l/OCag9q81gu
aDdujmVdp6Fi6RnmiBATqp3i/tkZY3nzyQ/bO64+HlQ3aOkB4jarqBzLXmgsSbxre4MX/j4bsVsT
B48Tj6X9ZSokkEEF86b/59QSs++jdaHXg0l5WzbxwMQa1Rpwkwx8G6o/azUmOvPz8T3KZjmAf66c
q1tDZoGcOk7F+CL57ctzwz4wt+qsBcFtrdYsRGYyHAZAtzMbWZ+zjDk4wjtLCgQcRkiwnV3CDgd4
DBSprSb/GDVg058SBlxM5scUCPHRBoovon7k9ZjPXkE2aAXEhYaAUNpdbTyjE9a84z0EoGXEs8FJ
yqedw4Q22wayUg/bRt2tNoFo9QX/bz1Dux6IIinhZd0tl2wV7LmBcckOqmF9TgfGmegHT4pfyZk/
FaY1EA2dR5T45J3XSNO9IZVUqaTOIg3/eqDUyyqOwEHmjcv41+UZs8K2acoHyaYOJIfewcl3cpN/
Ttj4/Ce4w6UZ1zOSNToztgJ8PKfAcZ2lVCoXTZ5XQWX+CX4j4COvowtQphyjmpr/DWGHkrlFDxHv
scCkt8yKqK/9H8fUllx/b6ETIdKwvexaTUqjhzfkWTWt1zqcT3rpHGXNpflJfyxgSpI7bZCwFJf4
hNrkZ71xeV6Q1mcpDD0Rhw/ETqdpztv8lz/os/wM9mhkkKaPKTwATNpgHVhzf9LckIdQJwEAN7zP
cFjlYXGh62261ysrvZr0yX6ofO+eOQw/aIxHvV4/sZOUWBeHn4jhG9tjlJqTyIcm+zIWunx1hmJ1
6oKLNMFMxTMjQ9oEwNwxAvU44KUENwPB2Q1C7qNEUe8O97pT8UOUDPapl0pgjiRc+OiG6ky9uW8f
5w4pN46Ai31oqmL+EnTos8yy9NrGsQfkC8ib7xVERvr7+LvvN5NfV+pNW+1zKS2sPRlCvKO2j/KA
phnKBpRf6JKS11n0vNTVMUt+AlQq4A6zeF2Sn2V56JBiiJaqZNUsZgFSRYNpA8/G7Xyh2fIpTusq
OX4P7PkELLw0lPqTmYScj/6SeI2CiJylEPTxeNUgUCUQyRZobqtbuuNEETvb9bF2wg3Suie0eGKl
10nbH3DG4e0iJmgWLSz48LIhOTxPFPTFMiNfmoh3uQLu+wA3JpMExkT/pxWpstuHOGum55NKrhAd
Q/DTkvwQRi0K5yfgj0RDAR3T1bSNOZEUP3a3BCc7c+9KUhLloCAE/HstyNaQcflzumJ7FocCp0fa
QoMIyDtRHQxKeHLWddObWDXUveYWtNU9dSQLPkHHqvnnips0McJmBlD2SBCPSYFwp9gAiAdF8GSv
zk2xns9Gqb3SdyJ/V0A5LVftgJLnp/p3GJtGUU3dnmNyTOzTv3F0n4bUceIL5SqdM/D/wB5K2oPe
1QSb8XlKgHMe1diar8esoR3HC5lla2Nxacbm64gy/plOPV6CUCOQRHadpw0gb6x0KoFVIZ6QZ1pI
M21SDGYI3sMcjvTs8P9T9udcAJgK9UF6qC1gQ50W+Ev7o3Gn9T5krL015pPd2ghAada0KZB8XCKy
kTXDIh0A7rtrpn+nAQ8uw9l3cVy6xBMc0gK+KFJoVhAEOSKVXpd7leWD/dSMpNJQa4DGoFw1UCyU
CIE7VAq2+c+80xGYrtoxCxf8u8+O7nBVixgTGtQjthyiw7vwmKf7bWLAVU8v4x+zhdmtObTCXnil
kd1YA6qHtwC24isIUAsXmpBFBpoNVwE8bxNQdio9fMCB8W1o4Pc9bo4m7O8DNjNJkyIZTXRsfQYH
yA29EnBIrXshh8RkTs3fA0WUvyYQG+dwYM94cqDHCB3fFkYl3RSteXLXoA89ioziJDHYEzcZTQkr
hefUKtvlYJNxZbSJW5nxEG2RqkwJvCs67DB0LpoHDCk4y1/GBCpwSoJRrjlzlGHf/jn1qUo7yZkm
frFaa2ezPHxHsvxkhtQtPwkLK+3iTDfuIR4JMMEAt1SxZmtGponhb5in3/hKo9QT5hvw6xjFVmr7
kyYsI5D06G8KwxkGkp9Yuso1Ugq//zxYv1bNk+87/NNC3DicFYXXlIxcJOICOhc/aaNDVFtQydlb
hOqoF70ri7MY5vptDCa0Yh0S5Ao6SwfuT0D0ff+MhLwfzrWFB3If6zw3Sbo1i+2fV6NfvJEld2h6
o+oQxnNAtN90+7L0OaIR+dbrZJHnn5olLSrFqI0OewGZKAVsdPkT1bJhdU44iZAY7GpShz5dlNxR
BjG7AOPR09x1npwXvGcDzUbb63UfDMHADLyr6vh73Otn2/1upFIEJ9YUM/L2Wu/mYxBdsgJI2cEz
DZNePnwS+UkST7NdJ7BhCq0xkNsI8k7V4Qec9TNcdStT0WOwt0qBLu13oHNeFX8SOXbvyjgTVQP1
tf3ba3ikB9VyTkm7gYs1KDGdTvY/Y7zdCWWetsDRXZ0WzK6ou8OfBbKjO5+BXjajh6vsGzu35zgv
U8MJ0eoNKHGqDpB2jhc2Yxiz991cTGozvw4Ck5DORdhNBizb76Mrs9PEMbURv7ne0XryAUVIN/ZR
OKayLeE4DxZKSuP34GD053hHV6IxceVo0Z8756AQYRCrJo83KDb3oQ192AJdyPC3u8mPg20P0gZj
u01bNQe5lFoZBsBINx3b/iOYQw9fjKdcDAnlPCToaRRL2zcN4XuPbyO05Ka6j8OSJy+Hn6n/T6WF
gO7QBeEDjNNgSu2l+HM7/ewN5B+jKWYhq27wbURAXrb8VChCNBBmIdnW1go2gi0AxuuXACb5zRsL
BhQchjNgB2xpJpb1d4HI15uU5vAdGXjOI9m32lFaOLuvYjinPlzejeljAxS69iEYCqEPsy+jqJd+
6rq0tVORGdvWR2+1Tc6VumpTUhLOKWaG0P+G7GS1vFpvc7YNHKcx09hGsIGelAKiWEW+f81vu3SE
zi1vNd0qDfBiqOJiTtG8btYHAHPLaVMcjdqLPTK+9N7zT3tZITm/mpiZ6yBayCl0YiodMs6VFHBF
t3u+vIH4JZX7F29ybZivk6qRywLlR6IM/6YWhJgZoIzmGtfFtIul574hNQE919CZBLUmEBfsm7QR
SXdIxV+6Trj8EEJ1HUv+YsTgLpWD8lKRQDXOJuhoz5DKIjDi7TNf4td13LiPMWryG8mEYY0VNblC
++YCZphNKi+SpM1So8i+g29/xJPDSBk4lw0iCD69sTvQIA2ZTkCnTwZkToaFypHUIXPf66fbfmsJ
HTA1pkYtnP+CDzo2byIwAcrCJr7XUC/vIQZjimkOlyFhgnR9g5A4ETSOLdrZrg1XL+se1VkspRny
bldVcIt9zgNOk+QWZr0FaQR3IXni/pLhA6FL97RLSIFEBP4IHWOFSIY57KKremQk//6EYiOy8yqI
YAlfNQztGxqwMuEOqUg0HQcqL5qEAM7W2wSWSWntostSTulPVwIMXSJR+T8RcB9tepJV5RGlA1R0
BQ4S5VutFZl955WhzQxpnQ4S+H9LpwK856ar5l8UveTap4evsj7ySJQzDqgUnpFG7WAcnat91nvy
8L0n9Tms8WmuHO0IInbsW/FP0tgXt50dDaVG7DqQGy9Iy2cJ6UN5SxtDnU7P4EfqTEc1il2cQvBX
GaG1TiOJ2K3mddZuXFeHvHJSrnm/XVtwYZJEQOHPREujodz2XGkTz+sgdnZdbh/6LL+gls/T5ZVV
x273VgO/HNG5u9sLT+DyRqUqrPwa4R8v4U4/5ai74lxHVJPICy58r1NFRORYoxr7U/9R40IsO210
kZ70jrFrFX9gwUwTwkYD1KjUe+RAeHl1Rr5/KEjT2+4jBSoyCA8EpGilyIw0ZdvaMQ/JK/tiwlcu
Ck6tZ6KzpSPN27DwNV3F/YAGMFGf9f5ZgckOim2ejfJjW+GffcLvSHZLGQGTITQVTjBq7O1i2hQZ
W8n7M7yoYbX83N7f7UB5eBgwQMoxDIVtYdRTCPeb6YEnK4e6bB+NfAadUpv+Ve2niqL2X8dMtRIG
4LDCcfBbKGgLlpo+lOQ+8NNj2NGXJnCIi3SIJiwOa+CQqmqx8YSk3PyQQ5AmIEd33gLdrAH/6nCd
EyE6/5Qzv5DojRKEw6aaVL9FUmSf5B6Pdb3ZRyFroVjoJeZrTWgRb5zZ6V8cE3Vt4eU9sn5tpzdz
6fEYUn8/sOftyyVa0SpT3S/eVOhDE6eI/AU/71Cu73VNqFgqJ2O+5GuLW8TIgSjZL9wYXKmraDnq
m0DJUJKZCLt7dS1BUBEudiMryMH4LLsZO5AJ6Dkf8bKnrMfEt6Ous1TZkvcezVrc0qIVS1fD3u1+
PmWskdvnwu3LPPKHEt7vRPdN00zIdZajxpTeVtr+9ctckQz9Frrh0toVMttlOLrXVugX/QPndaiQ
YWzZJCIe35/BLFhVY1xGTyxhw7vV1rgXiyJNkO9WxGaxtBwSvXtSSKxX4n84dSB8U+sZGOcyRU6o
ySeYaDhaxxiVWafvBMhEkCKeg3DlFaDS22iMfgFDCN8rydTF/G38/Udj/2ZQ0CJqyXBTVnfysJVH
9UpjLuETfVmy0tN8hQnmqw0SwKQP25touANpzqRVGJ2qcimOtq12U41K3v9XPHCW+a8zq6JEsPpd
pxZ3+Zg0WclDOC+QGoOgGJTpv94QAiX8V9dviCy2gj9SpHzCA3vRbple4W3Gf2PuhY2qurBoB+Sa
REQrUHK0p+JvThZ+6LRAIrMKXj/QvBoeR/acTcNFqUhsMyS8+nSIKAHdveLqErbw0idwRvlSF2O6
iT5m/Papu91ThdolLmXQTgUo3GtmrSTKw5T/J99xTPsLFj7351HXFPj2XYULlKd23LMSgku7yqbZ
eyf3+uiOsnoqSierNiz4ckS50+YR+e3h7Uq9x9OhUALADkvOpx93hLs46MbLIcrUEOEVoqGJmLSf
wA2ilF01RPSfSxZ2nDmSEjEkPjM/gX/pourmEfrfr3v8R8iJQanM5e636Pp7KaAcfc9I8VPzRdRs
27yWs7Ug8OF1YkVAzUSQRldJJvJIjBxTFHSOp3/q6Y8G5kZY/PrFrKVCVNUrdCDtjnI2gMIqbBwR
thjbClEQL2N8PyEwCMbBL2CJc2NDkDeTz0zEtiDDrRIEksL+BNGlv5ygE2YV89QSsfMCPq2lLgZM
AfmLxeLvaeEcZw01EFhSinrEv1QRnWNqmc+SHWJQdI5GBr6sJtEpB8aYCcbr4kE16xN9t2NaSV2p
6VOyLmPIZ3uYLKuWh6n5KyvMOUHfsEDkmIuuJWQO8lW9/gdpnAhP+jovYu9FBxGfpYuK476v4I/Y
TSOZc78gWlUSxiCTocLmlVpDU5kCagRcFj6EqwI3QA3u655KPMIfirmtyniqnpCuGknJO7w6TMwU
3PoKYYqQY33MltZ/ceq9q4VFBaS/ncFxCqqWcAVZ4udiIz21gCSNGgQdi16yDqL+6Qze3CTFI+s3
feAJtzx5RrJDtV6iGdh7TcVMSKGLEE07w5RNiFxqjWcAaJaRB/N5GeHefXb8BGXTOvBlRqpTzOXR
I52RTPTj3PezyLyi5kJzKECF298fx4In7bCy3bXMUR8bitt4IL4GlXm+bR2X/AuwbU19N0U0mDyG
T7S0GNAFaXBJ5wgPYpyBnllLIeK50FwHBvpW00mNzl9EPLC7pmi8QNGnpeNH1l8qec8hguRXbUcI
k7O5oVe1WkpRvWim37hkxafh+gPLWp0B8/5lvl8pWC6vkG76fa0X20e6xxlnKXr3E+xn/6UPInWk
RJuowNTuRleG6t+DlQYMA1QqKhSKrD7+bnnraaYRNfCSc+ykd2ipyL/A5iaq5S3EYvLMTUgcTZ6/
h6Fer9OZX7OV22M5ZF8aadO0soAAaSEeLpm1EMJy+HAYE9YVQvwncgKL2t7JFI82my4TzJwdd1Rs
ZRJBBlBEplOmvmYL5HgFKjHPn1Io0vH8g42DCOEFsXGXKLQVPQ6wLXoYFtZmL3cM2dkn/PfhJ+Kb
0u5UyWCQs8B5gGpnjO0D1OWbUNdtgMLsAkfVbCT5QnQq13enhvnDmpV5ySQNMKRXJ3HQfkkq/tWE
jWmKpjxkwnV9oBs/0HCwe6ptANh8s23sGg6M4pLFZH1wR9lvYgqyKKYUEDOuKM3tOehBU3+gi9DV
fX7r9EG+TN46NfnbfT5eq3We9zK6oIIPaycXxZ3NvI6MoS/rUVAA+mBuz2Wy1TA7UhlqtB8mQ5Cc
8Bb4xtVY7vFz6fUWKaXuI/y1gUgNjGUeBSyu6uzc8qtkJuGSBjKiZGLV0k+z+Ttv22nqOS9/JiTt
t55kVZ5hMlWZ7g9ca/AaV1z4NUUuRCL21jPOfb90q2dBKZqm5jiuoVYy3UuyZZe0OFo6xa+u76V3
DjlXF5B3qTE6/lIzvzcAfJx9FYH4piJVZ4mw8JZp5wDOHbHZQoEBzGY21+kkn8WDacnkFDUjSG0/
eapS1JAYZobwY2LBuQJTX/NajlnylvutLJOq/Ydc58vU1QwXTEyf1g6LW+RyxOdXFKHTgYYzbRjv
3ddpxO1bu4KYtvVCYxmWHeTYY58OTVyxHUYJYJLSW7aMcGNaL3ULfAfpOeekrahF7W5e1beHDYuM
dfQsO+1Ad61ufr6I6AnXMXndapcxU0xxBHPqlPhT8oVL+E/7JQHJQbYCIH/FFf9exmH9Z9vl3uyE
8ifXlhlDkEr8mZXmjwwJPl5qQaHoVlEhVgt41hrDZzPuxP92H22/isUtxO0eDSc+mHB5VMvx+bwo
zfENQUEZ2X+OFA2z2ng0n/WeTfnlus2+4VfxoZ6Y3L55tVMVAwwVYXxizQEKPHZYHAfLecH2Ef8c
eAcwB4KlOWyTtxoz3A67tko+xumqdYcdHcZOAI1zg1uhPE0qaPZG+6zmeAuL9kCPSW84FTm+bgUO
9Ov9GXy98iWgWtsY/YYYVTTf5merolkZmREpenhVPA9CGWtedCLKFA24jDfNNDQTMoew81P98brj
K92lolwb8G11+DXsrYvpsV96Px5mousUQPICuCCJyWflClK2/F04nsyJ/kvGGFIMxL2XHDbTSahM
YzjMJn/ILPI1+YsL8iR25QOvFSiGgVon92krrDKwZ2nRdJtT/vShwBjHADrUSwLTxfUHhjcw1T3S
I0+MlPFzxiUwTHUuu45QpVj40HWrc1QgWJodwNeIr6rYQ1QbZ9TqU2CkY4AZVLVlrVdVJZ0EcixO
nd6zIMV91gJmONRgcqaT6W8fTk3W7PAK2UNL96trBp6aNIh3ivjzgVgSUVy70WehJ47sKcF/QMvI
SP6QXLzJZCZoUFPlsYbCEqut6VxoryQ5klYnTW6xmWiuLlZqfHDS3gQ2NfaCeH7uE3knOVRUhu2s
MyCfoW3ojna3JFDxKOKpZJfC1bAc4UHyXq/FTVXfK8YocKePIHpHrZp0jV7fUdCvd8N+sApdAfG2
39ssxBNZ+V0oReEWDAKEfZ8Ah9aq+hju11QKJGY4RHD27+0wAI3+gcqaWkMzkw60AUVX84kCU9v1
27iN+tx/Rosfo7ZLe/Wjh5Q8vzyg3BpGZb4PVLKFUTd8uhGX/6wPrjZehSNucp/cxh6SBY8lFl9s
bSL6VKUn3MHb6Qi9RZtb+iud8E8PfEppwfQ70hHX7sSciaGDaoKWjCPJzR7n0FlUJ+NLukox/VBL
QLPADqsArjZDLU/XRz8RaVXHdR9uxgFl0EsFaERSoe+donzx1DjwhcLL6GO6pQZOamcXgP7QuROC
jzOp+AmaGDq8Ht5vnFyQIO5sewGp4I4gVYqNq4DlQ5CaE17GSOoaZbNzIPU2CpRzF4+mscp07XD5
/naDmazWaO6852hNeFhOGyaNDCHLX3YYzWYoP9fo+4OfqRgeN7FswphCWrhtSTwMF8EOj4JkBidV
NOTP7FqJQd7o99W01/TAtuHa+UOuOJn7+27dOxeKi4xDjs+S2q5HQ9lljgQbYXgxky9g3wKtR1aU
XUtL8EW7WNWAQeyfgrbqGmatLduhNcGtgMrewilorrFVPxzphgSd7F8RtfQB7lPULBHGKzf6GzxR
ybglgU/QRLTtFUATVWalVABBkbkzWn7u9KORZQenfmed7w2PyI5sm66f3Rkd6eb24QiXjtDDgD7j
BJs3BSJGmCiM7HTI+w5t1mXDtWI1G8p/UB9IUXdwzWpk9X1w0hGiwwnkjeU5zIcxFBXLTB0xDhua
0dw+/G7wbhOuOP4RCtHYOOl+zAINV28t3Ne3KPoYTIgXM2XClQRhVssGAYmMXPEBCf9yuO4OcmJk
z7hhFm1Y00Bpk/DZjkJTxEu9JyUqhTUZhIJIyjHPMLEMz4YJsRVJWZExjk/s6Lm/w8IgxCPaVUpM
pH4BJPEI78wb2uzNRC0wL83VmmcVGqTZtnxUKnainQB9LNHDB0CquuJGAvQYtq9KYd9OewsI8Sja
DebPrFvlwQJbBNAkE4/eEHLT88YhI48NR9BJ7ZiG8htwT4DbvOCZMNfTeEUtUpObQThe+zRx/GP4
GJl1tBPi5mPAjh9Blj6Q+GumJRbeH2JI/MRFXmIXhmgfuKk3H4VBAZBA+P2HXSXHaTYuk01OWciF
4tknOOsyOW8BOl1JzlCU/ywQweTAgV46SfmMAwUd49Oflq4uefhv/jNjb16i7usHbpwTbYFMy6aJ
f3KG1FW/EBcHCMy7yPLPUBrXUFRc99u7+W2cxnv4ZtBSl0l+P4uxGLRhmeZMBf+gyFuh4lGuobih
GLSNSsgVOn1rENFUPO1UfORxhwwNfTdFRTJR5Af3T4AxFIIv1FaX2Aek7aheVs09YTeBJeKEHLqQ
owBbwc0OwNJjkXPEZoAhtdzXWIbRxHbFLY10wqQNqWAFemP7isSkkiyHX4zv/Bp/fsaPbNhMbSta
ne29cy2nUjnwRsjRnfdjxucOr8meaxs0JSsXhaUtZ4an2uxW+eu07lqw9u55A0NOU0XMb5kkhK+a
NDunPSBub1U2vI8pc3444mxOPDO/7zCN4KoHt2vmROBrXN/z6gFZmd713Flhd0eHBXOqM7DuuzAU
HMb9VAIBQTWE5e+4at+48ub/Z0qWcf8ITcMUVjYwaT46AuIKUv+cKeXAHl3VbOUmb/kcN65XwRfb
4auCB3JYUz9CKBbFIX6sB1JBKADwezp003uOpej73A/0reXVevXnm+nOMne+17L6Ol4nFpd5YYMh
oGsiy2039YYB0IneWkTHWbXe1NRbENQobqzG7Dp4Xttn2rL82RkwOgcS+rw8wb5/CVeAe+GYMbrM
KEcP9Z6TKmFF4BlVlNucWuw6mxlva4MueBKn+zj+gg/HcjTkQHSSp36Gor8YLkNR/WPKmq7/EYP6
D5uljiVvaLt6HVpT6ArAM8W+G17BgO7SJ44PiJqZW3AYdjtbjKiBodxFLBcqIg0HlahiVQU+WZsA
1e1M3xeKOsTCwivEKAN/DCx37ZPVud3JtPjlciW0EH4mJJB/ncc8IOS5HQ/rLOf8+PYOowcD3JbO
RQEc1kaTRZOwk5GYWzKE7wEpjYBunvYWoCuYfoyak/4DFLSg9RBQAzyjVFBlb4G1o5r8pg4XM6yH
xIeX37cR4LADqJ60X/0LRhWOyHzYB22igHKHw1VtPdKqr9srXSw1ARcpsR6hVs84hAcVW7kxbUuK
iHyx1DRnHqqD55XF5qC01AH6SHPy5aDP0oVOjBmeLEukDzB9k0f9ptxvHNLfZHk5LhFJjLmN1EM/
Mi1c8B/eBfcDvEByQa9KmHHWWpKIAe9FVW45F+VhUA41GPG/REQaBvsqYay281JmSLXT/OABtGt+
tJ97MAD8kDRcPrJUoaVc+9efcqn587BzJI38w9h64v0jsIGNvuKno9f7VFTbkMFSZdgpC93TusLD
QPZc0X90F+0URI/MR45Tu1TCY3bnhX7ZQIidx9Nsp37sw4fEU7fNAJt4l5VnR2Nvn1to/KbU8eFy
b1RtPXNqJi64bsDZfc63qhEJi3Jt3tf4qkQbRNrt8CFdO/EGEgi/3op9vHJuP7Eof63Q+hcXxLpk
fAbR5BVCGUTgo+hfNu4yvl4BvVAUyS3hugTaJfAoRebgKZrT+wgOhlbdk9d8EMsd5/STdXI4pkjg
JFXYhu8ewp1YsRKwB4+7KxgeRl9fiKsBU7DSCmrNt8QsfJ3xIcXUV1S894Sdpqb7Viqx72FhqV7+
di6xy3wmzfjhamz94p9/lEk+wVzEK+gktriPiS2PlbbjY+KVVncM1O10tyYp1yMffY5bONhE7ozg
iMa1TXAV/SdTJlQV1sc5J1NsQu+HKIP/1IqVRn9Xt/SZYQ6bP7O27NxmiJ46JCYWCmeAc4g5bNV+
bhkifjVBDrc+Xw5GVfq5N3JhVEMizjcNes2Zp+Nh7ozolpSVVKWxMSFTQ20FYWXXgOc4H0rYdwKK
hxBYTuWiQ23mp1MfgghpFtB8hxBgIupAd18O7C/SfXGxNJGYLsr5BrZbSwCWbdlpjftvIdY2+DKu
1Sr92OGwPW26Lu5a1YNVGKHzYaBGj0FqPLRyhPKnvJkMlTe3VDyvAFe3hgEaqn0sGDJqUpj6Rs8B
u8WugIEjOW/7kIJ1mtcY6RMVdX/hTgpiq9QOrBRP44oBEGuhyCWl5EC9wBiqiFqnSRzurWTpaGz1
/hIDlCxLi1hhYiLMGeuSUqdSYt75HA7RAYsoSDtEg8bBsjLfXbZySkeeJvFaB+k+Tio5K65PBPYC
W3uiBxaNR6tl8+jBPiwPWR6u7eQolKYFaqbAfbcqDNEa1vmPmQ/zYR0/Yrzz0YoqH4Z1tuoTgaSH
0qRca/7krYFwZdGzWxlMuakdqji/xW6GSIxjPAPPp/HTSihnOwwc/QtraJI7eU/WgkFmNHx4leyK
1oTvMXo4LaWZlSPPo6EappWUYtJfHtVvOXL7mE2dBsopAP6KGIsDrigl0Ho89xWgKVEh5mTK4ZD4
wI7chI8jdFfY1E8r85Ow9xJGx3yOKuASHmLUinZ2iJP0C/hYCvIEv/kZYRedREu8Ui7exG9L9ST+
bSWlqHbkvEmGCVdq54GACP2RQWlvp/PpvnF8Ihabq+wRYvlpjLdWBjQ10RwpOpLj5SH2CGkquNxs
m56ubjSxTrnfGW22fM/vGt2ndz419kAmAKIGIzLX8BLLGNEA1z601jw63MakA4hjfG90IU17XCHb
/D2I69ILxysIU0eHu2C4MVP8KUpkN/s47k+s5lIGSiCazc4OrulWS+gDeXoYn0UU9WC2UP58WPSH
gil5lJSs6w8Uzu8DjGqJbbBxLjT78Xw/SatlaxS6bberwrIsF7RgDfRvKdmtfh2odL5GanFXg7u1
L3j61ckhjYDl047wCNyoKXpvjhop83nrNHuzyCRIu8r2y4ZTqFwgT3nH4t0js32pJo0tmDrAFU91
KJ80XVoTwnT9y73Y7hIdScUvmR0O8L0YnQ/Zwwutc5oD9F9Y1EZwcIs7yaC+0m0PfKTum47zqCWE
ieF1xMxK8+juqJIiBabT9dbsQbmBrEE7UfARlYJmwrwdoqXvhk2bf1BR6UqZH3TUbb8sUaV1MgFU
QG5UBWl7vKTAcxS3P+lRu1Vywjre5V+7KiFLG1SUd8jgvj6TUKEjnMLfZV8V8zCLpj8AHqe3N7gX
O9hwVjsqZJkWtWicctz6i1/YhJrQQX2lDu3QW/OixUTOSotok54plG4p6zpAs9fuVhAyuP7l69da
ne3aTbRQcfqkhoKZYWMN8eYE0x3g8fi1Q2rkHgoKK6+Xeae0FKvf5bRBa47Whnb5jTPHAEt42qIm
n8zfRB1NfKPxeXBQZahVQxEqKI59DV7RtR036ycAMiK+bsQLnbReHAWfuHZGMNPI+x/Cm5NSIY6I
7r9coau4gldAK1ot8kLrTf98tgpnld1K2d4BfK3HO20PX4p+4WUEtNoY3/5BGk9+H8uFV0SbWT+Z
rIofwHg9Fv8IZ6mxrERBytytNoj2pJcGB7CIzKxPrEqwK87Y1Q/KkivRforcWD7bW0t0WUwSA4FT
XsF+c9Fk7+16sG91hv2QCHT/5sVU2Mj3AdNQgppPXoVEWqUsXrfKaHW1N9hFvZYoRYt+TkdzvA+1
nwJfhMsrseaXfZ2/UjJ7jOq/wDli0bG+gADZvp1jSzjLvOMrR7AAwdtbtRUJFyA77sc+6CLmzWkr
uBpvsUp2CBEuCBw5to3Ac29byMy7G7M1lATZXkohwmLGgvt3WSpnbr9B9ASVGDoGkwlH6fY2o1IE
vMo7DeHH66/8JHqH6HWHbFs5+G/yOKZvIBg3ZimRgYFO4+bF8XNv4n9aIFvpRU/Z9EFa1FQ/xFTL
CwgvXKIq1uPLGCRUTUBTC0FlrM6pEFJQ4Ry1MLOvy+TwLybG3BUbYNE/qxxVfaVhP5T9pRr9k1du
9PUqlUp5vmgGUz35OUTBkQ0TFf6EzPrOkPCw+TkH5a2jTmYbUw7ZVZeqDY24PS2OaPN4cEuTK7fN
hyh7I8ZutAF4Ocox+HTbua+nYZ9lIO51rygDAvSqJ/GMdmdQpZ7AOh5ppqmDjfqrmUmQ5vvRk18Q
HbJnyBgDpoc8Nb6WnN//AuBiHNrTa1Bejjy1araXD5zAcNEdUvTz+Ls5G3RpjALANu92TwPH4yWO
B0bmHjEhihlQWb/ImUkcaq0kc2OSPRX5I2msJSAoYj7heLOI6A1ammPzjs+eCv68k/YGtcTLfgOT
n+zFq9wDM/J8KJP9sW1XNr8+fuL4m3jXfqcy8UQhn5ClkKTOiszd9mZ1KPWXu24+xj3j8AYrLrba
AnOlgfKw8m+1wNHX+VBi20fpadsknGAUcwSc69yep2KKW4Jt/koECOLpUtc+3Hr0IrFhxF89marU
4gxoBecBfL4AKVpM4kySRrRHK7LYeJBp/uPAR680040W25u42yru2w9BQb/7AbCHm6ZUCjdMUXvf
uj36sCjcs5WwvJxYCcgAh7dLnbNO5MOGHLrTn0gZFYoRyik63QxBei6TeH6fhxpfxBUt4ogrFXAV
ED84Wn9WF1qFsVv/bfzGufgBi9++KN0gSR4rX/UYPzQ+6KLQ6AHaTRjexVC2bMBKg2mgmEIFVuqZ
J9jnZb25lTsq+ECiGmWhL+UNk0J5ucdpI4dc7bsAgR8u4j5Ls2z2cZWW7fdGf0rjXInGBnTcja/I
S8+QViAX+CrwlIw/6baUS6IUx1IaLQUQjCNY7E8+h1cg5rwDXgMNs8t0v9Dgiromb4TZG7d3aAku
xepLlPUkck6zlLxc+zlvsApLXZmBlfTDoge9icy0D2Ax6mB7bsOCa39t6JRXXKvBrgAZjiUWTpMQ
bhwJBGvOTexasG6VLmQYLkW6BSm1oKwx1yLUhu/GDkBMgaez4UU5eCosS8HvPXXS54aKKW0kJNUD
fsKguTYTZYwDpEKdN8Wzy/pMOtbgNIQDftcBmSytYT3hp3KLozRpmESAbSYj0Os2Q2KrTYIoobGl
pZIieHqTf7skxckpssZhYuhZgxtIfivjzi9NznGjOa9+xGxIcu1c8E3lXWGni1EKh0vSQAIt5W1E
CxZipIUKYXv0ve9yumclnb4gHMvLcbHVc8B8NP5WICTz0xnUxdLavRehB/102ILXuf/C0miU+idL
ZbsJDPl33hvI4q0Bke49cOdfNS3RuQSU+T1jvtUAfVs2iGZtTfdZaEo3VrrX5Kdkn4l34Yi1axtf
kvsnE27T/M2QGUdbgDD08n3duvS7xG5NOeZEBLMBN3L0dQewTkYN8/q9PVdHm7ate4K92+3d1624
8zvUzzVxqZ/aP2cD0zSX7YEhWrO6Ogy7PSJMV90O3V6Zk+e75huFMWfZAgYw6TQJdCVrFseFcFT1
8OleXRGk81/SPcLByk8jqVbQB+HtZuzIPZWhY+pxlMVr7UzDrJjTqPM16p6iIn3EOyjw+4S2dbZs
gJz+onMXnTrTQJkU+LFcOWPL9riKEx8v2zDmNMQW6+XCJNVDYSXlN0BXSuDWfQ0ahSS0Y0dllNCV
leCXPctD5O4oLFjG+kTU8ZMZtGudTLSEQ2N7pYFl6KvZKc6bHihLDNuG4DOtgO4/0/3M3xEQyy/G
ikIfpSUAd5NoBcVJ2aFVr4y+ENUC7DMhIdkCCG1JDkVvYQeVozuX95ZZTUF1OL1MzU87CF4UyqH8
xew9x6ZWQI690oT3qKHiqAnP38k31rM9aEd/E+Qhbo9eTJGgT5+mvtkYo3xwSoP76w/cW+44eWTr
2rvPvFWZir5dRnZGfNTNWwp3NL5276qE2XxxLu1k1bdML/4Bd+7Sf32+a1quZA0rBAPASkzEA8h1
cWlwdifFondLx0GK8l/R48nlCwM0S4+DK5M1w6fFVgnwuUw+/wnR9r1FxxAscy7kOjWEwfDYaJbP
23nQRC0smAHdBcEjPvGzEarACS4uM3E747gyaFenJnXCv4qVZ0jeFZPAzcQWVsjWkPzx5B3L852y
STtBZz7lojXiCw2hFpyZO6m3MxO+uAgkHs+l2/WJSUDFwf4E1q05iIM5n+qIGaSg6aHtRBuBJyaw
T7f/M3YUnocqsoZomChNnfMp0uTgKHQdTJZUTmllNgaoH7MJVFO32nKd2Ref+2oSsiCaHWlAuUXX
GWnjMSU0JwritfaClhoARLLJezF+ES9GpgkGM5tqEA8x6iYSCgAAHZJi0W30cvtb+/Cay6SDGd5Y
63aD+dUskC3Z4bAUowJb3lOH+uAfMhZYS0b+Y5twhMiAGg7ncidi0NgXAR+cKOzlPmqN7he9xBLR
8c5U/TCYEWq+hgrcxwzWRlapS9s0e79cTWksvMyDQyBVWF6er6zobOMFizPZQMkupVV8Cn/aBkcA
PDs5kYfhJbAMy/q3Pr7z7oc5Yfuh5phqnmg2A9osv+xNTzUU6YfWrGujriURNG8CONHMrzAr49Xf
5wiJ4/B359uAdbcPXRO6I9lmHv7e8vjIvwNbcrqVEmXlnxcJJ0v5UoMUUI0ycZRUuBmKB2pfSxS0
5sqXH0QZRW7K+CiQ8OKr3A4un/bKX3Ie+yoJbduyG7OuTIPVJDMrsQkzeYj0U+x1TbiTqmSQ8jrl
AoQ6nk5EFydwwOQka6+t1FKsDOzDqDsRrrbUsit3p4mkPRM9ixsTFoScaAIz6KRlw//QmjDk+Ios
iqidczrhf67e6e8fnZERxW5xrTb6vtjxFzm3sXxy4BcDpYWlD7rQUSm0UHB1oP+HBD/mTM9lUB5P
Y6UM1qZ1j5o0nLlQPqzykVRRjyg2lXKZZF4/RqhRHpJcg1oL5TVhPWunqdt6j+qnXAIL0IQh8V4W
gy+d1M6MRLnIMNgmrDBw0a2rGdXu1XdqCrLFK4f9w83H7sJL7Trvms4pw+jjOizamBKTlF6q09kH
XwiWAEbKy/i0x527TCUV+/+V4cUmzCVnvYuclKzGKF6UZPJOZRHikkshc7ps/Ecztfg0NKRJFGE5
cWZirQ2lp5Ib3L6mZMO2ViAyxFMPR1894AD7beB6hki4XbNtLf5cQQ7+cZmMwGhPj8hz9lnNde8Z
U+uaY8S3Fb8Fq3KcgUalxtMLPZT3e5tBWMiNiDLEzKia/TdQ20WzVsbGc3yyLyezJtTmFOvlfBDv
BRh7q5CGWL7U9OQzYIVgqO7ee/9IjOsTlw7aJ5j9VUVu5TIY1+aQbHP8IqKuW1taYk54k09kxoGC
om2M4pc9C/7zn3qKS9PbuwTMO7fRWhgG+WeH+bWRwsNtIGy2AB+D3pLadqenHiBg3y2a7rfnf/Qw
HRRvXrOZttTRD3lOAmMe8hc/7Z/PNq52iikUm08JmxnKZsgtO9hswDR8UIYzoRFuiQi7jAalnKcd
HMcbAFz+YUovVsERuS08kjeqegHjy29yJNNTnu1+2AfqcdtPeCvoUbK1nFt35jEj0GZwAi3ZflaY
SJ9dqZmMrIJ2yO/TRneEl1SZeGHMmbAsoEXXiGhOX4LKag2vnVnvngCB2NuA0b2n3/fWYu/bd9+9
NgasIeUY0lUrORVEXD56p4ez3hxiB2XogLZgkRRONgiKxLeB/1hzHv1US/kGGodyfaAJh1iDIJbc
8Hn19I4Jn9FFud7clUrToaiEWV4rpmsLx9w3lgkVYYLxFR5QrRnhmKF4ktI2cEhnzJe+GSg18xl1
eYCJgG8OHhKq4PxRaZ5v5RL9iYjWm4MPLXf0+k0Ol6b8ouH8p4s96iLRM+E4PDAciDq/lK/SEg8N
JfoQtNCRwFmPTZXWEowspGg2d/S+2malirTVLxfQ2k6DqFQspeenhjgVbN349GFrNkH4x14LK8Wa
GaIB7Heb/UuKCrJj3LZT2UV3/ubT7T0cX7gSNQCV/+Tu0S6KoDSa6YJn71fM1LPogwAVeWaFGTy8
fBnEVzAgtfZo+lIF0YrLYPNylfgdLHm/+Mq8EyJLxEffAdGUF1Aaud4tybaGppRnFgtLzAQRDhfj
pyITplC6K8mqgFBPtuooE9c4LBW6WymYvx31RLcX99ncfeEL0lPMpP09TQiH7maVGT41elZYP02l
xLo8R1FndXEgBcyrDCtpCoLufjo/8/gBl4oDcUpPALnwGuQZtl38BVf2kmdf4By9lALb3m6bK411
Y2oY+DncRDciAusMJ01W6jv787ZZ31q9qGsjgo4LqrD/b8Fd0wTzMnKjFXhZh9wnUWow0eB4K83D
0IVYA/cLUKJcA/8itCf/WisbbiW/BscvZonysWaxbW7zkQw4pVKNtq49xwF8lRNhfXxIS6ANf0Gu
1H8oQvNX6uqAlhEd0CzKYrcEa+QRahicCGzSMGu6y2h6VLvpNEhKrYU6fdg7NflRLwU3Ci4tuV4v
iK0SRP0ctgC2rVa+xWMxg0hYXQ5zKGaUB+QfOSrURDlQO2i0nKikWAxHNSO1JJcWPj1jZ8r5bw9e
XetWacn6AQcx6SIpQNwMtCR/scZRQd6ti1g9V8kl1rWSubqTBeXWYNhcdPxP70v+bjmHGOYSZBFA
p9vZA0lrh8zVF+wmnB93XRppLlwtgj9RUBGunuPhJQOJ9V8THx0gr1jRq1zdolK8uRWYtqOX7WKi
fnDVQNpLBcK1F6QwssOxNd+oEnMizqeJyIaz6Rnxh1ZTqrVjn1KtDdT63aHlINSLFgo8YLN19/kD
ohwXYyEetNADOfKZZCvj6ORSJMZCdXHxvtksjrGxWjjTnOKeDS4fA7CSDBzFs9TgFK2uBF4+pCAa
RQqiRXxSp+ymwOdgE1cvVSSqUwuYxw48YuiQTlhWLFKdAfHmLaXVpdFKYnRn4v4qHvu5f/+kvTwV
xirGD9vY6/9HMRU6+AJP4RcwCX910ZncRgXkwcdrtGVzQaVRbgg0GnWaQU/ANAaq3K+Z4+X8rCBl
DluKjczbRRoK81/8KG8Q8Cf2cJ5kKUOYtE5kGUBZ+H0B7UsvGHBmfOhCgrdjfmn+D2W8EGwrTXyJ
fxyMhJHffvLV7C54YlqzG0UUQMF2MLkwsv5LA2Bb5RfWbyFpOPyBbe5QFtV17HCui8dM411eGpNe
q5e1ofErX8hV9wJUv+YngtEDc2E0qPtnuv5SzM7e0CtV605NJMmPuxXRm9eOuRuijSkjn3LA4KHy
5fU8Vh7yackROYj7CoOqD1pxcYA4B/dRERhHsR2noNN4JfoLTQBDTBZfdiK0jp/fxB7TEPdoIT1W
rfw/jCaY6mwqULD3bVtrfEI8DrglahmbyrY2r002d8WiihUE02ZLMAL/X5aFc7ohvmOQX1/tjBtG
V3lKL3atSsJDRs5r0nhNCkIT/8FYNG8couVjrC68MjykHf36Zot/e1Y9mprWY5k5fCRGjKGrro/E
dmmCyOITS/qYwM1drxIfC2aI5CBDGDEliNiQMs5V1Dn4TicWZkqYmIPhFRAj3FiKRmvJl9lkYhkV
fwA4xquoZZkFA1Z1YZZQO9j4NPVOjldnhX1dydnV8asEjQ7XpXsw4GoSljS6USCs5VY02jUoJv8Z
7jTQw1+yD9nf0Kbul4UOMOz3RCij8TMZpqYmfjpATeVLiW2WVL6a4yqj0Jz/TB+lLuLGhzZUHDbh
H7Q6oDrH3mI1QiU89oLtVNMbHyJFWIU4sTIE+lpKwy3vgVLorqtjeMwcKqxS8KyJfV0cCiHuNVER
yy0buEKOfueH4EXVWMT72XEqn4M9mjp6yxnKqIJBqdDrMfVZQoEJfcNdPWPfuWHRNskDMlt8YFyw
rMqSSl2iPUZ13MobpCnO8+pTXwNNXLckFlTDVARS2ClD3c4Y85TqRrTZi8LMWI+2n0GuuXvP6RFd
+pcsGwKZ5tERF3e0iCKwTRAGUODbiFoMtdl0AiqN281bIHXZHadVx/T2DEDmHLyiSoArBV9SvjtU
UrpwZw/4QSDdG4+y3Fjm+vTpq+i5JcWnrhGroOt2Dk/7r46B7n1XZj6lQbyaNiIP/D+vxgDQa4QY
e3SvRG4BMMGsRrwa2e5lU78wJU3V4mCNWvr6+J3XJx+NJVEb3Iln9x6tuV1am3tibZZUkl5xhuZk
1j66wQhEOXfXqC87NfuKFmZEHb7JTmJNIhceL5G6PJb1B6CdtdrHKKxsVeBRjubnbWIOQBOsGQhR
AvK0K1pw72V7vcQUP82OhpVrt4F4LpRzZwpgMm4D2OzEuaq4FIx50TERttzm/ZabjWZTBLYgGtsu
mhej6Qc0JVYWsWexHocmEUFAGEhYKThepYnFxVQP78k9rN6MAD7Pnx6JY2OocV4Q6bmTnh1Qug28
lbDdJQNpbqDbCq8C+eZokWnxkrhgkvvmlPQBjABTSbEmulaPYGxTFDdECJfhkQbTlEWwd9lT9oIv
dI6/ShVCeGecF8KmRKcdYiB0sJGwVGIJgBURyg4YWhSjQI/AT/giL8dTpZ3DU4+nh6UKBKHxMb8N
WWPvbQ04FFtbDXIv61nYZUuf9eWLr68i62NH2g34j8d8AVsmNqRSERE2rukiOr19eLRsgpcRI+t7
b6DEcIn1wg/BrTr2gs7uCvQZFyj8D7yLYKZHk8OrJaavqo338KSIb2g79U4+8jHxlrh24Mwysgb1
kmpzd/xO3qo8WrMZFIougAER31MlZ8CZ3pyC83z0KzCEUnA0aX7v1fXG+E12cGZtsG1Err0VXDTL
vYlPmM/SVoWMoQYQegLl2kkh/hPMETXYxj11pLTJXWGorkYpUEkSyG5bOVUR1xHODPwFMvieeqPJ
B2EIwJXmi+rjU6jGd8WHWL/SW434qto39oDNZSTCslrPikeJyO9yZAXAiGGSjBsX5AqnkzHeN+sF
pkaVDT8AXzjJpvCKX7l5x0A2fsq2XE0kRi7SsqaSdjMinapU8AScn5jTlUaZUons0tQ8H40IisAO
PmcWNnSVwJTp3vR5KJv/J6uvnFMQe7d75vK9dgooZyUcmFnSXyCwmnddYIClzkX3SGEkk8E0g9qu
ZWmadKf7Y2zvIx39cfOjarf5tWRyzK3mrBoyiZxeJNLuEywo4TeyWYvgYia2Y9A5Tiwy3Xb6fKfD
1wuMd1MDXaArwLP18xoL0xzbgqrwQZK/mR9Sxx+8eJh39XBmQfHIq2XmS+2WLFoJHM1VbVqg261N
Rx9cuRgFcEjU9CdwhZ1j/kmv2KXF5liW/zG+n+36eWM9gezTw5EMRUCNjv0zv5gfbl2iBYb0+kAq
m1bXi6mUbZvUV/xDDxp0WvbTsW2yHeecPkaataKLAANa0+gxImAn1pNe25uOSn8ZHs4W6i9ltLAe
X7+enqr4RTRBC+kULHJjAL21xPFhmezdEfgM9b8Zp3tKD5NZdkZeVpH33Lj8yUW8ZYAsac8cEgQ7
1QiPBpiFh1nrxGrNPCZ+5K+4gblwC20689za5T8v3z6cGVJ3mdrxKt9Ny1NjwlSKyySqBqZ1pzVO
aq8cUSp3qQki2P2bNrRh5ugZh8cxGfV7C0Fqv+KaYNjrC8naSYbJSm4r2qL4V4iQ52d2Ts2reHjq
Y7O3lsgg09awgAb9NUfh5BLCBI47YE4sZjpwZs9PHchKlBqryMvFYzUAKXIrqukot7WKNJz7XXtZ
T9hh1uNYvAXj5nfEV84sOhLx8Q7JVjzvHiWH37pRQ0c3WdJxfMEko5anVNNv4LO/eISwL8iSaajj
NQNAzl0KfrGOpdHvbeI6maOwu220uH26411B39ekv+px1tM/Iey9JQqEBPM4X1TLqqPrL5DHXVQy
ZhUTvWWVwUo6WouQkf9P39MyxoSSKjqLXnd013aFfhOtri/cER+5YU837Dfr67NeD2hvGLLp0hif
SnNNGqvHHA8q81E0e6naIOXlm3JbuXP1vGeeou9RtNeINmJy9cGKDTTPtTYlh1LXk4dB498S2Aul
dNKybhZR94prAbTkn67tz1PFKIxkVpM574kyI0zSUQeaVnTOwY+XrpdzrkfGhKWKmsF25wEG3I6N
LZWvWDX6ljJBSOWan//DZuTH9JRJ8qzbRUAb81bkMqJbEeam/9L7QM3OReuM10cR9FzhcdUMdOjX
z4gKpksmGYMPDI4mpOA1X3RJ+KABJiwUfxXFPsKARrMERoE0PYHIEwMN3lPoiBAwYN3UeJHmLPx4
PKZAbIWPpSnda/ePbAUe4eEiu3X07uZMHc4vbwdEcMKaWM3SoHZp7yF3tRxAXOjAggKYsPABsBBP
984+wG6bNprBAA8xALxkbVk/QN1c513jcY9M31OK8puUPyLBDixxamDlIXDe5pTnL7YLUuhb3yWU
0VWOAp0R1wi1w1ardbMOcQNm8onmwEtp/PIB7/rYlFuKvre4aG3zfGDaXA1jC9IReJgV9XDwflGK
LfWU/cxs5xl096Q+Vhz5PksxvH7eeW6xdLnA7rkhHmGj1Ie3ZeTn+obXK7aFuhegd0lu3Yx5Wzic
hJxfnAf+qL9LDZn6P5bkOATd4RUDCN3AukxndtvgvGXG6uiG+j2ypW+oQN6wxvXj7k49WPw5H8Qx
LYWRSjXK5CNfdGkGBf34s8EIELF/osaEilKM+DY+nYKU3RrSKRH0otEw4eDbUvAR6qr+7rRrbwie
NqUM1VQMnNtMF3A0sGwS//lo2Bh10esGZhe6X4C0P23NxGcGHzjcL73KWtsiKUNK3/cpfCT8xuyI
nZhTR+LUDGEQNTL+cPi4ITzmtt5Ae4ogqg0zMoUoh+Rt4xKekK/+b5GMIu005S7BOD0VBe3I/jxZ
QRfwa70o3Y/8GzpzDr7o3LJJE8yAF92V4rFfg/BF4wGqWgYNLDO4l8/6uA2tECgYnYg2lqk19Bnk
9cgegPJeeB/Gh/QtnKkU8C8EWKAOGNEF2QSahN8tCAkQxKALzgdH5cTQPU0bl+NO/RDXATKyAR8i
/eG+jzu+Hw7SBOPAZyqmHiSZqkJPwcg9unwxcCIyaJd5fq6FQ/Y3u5iyGNv/rVBaf4WN+sly4oUn
V6nBI1qmN1IPez0SVmS7PXlg79SlJwuaayAauCAmryRaCp7bpK9VzsKKBVUr1cckKrS5O5TpsegL
Wh1/IlyXFFSzyL7v52ecTDUAOWzbNF9TFRMjx1dA0fMvvrzFz9uEvsF9IwaMP/vuGAV03Jtd6LTj
R48D3v/Un1ByNZ5LQSsu53cnlcWHrw4SiVHSPjbYoRV41J8ZjwgsrxqUGnDqEvYgILRwYUH7Bdew
SOC044yJfZVqZDS+q5ED2Opp2nvFQV9sSshVyT2l0im0v0JQXK248iMKNOrgi12o5IBiysN2mpnT
+jiCAjdm2YK4xkeoITl+rz1sxA2CcNTVToNZ3hm/8zMkAG7gIOSYurlpuX6JfMmdlAAb0tkKjmsa
EymCweBWoF3Qfw+3wmkCB05hCRlnVOzk+V3G8HsLxq2XdTH2jNTKFkmAf2WEuwGomWr00/oQBFiU
UxtywHwrXHlWu+2TwTeRqDeH5K0TxLmSbdfl0KKja0hC8sEXCHXxtyko8gGEu9xSNPe7CqloKhh5
KU+x6aySBw0N4Mqjb6dhZPxz6+Hn8aV24bLbKoPEsfSMjyn3za5knwVs23Dd5cavjXZCvPlKfL+b
61XBMe5Y6Q5m0mkBiKs9WHOIbPFtRWWzTfrecIjingL6YcjaqJy3KjAI9xO8SdDjutcAkCjIMx/Q
njARFOYbqK22b5AeaFGe4ROlkDRMJgeWSCCv8n251t2+/JYcET0KRU7lqRoubj1dnjgnEauoFDwi
qYvWrGr281tXrrqQqSEKzWBRBlTuM75SU/T4l3YCbWYzJdF+1I/C/0i2B7kohtJCHQNHhTrnCn2Z
4deqrn62zJtBdT/H7izsftjrgzjbpw/B2HUKR0WvqwuLGH8Sy4+YmJa5+kOlC/nHIiRp/MBTmRPn
xpldrL7i1LBgIydIY/4JOjvosP9M/ZFlC9T/tjGyfl2KN0HDN2dlSIq4ZMdcOrbVLwgHENj9KAmG
FqeWUEssekKp9Hy1PY0eRbthdsJ8oJLonZo7F1xshFiO5Ga/HzrkCcqt0i6DOH9kMAtneVagN9TO
29UAr6zvCZ/t0t/pDPcgMFSN29Nb/1U4E/ljGMwA6oQpRUTjv2X3W6Ay8rmVUoICrnwS3UznMpkK
I+4+njzFaUcnDbLd1PFXYi4MXnVH588DZrcaSpisvxe4YNjx7eW5vqX2ffAfzp3sPYPCCKvWzWAa
DtE55qNJ+5F3162lzKivjEeLkO5K9f+tk1fiaoyO4aICwPYaAxU8abqQ6uFdhkQOZyRkxVpGetPJ
JMQZHH1SfKJqH5NVyDsqLZ+VU8aiy1ojgIS0ccTKe8ORctsyIaoMmzt40L25+MfWLRKgCSRtCjBe
EChPQY8bb0mhb/fhjPixSIFfrZmFMEozUBzBQGyoD8dezndQsSb8IKrZMMDdvJTZ0f5/KZF3zHz4
3/uMq+GObtX89QWnIl/i4G2l049DMKz4jwmZY8+sHr37krlJIeILlbdNH5MQg3bZK9luAUxi7GiE
5imPQpH4YGNk9baRqKaIrMGStJ2SjWM8dpL+A9qHxe6kdsbt1yKNnEThY37r0Rd0+V4qO8RrWrdn
hUzPPR00PZUBlFignWpkFb08oakopTHLSDf8heGdyA/i068bZJRTIzWXwu4t6nkHX+ED5/n2Iu/n
SjKrqt1sakD65NUhS3JEk1bQo7kwGm7PgIaxxF8CZ+7/hoPKgRFsA0QTGb6j3F460Uf8grMcYIvy
cXccPlv8UWu1mkP4eN85+dMO6RTMmnTX4Zl2Sg6wXV9qD1y9Kg61/aeIzKNQoUrn7QzJ58NyVMVT
kf5A1KoHCpWIswb0n/8UZBtTr2vMNQEfaR9TeRUsTkghoDimCnhMmepMx9GQkviscp+XaZrvv941
6g7qR/5WGqxsNNrZ64LwXexKLPHILt+032l5IMJBDJtfcNY+e5D1HR+wvsHr5yS51+l5ZxaVlSFp
oBvvOO9agGahpyGInq5i9wrmiREbMdj6Ox/vcANTaLGXwkEK9Q1K2o9J63eSFMat23/iwBTYl7it
uyQRKBW0VoiDNSVgPNzdJ2Hpybe3vvwHkme1teCzFnz7er7y3aH6Nu01rp43NWwd5ug29k+mxc2l
omB0XYnzAme18MKzZFlrHwM7Ab0wuKBIpaVX+7rUlH84WxkMEI+WwnZpt1sLCq4l84Y9s35QYY6w
+dNl+SIhyS67wnAjyqm8gXFkuXFRkfoz9Slp32z5hBBwBoLHv43wYyRH6wkNaeckeme/LJtNRN3v
ofjTTUYLJ+Shorr/gJe51KbpCOFaL1RzdqT7knpXOOfoynpHUxtINfEJR/ZM9mrwLMr9JkYKinou
SiF+sXG92AELXoZaP/bRfoEf6C/mkUH+/QZrx0NwnfvafspgAH+XWfZ4YXuPddKHHWkYPQtZEkCw
9rCjx2WaMo2I9+qnEkvPW7U4xEmp+MDSwM05zRRd1wSdN190fRJANGZsVsyLCrc9V87Cwns1+Sny
9ChAqemk3E3bRt3RhhRa5l7MI4nw4FldWzjKhG/Ts5Y5oavholdZzd2SGMmEYbjYyQ0XKLUhwv6K
GRJ02NxmErl5rE/mBQ0PlMkhL3Xg1ZKJ6RB0bzHpXqFmYdyJspBs7LeNwUxor9u1g6WFcIyXHEep
zPmmgq5dKKzS8X0qa5KOMJADMb3oDEhRVwEpEgDu1R33j3Q7KRu9dvGPoG06/zpP6GeQssnjLsVR
/UvLOoVR1TQBOJ+UVGTbyRHbo8iWy9vDtD/dOUWsixIW26mAvwgHiIk3abkFJgAtPd80JY8fjNqo
xzZ+cLJ4zM27F70nUtOATFG5s0omF7mwp/mP6jgpan3qGmUA46P0w/Kh4YIqNBqbUmTMczDv6Wzz
Epp4qHEfnUBsctfupRrmbNa1Uq6W9EWLpLDIE40+Fr5iesKUUs/fiX1SuuEIFSxHgT5tAjFQbCNx
bDhGib5XJ2ecKgwY2MGZuLt7dW7JQiYf2tBumzFrtK9wwscX5RKAIpE1h6w9TbMt2Q5Y+x5ecq2R
adR0BmsJMBERRPz3BQ/9U4GDX0YmuI/Q8khooinwpuiFMJXPHCdXvlB1jHvF/wFkEzfzM+FpC+Zp
Hm56Z+FVqmGWiigLuBImFJZlro7GluOrdcwJ3s6VMqCyQYtK92XMq3TFQ5fwPuJM8Mhcj9Mh0Ist
iDNI69fQeRjxHkDVtslVhkQHP00f8BfICWkRn+kpsS/uqOFPI9hRW9gOqg+Y4ryhvwOsjqBQUI1T
05IegyFOuGs3Wu9eayeVcRLQZWDTTu3hLSLLFxBEJAt1hp4uUhnejc57HCSt8/hQAnWVxTufSLAA
S1TULEC7o009dVoPmAqW71qsUDW4ErZ1p6KWL4NxLaKg/wXE/0voj8cvAdXFipPfmRsL2IV/4kVs
qLQeG/2VkzGIXQYnHWUoaQd82Ub8gHBGUfacROrRhGAwmRm3maUvBjtN44QgyLlynzhm87wkG7hn
MYFjPZ5t8B8vGDi7nswd9PTrLQbeWx06hBRxdup8oBGKR6cs0TZTKdwn7oIxPF0YE+5mD8+6I1vm
C/Osxfwx5o7t4DdEY49KAa6QEYDdvsl85UJXXLUnKCV10w0GmxoWGX/JDzaaZhuwAgg2I9bBGUcw
QR7DBpS0gfPLXSz2rXVJcOa/BzyvZMFcxQBb5KK0z8PxpCJdYojZwdDBdF0kB1+asXk3zeDgYkat
T3wwo/6C/RSI9iV00CEAfYl4HowOB/qQyJoqFQFpEq/wRTnrZk2+llnTJ2SN2Vm57MA/i+75VIdX
kvfof+B139SDIP/Hn2KC021wp31rpH+MgbIeI207DIfoKNrElzP60EGEHpOWVt6ljB582gMs+YNT
67H2xrkocIgHmC3/FNn23e+YAywD9heui9TwsNwbaNcSty7EqkL8PmCQrGgv3wEjoiKHQ6dqeOAP
f0SH98U5AyqjwoPDIHU1ZMGonO45sTYOJ3wZH994K30Z+APR2yZJtrrd5nm/Sy9vyutxUtBRov5j
dqyvSNfyzdApyN75qipzvj2e5dSn9Fg/taLoN5zgtTxyQxs9Lvjl+sbbubxlQq0rdIJ+uuQNq+Sq
xGuzuyfiFnYDxgW/Vdhx9gbUl6r/fo7viprzkskrWoTonsqsYZ107fZ09aWTp2zYEhmXUOPHeRv5
5KlKdXJ36lvC27bj98yQp8e69i9cvuYXBBClzCDQJcWFq42HEtEsiFhEDygDvQwGF9o767gpsMHk
ZHMO3+paIP+sR5DT18dFPEjkGbliCdfndsFFVtFlx0sEMQEVSXwOHbBSij8mztGOXtTXQuj+aJYj
qkN4dWxg/4HpadQ5XGZbPnT98DSWiT1AUD1rD754cOdG0jwCw5o2UB4crEUXaCZ3tEWbuuIWK5gD
QDantlIFwY9kgMRr4LtXmEw124SCZgvlXkgbcwz8tIjSxc+xrqsxLUBn8GqkdQRvvOxRJwodaHvh
V6BvY0+YSBinVEUXTt5SON8jxd9+Hu0MAwPck9wztD6eFA1+azPxAX++vG+vG+fu2nUOxrf1F8aS
qEmfdQ14NNRK3vp4H8avAZ1nLYSDQspppQdS9rbA9oI9Okyx154AA3MPGKKD/BoIEbaUPHk6tTLc
Lym5WSIFo23keV+WIUcPjt64jHx3SnU2hkgBkQ3j4xZ0LhVNQCnSlUcXI41fo/abi61RCSVkOEEg
A44rSkCqP+iTO+RgrvwTIWQYejgRKWYE4UMwGqTZsoZnFSU5JleQLTfR24BG2cCJ6HlLRBGvdju4
xIHi7ffjCtCFqpXFFgowDFG7fHN7WUEXcTwhi6CssnClsELnMEwcyWKk3qlm8rM11a9qRPBNBHnv
OmsWbsL4Ltj7KFRW4rF6fqzBJmf32A1M1XsVwIQuu9ZTkV+nck2bD232zFIVQd3XDpsd+GDLk14E
X0HLmh98wwPqpDztBX+fZV1Uo9O1VmpEYlSeWqLnoibYNFG0ezv/qNNdAUT6KLhkBjZMdweCy/im
2STliucJRjeCaGlTKWJgvLPGOFdSeFcbw1DbT0Ff5s+p5fuAghjyh2bIXtsN/24FNrTQWNtRALqo
bnONR6gHVHEFtM4PYBcMUDfRHngQ7HIhbrAm9/u7NW/BX9wGt1YNZ1LqGTjpHouP55NRNsiqPGQ6
U3oUecEVbWGh0LlnwoiM8h943byuMUq7GDb2L4JNVa0bnzv2cfwupZWLboQmjrJ3pJ0r4hMlfJ2r
oDbXSUXLtmIhrM392E+MFZKtE5vc7Vxafr5i95+mIIcVpTk2xt3xG4jBXoK02GzmogjrqJappEKZ
p1tq2dp4VKQYR7gNR9DL3ygSqYd9JMsKzXtslyJnc3d0Ra8DXA6qO7Bjl+GFYvM9KRNwN7dxjpUq
o1xOVshTCKB4FMSjsku/EO+fXf3Zy57lC+lss4cqYz6ZuuND52oC5CwXa6L/SkkYb4stBUGDeZRM
+cKpFxho7NZ+7Sl2OPZj+/WAWCppQIIOV8p909avt49X0IVrx+RJeCkWenm5kjym6HLD9pU5pbkx
02fwMQ18KFKmdSkN2OKzIlkltDcqbaEnD7SdRUjTXRUWtJtr21MzZGNftkVdjxf4LPNIy/3g37WM
vzXUHi6nPlPTNLq8EDfhfT6mmgk84EUCSngEPoI93uY1vBNI1Inr37J19dMJ6UbM9V/KnGic4OMo
qHDhSpSCoYl5Hykvh8YXuGmzuJgtrT3eSJw15cKOOztzpT8KG+Zcg9ECdIocyDrDj8cFnL9VmTV+
Da5msWbn5rCPD0/GBrFimEBsI7P7E0SflkkVk9XSv2quuIC4XlmpT5+efsR0NoTHhCB1CGcuCC5y
70Q/sgWpELRXWExgpFxRLzvg8kPlDHAsv+LMTHPpF4eN40wY8jnWWrz6fHdCTPj4gIpI+qzhRkx+
ZxdyC05xAVXsP4NInOpHo7OS8g75hen0z+fadUvvSqA3gyock/vRDRaq/iWwZYMRX3qdmyhsDjs4
VmYp4FE80u1jDkafS2Mox8gQ+hLnUiFQTxAAVa6kaCxGu7Lbxu3kUG5o5AX5lv+7GvdH0SGGnbdh
bdLjsBQhsd9pSeXz9XIxPsJ6EhpVYVNQ/izsdbzlFlcXEm9FeoSdVuywgd/wmEiSod/+AcrU7rMt
UL5M7quXVdmFxj5Q6G4WLa8/MwYJNDHCPFHdbVLcXKWRLqA1vHzVLoIgpwc6Tk7fYnCgN6hDPo6z
7EpnhE+BtSvuinq9Y9sJgRgc8DURF9CtDFwWJ2VvgMplLxpNX2h/H6rkWpl/QnOrutAuCS47pZRA
YeRhhjiqevr2RG+z4Wtip3R9HRqNa8leC/6Ae3KXMzJAR0V/fGtcs7q5snuwhfCAU9NM7cYIgmE2
8Vh3IOpivo0cKd81IVNdlyiv8htlqkwL2geeB+bp86+6wo0/B4icb3wUXWXfK9tuWy4qwt/HynXX
8MsPSsDG+w24pT52uljjNsFCp/dtlkykE0OPtv/k39wDZsKLYqk99o/0EURav+6K5yLTV0yOu57h
eZH1pkHpRmm5LxL/8/GWKT18v7RBEpO94phrjNbifzWPJ7UWxB4COe0gOCwEUHnBNUXJGsoL47Rj
7BVUK6kUY0Ir6B9FU+3wR7jKkz4GJRCcXl4iPFMqqmFfzRm2W/QL1VuHTBXy46zPquTuVZJZn03G
KCCmNlY+Mk3s5I6S6FpRU9JSmzEe2kyWMBZi7Y+BRgPA9O8l0b03uZT38aUcp4Eku6Fcu2igCeOq
7XqPMhDLiJeVUJJEjf3xHRyY9jLUD90aKIMTaig3JxGgmfxHQp6o0II2kKVTmJ0a7e++h0XT7RvM
wJRhF3SXS2eyfj35HbBYU9TBUnbZrBHf6GbHPUjYApUIVySMOWHavFusRPP5gfzVlw/SUArQp/Vc
jUTDKDt0E/uMvUrbDmhv9dcheXEjmFjr2bgsdIFtMirErPqQhNOwJinwKnRd5CJNZrsyJ9xwa/U1
MtHqi+zPlmvABfj41FLT1n/89wNH6GC/CAPcWBoB4C+/Zgmw+i460q0K/usMgfIx6ptPSiVPuRfO
OwPHktex6X/67PfwMnT0Gfd7Ylo6TQ+1R2X9ia+DlGc/SKZix4U25RHOM6HWijwMxxk+1S6KxPyK
rwEuKiDEwIydOpiPuP4RMXCTJNx7woX0dwdyh8JL+u/OhHvSYhvZ1HdvoPH1tqaHRyx2oeo/YgS5
g9VZpvDqMs47oJ/fM1PWjcp5kWofHRHqNuILbGQ9g9kGOi1BQvMCHPMdcmaSkglbWBZnrorqmgw5
rM9aKcdjLAdO9pBUd5I7hU2r8wkUiJFJONTLm2GTXtQu9Dy5lcNXAtkbW6FyLA1uKbs1v47sYYQ8
e7CvsB/zeFd2ez6Mw/M6T6Ihmufppz3oIGPze4iDyQZv5TRJM+4henf+LW/Tzg4FyS8ziw+LZWjD
X0w6bg8mZoDkPVu/Ft/X+iyh2DAFn6owVJSoxDT0rVjUy3SxxZeH//I34KoaXflnmic88vS4hLGW
28VdtUPkxhkO2XyG27bTSPhMSjKl0atpKq3tDJf3DWemZ8jzKbcL9T5IiFcVuLucld1qPR+d/oB5
ldnUbBxwEsPVMyIf2Sffg0cphXJIsF2c3WABB8ym8q89sKZI3NnYeCry+195mBW8RhdZ0w2CLALY
VHseDVPDkOk9QWfRXfpm4OlQhPe9BBBeffmPVz67xBqcbNFIbYSZgA+CNqUc2/ipPt5om7u5QIrE
JpYqxlvMRlqDNKv+eyl+UQOhGJJ3gLSigtwL4aGbSpNdp1/qquAJEcmMF9XAOmGkGB4vxc9TcdM0
wSkNh+SjFmURT+CThqndNw/YEy5UKIg/KrPbYsd9BVnnojQbx24yRI5+ddm2kxc7y2QU0IOEbZFT
XdHxSUlZsribsCDGnLZqFuD6hvQ48QSVygKkTID9TXpoXuXMMTfQeNOTvp929lLw4bmeLYaFxGEL
K1v9FEx7P3eSZjGOkBtBmyA/yUvSbpyA81P03yRiX0KUydSqkVlTr+8qIVIfE3/X+X0mJCCzCQtW
nlDLNgvMeTth8gVV/MpnCCYOXYj+pQ33xykKr1KSW19majB0+5eMoJL5hKnnM1xw++mGu3mF59nA
uaX97xqbXh9T0J/iUQou1/GQD1hjs1FMe580L3Rfhzv5Ssk27gC9iFj2SH7vl6ktwtMdJ4TPA0l9
yyHw9Zp63bpTm4sC48jEeZoZ9piGWXw92nDBN4TN/da9sqdtvz7n/bZYdHJGOp6nYs8AjM46ysTq
d3Bw9vRAkB1ehXe8etEsrNbpBF5ZI/sdOAShSE1bx5FYcYPyQm3Mcm9hY64bAyA3mxegGB3V4Yx5
YVRh1J/Kacnp154xqgiJb4LEsz9lLw8yQ9WpP7MUmg9F8P24NBHdGJ4SteDsTkyiADLeBMFc/gDH
jgIFXeFjncoHx+vqh8Rkk9XXYvYyVoO13eFbhlksI1VahozgCVDxPyZwVT33MBufdFwgQgYIME3r
SVlxU0MdycE3R5J/eUZ5EACVBuMEyKuaR6ZrQy0LipLk1chmuCvrFC5qSdl+dVUC/PDUF8C/qzK1
wWw65omyrcO7W1dAQ9Fm/LFmzRe/IPkvUvgKOAO248jrqdPOcAlytGtl9b0AcD6jNOo3MH6GerkI
NS2i+8GXxg2HGOwHq231VLHHhuZ31AQuhCfT4wCGJw3bianHE4VOyN0nEIDNn2mqS8ylBqqbJVrb
TyIbT81WhQCxEh8OJ+N5a/W2ZiFN40KSySkl9sXn8XNfe4UvQYNp6o8faXtzNOFulPbaQDgSy7aw
eQFei+mIQmpxjTr2z0bJ6vY2VPHTRmB/sCCia4GjIZIgkeZGiabAS150sj3O/t1KynSeNfiTcd6M
625mim2umPLybxbglub/lZRn290720+7fcKscw7kCmH6ij1rvFlcaxPjaDAULw6IlAJmTY2Hk4h5
ElsVsJmJx5rvsFy3QlEshe0QfG+g+txIOSFm5M9soGyP4sxmCJSczu8X9bVesi8s3OrPHNzCIdts
3/2w265vIoUxxd4gl+1Bm0Yu5eoTdBEvvokSSLKRucOzwctuheLkrdkWbOUsXHJTA/UqtcnASoVX
nkNJyWYJ2MdkJHnIbvz8otz+XM/wen9T3KrfU3uLifeQb0tLWe0Ah21qkruPwxkTwvXZYhgKunec
hmyBm1Y/zATqw1xiIrt21qTASie7tcracCrwj+GgGNOIaQqvLtiyVZRUq8MOq+cypxGuvX+z2DrU
cwSgPlQm/7MgkhGqoqFaZSlauHbxk24B9TcuC1+V3UYqKRYpZkVu/pbNuIaq+IkhoP/Zr2FBPcaY
+pIwf3L4OllQvw7zIncDiKlHhTJZ9jwl88vFsIrefDODTNfiFLGIsLcT20MKG0bgTd+GhoHSl3tC
htH73tRbzI9HRqm39u8ozlMg61r252Z1XUhQ6XdA/jBGjySrwsU72dWYiQ3omQuC7wdaf0PS6hno
939K0pE2cxaGFU9qvcud+a7ks+gzmfgMiJjWm+rEgVgE38AiMHgshUfyxmAdB2GkpaoJm0rBbfdd
GxVHjBGywcInxycXjzIJdFi/11Xw1/hy1HaoGNDLqNLjv3Pd7g4mc757FEkwIdy6So6Vh5CXzoPL
vKrCkc6Fz6FsV85NhX8xqRaw1Alz4PIfbC4Ym8xCR0vnT+SFJTwFwp/mQ5inpGfxpHXUL8Nziu1A
pcqPjvWTrGypfAsGJYNCgbUISEcoLs87EZOCHtxS9Mg8YUgJ46dXLfKG9iQBtCe+2X0aMPhUG3RV
nlUm9dGifFYzR7czeismyreZoAmkPphe3VHb/svwuQs64nyIT2QOTJvyzL6Z+oVJkmxYDCtE+SUc
Vqra6nq4qFu/6sVbwO2vpbzMlQs1Z4x2M8GL+BAajqOAcVNWsY+7KVASyWLiWPJPhaozkUnHh8ck
lti+6quXhH++q0J5tZDx1Uf8qTZF608HhEiBGzmksRFPnNg0ViVcs8kZfZbSvEcXXxhtTwE+kWyZ
wmFJ/g8RkyXjxFgJxBSbH/g+iq2xXKtwKPWN3T00pRXuXBPSEX7IvkKfvNkxHirpBxDbQYjEa04o
bmAbEtYD0X/Oy6o9ABr86YUoht1+2mvlUVDmT/bJwPttUBZ1N3nBGwlzSwXOR26l3sYDQWvFMvjq
7YQ+thJfYkOJrtvAXSswC+WjcvB3wz5jKxYt1AHGMsg4mB04UIl53zxA5k/mX+RF2qyAwjtqCxMc
oEMBfMlE8E2zZtaqxDjjcEjFF+33O6bRPaB8pzTeI+V72ue+YdB3Za5xNe6U5VdmilgWRLmmBF9n
MVj2GPmNI1AG/C2ZxBKZYnWRYKdp96Dj4fn2fc4vGXmC9LW8uRJ6tBd2FAehw/87hce6oqi+HL0X
NBb3y4N+Y06NMDu1Ls33dXvsqsns5LjkjwiouSLLCf9nV9W2ZhfjiLkg0UZxk3czt+Y/0xnizcxt
dYxoeO86j5BUZMDa4R8I/7WykbEU6GZl2PferOIWc5UbEC78U6LgWREGQFCDgyTM6JmTD7wAe670
LNIE37Sb17E1UE87M78YC3RpZkv0+/sA4l2koQmBm8hgYFWHtFLFJIbS7TNQOibAMMCas9GczuzM
lZ23Bp9gy1bUQtXWZzb0oA2pF44W6xBJgQQlVGzxCtRP7HvTlZLnGiBa+8rksyPOMt918L4c7mc8
LEjWJSCRv/QFe+ptnTYPFugwdfAfDRLqR73pixKXfjZPGrmmsTl5Jy1Njb48r/H7RuIhsWPIcnp/
Kn6hlTYlvVroAFJtM4JJbENNkXiBJtkcIGQhJVW1VGt9Jll9OfxpHC4A2eHql7Av2fGaOZhMhUI8
RoxY5TieG7Wka3AuXEEnjJ3gJuVNkiL/XwvjKLicCjc4SFV6iR5Vbz11BiSoKDGJ34bl/DFTknBS
eSRdkpoPVZ2KFvfDyRUiuaDElL/MR+oPbpx3kUmD5erzq6klFyIOxKDsetLKWka7xmNcaEny8Crq
uKEjaTMt2H4fqsacus6UhZBXUL5/hQWoCy0qG9t5t5XUXws3/KbnqH5ZCLNU7vMt1yMJl7ulP44M
LDXdRsV0Ozi3X67d8IOQEWdornXoxFvmbT3EXIuzBbj/3PRFYTibSaWrjAmZcGfIZmuSUsv/H60c
geXzm3DzIY70ftNhbj1h8ElTHiI9gY+6qZMWAxyRy1jNqU3Jh1VC6DIbGy+qZMXRuG7PSGvV6weT
Z/Q6y82YhFuNPG7vFx8pGSHLhtwRL7VOUdylUpqcF++27bJRO49krP05sD+Iq0l9MBYVeSvIwnAq
XjA9tdocASGQAGiRcNvfa/vp8uXUHmfReVg4b/vAMce4f6xBIo5hc1P2K7S6g7zemW4vsAIum7Pp
NBiakHW3wh5MudG8ixkcaJhVMSLZRFsQRp1PIAFOoTTBefud7Poo4IfZZ/+TH43Iinh6wVrbQYOk
hngCGSDUasxQVPvdH27puv61WlF1wP+8OwLmeAQUb9XAh7CkSRhLZgXBCJCo50GSyZOaFHwy93hN
66MlaqOzPDVbjvaXZDACSn9r0Ywo1PyT0I9rvcy5vSVFsln47nzZDoweXGr+hX6lyrwulUZaxrMj
dPkPnjjrpOLc6hVUwy0akqP8hhYEN3kPaL9uneAoKyrlGp4GLjWKCODVF57IzNYyqVa7IpjTCQVO
w7KjzqoYNcVYFRpVnFWBRzIznJsN+3NfMFBzIcurnLfxsrEQTO/J7OoJyrJR6WQZXoeij6/dE8b7
+yr7Yhu33pPJ4XlhjurdtTmMFzdB4dIzat1eicaRdCWcPLmDkFSQdVP7d8+kNHHm63tfl6fv29tS
0Jf3NeUIRHqIZaM/S49oy1gAgGCYRrVp0/nKB0GsrFC3RalO+foA75NwoD4mSfMv7HjwI0iK+tBz
2QJRim3DmN+AniVEuT+Oz0QjYiE1hiliP/UYy2U2yiLX+WqkxpUegpfGvBRjBsJPw06cMPlWpYN0
SY9yD9TiRXYnR1+wykaQp+MSJbvPZvqOvKbOcjz10WHYQnmtQ9KXXaud975sP5jyL7D9ilR6ym0A
OcpqObCC7+Rp9nF6BZbjpApqQC1Rr2swTuBxUkcFmuy9u3iJMWaHnhyxtNu+gS4O5wVQo+Vlr6o9
MfpoJKXLWz6BBy7eLgq+1htwfcTbzQUpNPUeGtZnnipB8DwIIyZeRcY4wPgVyEcf2F7UdE6RIh8j
cbT7FAHjf5UGiiWddNu51wxe1w366Y6RLQ3dzwAPAjc2zeBc7R8TWCTQwUzJ4s2Ytfyn8aJzxRX0
xLOJykR6/7e6gg9OU+bkUNi912ISBUNvgDGWUaKQ8999fbElOzQlEFFbHdZksmSeYtppUS+N93ar
V5f8JVafI+y7UVQAgWtKswQC5VQFbqna49dOf4S2timxGXZsU+/8PBPwWkmX+1YeTc8IY8N1VEJ2
ZLlSwjrMy1o8rXzSYIy6lCDejsJfn7OxaHPnDea56r3cWh3vI0g/c9HQ0VsXxt6JSrZQLlw5OT4s
o7zQ1xuNPOoXz1KFpWu79wl3+U6z7HM9/NdBvn3ciRDFr1FcbzY5t060ccN9rkUDhC62aa+YcDp5
yxT1hf/z4vZW7Mux6Yv9Ayw0/dlhFZnQPyOFvhzj2WWResrcAnrU1jvglsOZrT3C05+9r18HexbS
R0ZXb6PXzuu6AFE40pDGfiZuKQflLEZyggXyCSP6lNZt1dzTCACV53g62iwlw7QSXcpVyAVK22DO
YDQ4Crp1EhmL8AQwUptFE9UWSU9B0nsYBLsq5cAKl8SvQnMnOt8/12URgl/9A7hnuQ/sdzqDPart
lwsDbQHo2aIWsRwy+pi2lF1ritAU2bB8qU/W23GntpTxiGJL8k5qp+uVkp82khrOfIS4X2mMY51D
wB5C44a5uppTtDj+HEoFnbfXxwJ1MPInzglcw988j4UWF5t24zA/10En0hsgalWD/JoJlPoA0w2s
kmeAkXQfFLAdT1gIGu44ylnkp1Jji+34kA6/7BBVls/P9IMjPKMRkRVW1dpsprI9wq7QqH2kQ/bb
xFL6Ky487/KNOv/H4ayy2B1V5nZ5+8aorX14K6Vt0EaSu6NlMxbnSe0qIMLvWbDOCozb1jcOy2FP
V1MGEEK5YdfN0Xem4JNZFxXJfDXvHa8N61foovOJjbHnv1BesZkFQaR61GhIGcjUc+WOm8pUp8ld
j9mm3N8GC5OsbGlhwMLHVjaUOV8gwBI76qhBdDm3yuUx4EQM76Ao1/pxwQz/tDnl4YNqxrZpgObi
sTu7qp0xWywn84QGLqYHrebNc7Fs+9EAsUEec5Hg5JHQFTKl+PZ3BeOGajNhXEA9Rx5VWXzAZjL2
hKV/Ap7+QB2AWToa+BsvsGGlLqJE5bBIiEjDbLvR2qffEcwmXfq9eN1VuUQbdWQYbES5EG+pl/zg
VFeHwGfdUaoMedJXYHSn+EIpyiEYbsj+uuVSjo//6sLhPKlBD0GfLMHwYe206DRwhgSNTroj9i/U
BWh37KSExC8AAYsalOUXxDIgpweqwNLv4FI1O/Mv6qmK2r7IovftzVEz73s6mmaI1SZ++RRS0609
CAz6mmBUWla8E9zxLmVVECMtLhsd5y65D0m6qx65NEf2qItKTneC6OxxamPzq0TiqQoFzpGaZUHP
OZiqj/38JeuMe2j5IFDBfBvRkaTGIxgGk4kXvqH6zicBYq6DYnhFdppfxzG2EHlS6oz3NSl9jvMP
NYITOqa8XMxnO6jv5Qu5tcROx4CFewkLQ2r+UVCXuiWcfIZX1nLKNOGEuYJ0i/JuE3qwrw01Sd7n
Vjhzl5JLlKB1TavIICuDjJ2+8wZW3URntqb2kHnrg2uyHrNWOgt83VGb/LF0mGqiLAz0MYIMahfo
0sT+1UqeZq/ijsaLcM8zjMz4QJeRcbhs559JgtwdKe3U3MiW2+Y4N3/rNBeazS0popw4wK9vQdUY
iuoTL1WlwlXUaXSXXAV/pv2n15RBcDjgddlCZ022K9P+hc+ZvmPPGmdofyvyg1w9o9nhLltu0+2Y
iIDLQiIs3fS7MCc9fbyZRK3H2fjYjrdDzM6eCR705PjJtYalWhogOfcOUz6I6B+9Uew981G87gwO
Nh5ob4l5HV6Ie+rQJEQlRbGqD/oteDP0xrX5LIUrIC/ywJKNm+9S8LG3jimvU5b7Os7mJG5ROGJe
pZCQc6Xb1RXqfxxabOc4wjJzY5Dwa/arnZ+x1A8y76YLXKryaosxz00K6ZzELNhevEr1dBaUJfSc
l1c0V6xfpy7ZWoZDRr1k8ki7XWLeo+BLU8aKVc3WVZw/vxLPN+GkmuRNktJ+1k4jkKPPpbTAkRz5
1xBN7fLkZl6dgo3end5XdQzSvkRND/izkeihyDM+Rb1Ccvs+gfr5nK2uKvsaBfODdLs5WXLnuuMc
2Ur25Q/9ZAritLgJsVNS0A7ibsJ/gRfoM4tuUXpAlGDq6IcpIz88BK/iZXPBKfVPX/8tgOPewdtq
GuqapQMN/J6HPnbSuvuwirJadsRfrgGajCyltXjMml1ETDMqPKtwQW3ZznrFYM3Zvsxwo29+9iLB
ox7v3rmY6wJtMZmnJnj7p8cECtTAW5L/uA3g2ilkCvK5wUAQ8aXOCNAAofmVZnLWV63n4A6DUJf6
2TXKxykq+ocI25F1Dm819rXf8CwEEpV9UG5SQ8naiKtGdDchz2XRGuPTtvXCl9DZbqNeLhpQonSN
Gyex7sqCxijgEl0h5b7EQoe/wBKA4U6EsDt1XVzPyQz8mG+77pHPtC2l0we+3eWNNF16GLJRMiP/
GEXo4mODipDAYjOp1wqhKt+Pso0+Xr5cjqfSY480ZZTALjbMY8NIrDjK7v+bkkuphyeoCtIhd0P2
2eRbr10D6KylKbWwIwNZ+uDv2SBLkmd8/uYMUMN526GoBqkH4JYFVZfvsvWNVAbEhTv4Cpp3BDqa
DKBPy6yCdsYHVT09blZ1G939LrDGz4eA9iFBLjHdYDJz4UzOXFOWwqJIFgRF27GRDGbuq2qAuCLM
bNpjShJS00cLI3P8gvXJYZEixbkXPDKKxXyzXFCs2z0E4jWkea4o+mnMFymg5eJ3in6pNtxAZsHx
k6KOjKPi4fxPetMrsUalmYlfjm4M3If9zwIywiqthjfUSu0mTA3bMlWv5K6t8Q3X+wLxCZYmLVWA
+NGCWMVT8FwUP34mt3pmUpBDkEC4GZBZeUD8pFCFhYO/SQBuXdrp8h3ZG+lHNaXr1OQmQhVbZXkK
EUw3Ea7lGBLDwBopUnUCD71id1FhZ086xMkIu64LGTpgdZz2eEBr4M2K9YoXe/ydvi6Fn1BOHf0S
JQ/+G2XLDQjnI6Bn9SlzQ8DK7zf0GY7U2rogtwwQj0zIPQHbjPozE7Mqu9BycMpjV7KnoJXYvdnG
gCOSMU+gEqynWs+x0qbHebol12FTM3uWBtHcZW55Y1vKkYy1xn5j6Y1OWOIz66jXxX2jGkHriQ/j
xRVsEX60mNQwEh8wdX4fiM9F8/2Ye4pvPiov2hW6k6hnVjXBnyB0VYptzo9ahZujP12c+HiF87eM
MdDUxjmhmlYRaL04SawPXyYud1s0gkTIEHi5z/j1p/HAtVEgjNZRexM81DG0fHwQL5By6cjZ4sBf
ODztWrt8Bpi7gMrnul4zF4pPnSCaXU2ILaZkQ6Ma4Hyl+zjlSBRgL15wIskKL4FwI/PpDutdDWJd
TAjKRMzzvxYf3BZ1bFcRc4KwbpnPqF38TzDPLEARAEwtS52p5dnAhUReatZnH35YScQP/eT9S9iB
sw7iaPIq6oFc3lfuUkYSCZktb4giNfWm1BsNvtFkqfrZtzIQXk1NG74C4xr7lrmLw8VYe5/Vd7JF
kf8uwWsLBL8L3P3LWZ+CB5WDbT9I4yVS0uB7AQrBN+oIJawj/5n57PGn5lyZLsdmyak45Lzz0PCZ
qHhK2tiGpPxStOGhyV3Y5qfvO6onIU5W1/fVkz0UxtoD2nu0vDZtLtfRt0GiK4YxbF+PLfuKU/dl
xeLEhaJcf0o19erh6bHImjFlM5n4FSDiHP6KL/vssYTtPA8yoDmY26nodNmd3xN7o3giM/5fmN0S
PtaAhKf4vp90vXkmKO7QJO4kwwUytwEHv5m5YRrBhpsIxX0Co1hp64qy2HHbU5ffkePBlaCotb2R
KCqWwAeiccVp/KfJvJl+gE4J908//F8nY+1SuHRzk9RgHOvouY2eukH3LlO7Cyw1aZY4UUUhykCp
qV8R/kg1Tu3ygkadIiriHJ6wZT3DjEWkv53lzQhCNkVjkSoc4P7fCzJWxezH/1qhMPdx15qoGpKE
XfTLEIyoB5eH3xDZ7sq7NPTHJUCt4pHqPpMgGddPwqOoFv4PTqTAepUNrqKbxPgb9hQbCUmln+u+
+CZqBqGQa0GHz7ayAqfPTM1GQKR7btHuubAAoyWSbS7XqzvoIfR2JzS13m2QIhZk4vrZ+isyF12M
4RMkRka+i7o7I3U+7Gr1BA3OeF7w6rBVWqT0KsIs+olMyqzYT6VQs9dJy2e6DtV1O2SsOm6g5a63
V4AVzqueMDbJI/zRVSvkRiOM62BdMGq0/hhayaYjdr9nNcq8kBHhgSFpBu6ZKPJ0UyDTPiYv9+lr
GK13w8dFr/o9s8/i86Jadv0gv3uqtcu6IDHANlyhxKerfJi+3AM2znDPQgWauDW8W4tYkaHHdtS9
+KJpjyWHRa6GTVk1NyrA8Mbyp5ZZ26fzPe6yhbwVsQ/nlBR1kYGhJ20s+TSfwQk8YqPOvVqvliwE
TkX5/atIncIDZKtD26uGKkSM6UN51DCIsy4RJqQ+TiFo9kQg79KEjvmwp0OZ6bOmMOKrTydYwyp+
AHwxTYVy74BvZRk2oTY5f0i36qcdY/Au59UrXbAZrD8j9VqkQyEoxcn+G1WqFdS3qaRu7pJD/ipu
8rnfBG/kNhZ6PoQyrZrliZ/uTjy8G3W15D4NvVK7my51Ml+/m2LSxfXGR6ZbInkrOkPL4sbGN9LG
WJ8jX+Keqo8uNbUcJcjAvG2V0Sh6haSZn26NcyUDywe8MKNeLZHqPRRtW3hVRrOdxtLbRWMziAcP
PcPSznNO/8j9xY5AAuX5mVPtpNO8OC6Cq8FKjI8KdJvvITHpq5PVQrTISOt2NEJk8WbSc2nr45Yn
Av/XtGJeKWPlWzL7PAMLbKENmk6Yq4lqjzrN3vb/3LxMeg07XS4kQ3u3CRbaQZknoTqk8JTUOOYF
xlC+FgqVnKYn75DjWppBfdIASEJzzieTEbIJ14u2ZXV/glPpNKfUB5inRZTELlPNUUnfNimlVdOB
wzFEw0+HysCh9dm5bb22bY6ZMpFHtkekLOrqO4Vd9Ju7rEJ0GM6zG7meo82g6G4x4lg0KVZoQVw4
pHdX8Bz8yzkHVj9S07MPMEdVydk2XF4Vm3AjXheTENxM+L0jUf7BVaaUrTdPPr7fZSbtYk4C8v+v
c+FX9o/Qard49C5T+lAtTTlo8TOqBVa0kuOoTvYiEHfOY4AS8FR0rTA/zwoZyRXeNm1N9HGkkohJ
P0CHTztWC0jhqohJTX9jlc78DG9Ig3FxZpp2cNcmJ09niYufog0YY0JRRFigeaEAIdJlu/mgl+7X
TdLopb5y8bkMTexPCRutq009MmwonsbNYPuvZ8MWS6iyQaPBivqaw9Ys88wbTSOx8twTIB4JQ6oy
nk3rD5hq82psediGfb5AWUbq5j58CySnX4YUCGREMtFbKkgR/EC9/9mR1VkF/srmGqm9Q+FcQD6g
IXNLKtsru/jYI/j2ZxShHoNywlLTStJubQDhPk57IW4lDszit6nnf3fNX2cZffXww98kjGqyktHX
t+CwWPIFZoUKI0VJaXE6LQ9EjaCLBJt9I/785RDbolqMAjN6Uuk0GfL2LqnywdvA0RGoWc3NQI8P
4LjBTfZTFbsXr0CyqlJETg/RuYsxGRoZyn+r0J4Wym7XIicv/wNPV3oWk9N+j1fT7nnvzpDPQRZ4
s5irmLJzZ2gR0a1oKE70oN68oJdG4pZxubiB/gEIe47kRadZjR1EHptrS3HYmRY9210b6wz5c661
XKyAXdIKB3wdlnU7mJOuYIvH+LIPzI2sSUjc4eOmC3pAEkMxWHpUB/re10Uoya25a3vzxyNPh/fO
bd8dqShR2VCmuPuoSiEj3J+RJtbPcIKYZX6agHLcP+yZ2ZPukMb7pAUuPeGsj2DopnFzSy1k0Avw
g6VraTF2chr6//ZKFuJ7pZQwpUU0ckHmrrGc8xCVYbFmO66yywUme28wSS79ofxMLa760MsZWH2A
FzSo70/WwD2cidMlpp6P0vmqa3qGwkXb/POYTdLWQfJDbnYRTqvMMtaGwTafnK1iKHkRdRuax5rI
sa7JA7kX7tSWVG47eo0RlkH7ZkhNXxHJlGgvvmMCdTtPtNFBGhgXOZ7ZgctfsoHluCL+m4gSGFMp
RKOW1sEF+yLgoUoUBYLxvSP7DnmaPlsSbjTr5GcUYQlsVmTkOo/dUZ5I2SWh4iWcxQ8Jk2JaF5fW
FY98aksSm6NC2jgKk7y25gfRIC9WkJNt7DpaTQtHD2LDvjKU0CTtl2dZ0DiqdJyJb04D07kLpc69
pq7ESunbOp811J92JXBPw/kYKXkwOdlYl8zIebs2CXz/CajKAvpL6X1xS/riJuw+/aJeMgh9+Nlt
/1aDtZznVJswDX+mrl57Ey/okow+gZ0Z/Q2SDXdj2A4RmK5eL1EuakFNOVOC0QMEZfnP9ru6QC5c
bNgJodC2454Zpf2bEc2n2of+RGN22T7J2cvLd8Z7lV9xBJG0jrBes9y35zhrLnC+SJZxrVIj2Js7
ppEMRGP/BeLPGWYr+q2Ko7CFSNcR+SJkrdayj0mp0AolQGs1K+L5HCwbFQmSEqSl3oW9zGrCJUl+
BZe4UQ6LOlSzpxtLwOvox8EDClaHdsyD+JfAULXoIIT4Wg1jGHDxpAs3PnSRrmprKL6d8MFNkqbF
N3vFLNysht7mAnPUKZ0NIxFs6MLvqC0AzfaYZOoumnn5PpB6bMntGjGJqF6FiFZJ4WU9Q/Dmhkvd
7ECwQady3Ds3i9O/iZIMmHsoqmviGgUvRUIn4ERPzmmlV11CZU54hnvZCmCJacoSGMo5qddynL35
ZwYbF89Spji+Jr/E6qsQqPB4WgM181RFhqu+RI1cq47AFc0lGusC1+ZiXfEIGwJiVVmSyvgev6kb
bXfLmLTZpZ/jWc5qIxZRVRnOTwRFT9V4BISWrq/UGN+bWJK+rhT6w7ZXtDpMk6PhcCtIp0/ugKjr
1z2oc8Y0rH2tY5XVvlMI+Jvex+VQKkYOQiij2ydi32nnkBL+RFz21Vry6sze0cO8nDjmT3/u/VXI
KY2AX3XS9HZ5MRdR52LEoOY9wRIfhlRW1Ami/NhxVz3RQ3yElrRaPltrIJKgWXO7H2E33YRb1pb5
YQInQHF0nxOO6QQLG7b6Q4lF/95Tb/uWjrartrFpk4sxSmsnUeWMk+JrMK7QSnv7MQCk3Z9Z5Cwk
3HyzI3VAbXHEBTA9jSPAgr7vUZVtA+lwX1bLeDgRdkD2SFMeMkooxY22UMzIWt+R+p08KuR5B69Y
+FxN98yOumxpn39UHbwn2voyOG1V75ESDGUVRgObdt4oyLpNV7RW7IxY80bhB4+24kR+LIWNuflw
sD4OKZV6FM4ZL7fgXzzVueltidkn2Y+bh+KTW+iF9iRJkoKrHSUVuQMBR+TIe5WsxN8Y1eF9D58J
CYin0PJgFckK5dbltFKUZO2p65z67ki28/BfeanbSu7JAFUHKEmzzPClvV02mBpIvoOw/WD5h6ds
totaxU7/UAe0W8vy0Ew5vnlRC0VuMlnihNjhOKH4ejwHZ+6BQz7xRFh9XRZbwCLFWROrYbGl+jns
isehf03ULyuIllL8sBdahkfEwX9xfxiUhFyBl8Rkxjnjsbt/+QO94ik85RvpU3SaK/YD8nhNaREK
T+0cd4ZBumInjHjjk7/Ek4BaLcU0VuPXT3vuyN0ZY8edyEVPYLdG1U4SKjGXGGK/HB1vBM9pi/1Q
6oWc8ACXXgZr0vIuJ9R3HTi0tWIUbw+Z52q/h6AHeuqlTFLTzslJCKMwSxdst+P3MpEvKPKB/42h
Lkjt06DDv4RlCr4FekIFrGfwH3l6/O994SlyvKNUh65QVI0rMS3+YW9+8+geybrgUse5Gi1Kwc9B
4E9wA0VdKdVh1dia871gek/tfCiaqi5IQPF/lmLFKSB49bu8UU+q4gIw8bx7JDT81TD0GZEOXRdP
IEzaiNLsWcnseO05VTObXHb/xzLKdwNGm3PQHSS4unWPt4WvNAjXsSNbep24sjXE/FANHKJSbBUa
5ZnVagsYFb3lrBzFGzaSvv3lj7iwD9Ocmx4OOtEffbNlBLn23RR58m/NKEZvB3kx4TLjbJJ78EBH
vfyUEa5JrIG51MA6tyhLi9K2SnY8WAR6twfK8F2VFoj6FyxsW6AJXVvPvnXhhvvK7vjsqy24DHr5
g+PFdIJcIs+Dkh1vBqoS+KimKC1sVW+Bf+Qb2oBUY1iodEptapzWfaXtSItTtFXxdTUEDXEsDIug
X0QSNml/zyhiCYrJTkiB4Ml2ThRQD1wB7FvRC3QQp6Dduz9vUyJVHihGH/6kJhWH8r3ppsRbsxAM
EHcMVhh8aYxjYBbG4W7qMjKsFzC1UQF3lNj9jc1uo0kh3Zm1XUQgebwGrXQo3A4PiZMCPkfLrLjA
Wic7nXy/RuoiX6B7BQqCzbPC63QGIHszG7KOG7w1ABrZe6unguLbpxu5CCOUzl+CVGhkRo8XEldg
Wgqw4pYgSgvbbWQvlJd5wpZp4iRMVk1dvharwl66abNV3RYNerhEuoEToJZ1c55qGaIbP016zjSm
sEylMqqx1KvJMa61HaJTM3a81eTNk50PXu49E4UD/Che0HhDlH79kgkDNmUzoRQ6lqCWZZ14BcA4
S6nfgpOtG4HFwhED+e3Zfhy7VxHnuhZl+aRpXXUetbt+xvdni9XWWxR18TJXkYr6X5JKyJoxQGRy
MOPwe6+b51wvABgnBtSlaXrQajegtRzqJGho1I0ZgsCh2aH4L3254tWu057CElrxId7FZZDrfDgS
Jl6vHG5GoJCj4s92u1cv5JOXAdBNNKQO2Z6fuXlLfTs6byP2YTjcn/uCJ9ZcGBtMsIDW6PFrm3oC
hf9YJxshwGlGSoNWlR29RmJisDfXkRIk6O9suZHObbo+OP6KxLDPrSQkkg6rhRoD9pYxrfxNzhgm
jtdlzW9uiwaNcSlw0gvLayQOyCjUDNuG1bpXmbAU/afT/EscktMfji5X88mAPc93yXQFsOj1slEZ
IVtyf2PjdfJU6RAfa5sgvbov79JH1D1I6XwZz6Isk2UQnQ8m39ptuUBjF49o542cQDhdxIFKTlYs
Uv9/r6udrzFvhAt61uDi7B7tEr+b1Irc3KCeEvTb/XeQBqCbBSKmORjE3PDkdcVyNY2hxGWgPae7
RlB0xUa4ZS3zh1aky2pSn8a15OQqQvBivPr9pDYSUwEx38cG9mxJDKmOwYvqWFGxNKSKZf6kBJEH
Nf71+SbDVW3sBu7yx55BPoSP8RXiTKI4PJhVEKk36GpRvqeFYffnrqgQdwtuKHwdbnDgnx8y62VG
9Y+QFzMkonvffacz4mPoNQBbvZtYI5l6ToF4jAFDZcFJZxG5G46P368Fh8XTlxYHxs0y+cHbAwfY
trkHfHWxPUGEEouG1ywN8uWlb7ax+0fF3EoOA3NBFJxNc08popus0kRkStRIMeudRSSpIJgggcIe
gOzwIMbCXmCdy6bMZtqxxHsIMvIScPWbG64OkTMpz9ORws2wgq5Om6o20IHb18wmyHbfOTv0882p
HO+OAX4r7rKHBj9o9utdbI9ODJH8wYoF/DAzQYOpvEFy6fzri74CNdYStWeyYm+eF6Pbe0M5iwuJ
L1pafoPxXgd7yPOQjMoERJdO38kLVjiCYKHzKXKwf24JhOH0vzrapthFdH2mNFqRUDNGwAvn7SmQ
ph+3OEaSoniKuBFGLrTcz2ctov9XY/w6BixMzVqyIUBIghQ2qrJQ9+x8oS0Af6RVDk65dkQPtRnx
3gKxesFnNUvk2/5cCBBVTwVs5dV7cHIFr4e4JkL6J5IXcRUPpexlVKgu7luKyvu2NlPoVFHnfKqM
EwyrSb11oh/TU1KNpYfZxqj37ic/P9FbGykkWR6XvQwL+mnp78Niuw4jo4mGfVdUV9FTToXTiBuN
cLVZIvZ5y87aFqEjTg8Ic385NxqhWkanCV8CTnN7DpXWxI5wGqwuE9Qv+jow95lk9ajUopFo+0Dp
h0tmP/i/8kZeeRQH5QxSpGEXHfuyEPH+ydsOnhCdk3UQWUnM1qhDC6mib4Hbo1fbFkyJLY6vHX1o
XYqoK6nsDN3cVOtcQYjk8Nc57YF7+6N6XyzETMoYoLqLKpEu1MarFKv42Pp1BF6hY9GZlwSFqRc9
kcHNUmyOBGbeoqauLhN7wNet8twNQIWhbQwXv5FjkIsoKDc47e8KYTwIt8Hbqr+3hVcmXWnw6TEt
LbnrnmppexqPkA/MV4mlb7a2FQ4g4gjNI0/76i74YXE+J9YXLl3prWfYu2AvAAJHqyp0EB0sW9WQ
Xr8hRcIwHPEaKxj1+6rR98tB5sBPv8QoUnQ3nNs3K6CIuWy48Itx86iPERvVgDWD1Iz0Hv4ksqYO
pSuWjCmjT3rVjy/NVTcLgKJMQIV1zo+3zez0DpwLuM+FHQZnPl8JSX9q3BvRbamW24KCuJiieIuE
c/ELDzdaV9+aA38K4/cNBhNPn60rMGQmyrU2wqAkK1+Jh5BSREr/n3ZA81xevuMoNqZLA/hjPATE
5y9K4b0UkGodMQ1VJhmBZeVIIDpNa1bt9ancmZoWpgKF5x62NBQv1Apzf9inaCh09B9WBT6EI/cT
lMHaZnP7sAvS/oUMGHpDG2sYBntqhbGYAu9cEXzWwJLkg/v6scugDkFHSJUXw98gePQ6nIKCpkHT
jgi0XW6yVvUpA8T4DOT7QjHrubRrnd+xkCa8I9X6CfLwvEUHpuEeKwt1ZxjpnswdxWIQVVGysuQ/
Cv2k1cgQTOgFEP0nrbpFH8lJm1pac35N6WzVYnIpl2jEZGbEaZalPFZP8OJxVLSpLU/IFl5EnzOE
W1veoykctWH3nC4LhPdEMErgSBoNZ1aOwspWtQ/lsHxfsBx8vIeDkNqCkBNtftgswDuzc2wRBPG+
nooyhwsMfh31o+itCI4a0+7UosnKjsuh20IqGr9j/95i8C6tNO+QONZBQQDGF2eEQ4drX29miJGA
teexe6cbKtmSsFDdjQAlYa8MEyaO4M/ZqowswemwpxCASeX99REVu6kOVI4ZmXs9s6J43WaV6weF
YhEKuZsgs6b6AgXheeKKTQeCANLV+0vwKPHhyDp81Prke7BQQj9LBPMYvvzJlhdNK3rdrfA8+RSk
hdsqjPNsSU5EdjxZdH8J3PcQcUqJGpFsumbQPKEfSm+5GrURnN0F/caa3yMtsNpB/TatO2YQD5pe
YI4POgkuTEhicROtUpnb205Pe33OXrVgXQfxYAvnwesXrf54bkrHdWZdoMxVhYmiUmZIYVVi14+m
nPLGdum3Ghci9vhYKrVXwFwWVwesIeqhPnWBBdu8crL9BS3unJivc3/YTGLxrQur+ZkVWX5c/9Si
kefmjHsB84SJJI+dA68cWCWayk/KWMDGdckr1A63vn/Tk/YgW4WhS6rCFEzJMOls4GmScKi2+yCi
rnFdvxNQFnchwxPIiamzk1XJi5lZauR/61ScAgdzKJJJmKR81RHB8PYihcOMo8Rlf2003yHtUdO/
5vRy1gxB/91qr/tcTbAIrmyCVEk8dAgkVsggVTDqQwybV58P+7Va2WC9JY5YhZUIW/Huw5XveLG7
lTk/u8JiV1cMO/zQnl9u/1g1g5WyrcxAH9uxJgC1jH1NAsRK2lv6bwAI3D89SZ7RQWfHPG2k+4M/
UiwQM/uOwJ1Hef52I0qRED05wQri4xW2CkAR4Bz4sA1PiOXFLrkH9PjfAKj/qZ+ttdccJMIswYci
KeiZYhx96PZjGUcMbIfZdaJi0BbPY/iG4ZIDHnqOxTXJxy4Rr44/tdYTKd9idddgXrd3Ngneaxbz
PX5r71Di5S7OBHzU8/eRuRNf8p3fOU6kDVHts8Vk5lxfLbO+A3xRJFK4S72VHlvDtzCjF5FvEOsi
PghOYMoQb4LbVB/yaSmXEL14sb5xCMcTSivE2Vr87NT+K19J4HfnOELKe4gqDHDYtWE4iH00heqG
eQN9riMbgHblix1jSY6l29V3yMayyvt+NMmy98u5tP2D21yy+bb1WDfxYwFQ0xrpOldCBDrWAOWT
Tx/LgWFxkyLcVHje+8MjzKsZp+dQQPcqxcmg0/CyPZ+ryhLq1By3q57OUB16o/fmaB2cNOB0ZTN+
CdmTTvrevwGKuBujJG9lClNu/uYTjlqMjJ9dOUA96+owKGDCPsVq+INdB8IwAjNQBpOHwuAtTJfO
yVk4cKo3ZULuL9xnOn7cCakT9MUxMojM0iKrZQIfpGKAqR0wXDVbwE0o9L/HLLVOxxw8/pHfksV0
I20lctsvL0q9ZGzsG69WFvT11M1fxzkZeyoxn7uATx0fQd1rHXHgzZi52rQJAnHSo+xyNfH22TIJ
XKEkDOig+KA1i/Ksl0OyYSDFPrcGovbSYPkK+IE0xW2Ga5JOvX4MuiOGrQy+WCbg1GKam7vZ6N3Y
Na5RKCwwoZTg1KFbI73k18kWW+fuGDbJ2OaztELy91P3ykHSDhjhHEv0NUXgi1RbXHA/fyTYyUsW
AF0nj/vF3l5+xf255hBRZ5JBalOu5o3jKZfry9DRRic3BF4hLet3AueaqK7HkMf2kff8lfzzOViB
xVSWsdL7YqZw2JSOrWwlGawhapz/k3NgtQKFo2bRuoSNPJOZQ1Lv+CpfDyvbV+yjeElmVhleQYJE
Cewxz9EEDjo/QB41XWdCVnS+OA+GxfVSXLBTEVbpSSvRoo7G8gdisLyspqg0WOTDV+li+yRRDS9C
Ljr1K4fww+NdD4DxnKXCC+GZzIYTBbqF0Y//Nx4AmvhhvQKI1AQtPwHAP7JMBQOYyEC+GqNiVbwE
wZsFfjDdq1fZVTzuHMjmaHHMaatkH5KXqFeiHm4C6Hq0HO8VPwjeMJ6/Gkb/VBgn/qMfMH4BwNaX
BFeO49GydS1rsQ27ENsKHln/W6G5rUkfpsuDXVSorev/2cSRug0zsmRi8HudvKmGQZDZmmlaiIRw
A5kzki99S7LbBlJk38OMWo2ClAV82Iiwuea6EqPqeWhCMPnjZ83Nqij638lm2Z6E7erq0+wPTmpz
zIarhOr48JiOEGLld91/58ECDImm7Wg6iFBaVUNE/6BaFKB5jEcP72VjPhXIJGNZTGfirq7IhhPH
GP1nvmrg8PiHr18ui0Lz4BJBkEq2mXzrA6r7prdYkoendNEGAHCngFcF0eTrOpHhny8xyaZlrJqg
Gy52ZqTqeDFginebCS5j6q+nQnCCgX5SPFoJCERXoCxVU2B+YhirGZixFG9BvPh1hlcfukb924A9
k2YUD9B1RzJczCMT/P0j7bp8js5TxMwq3BxDd/69pSyY+ZxxKqXw1PSkGJOdcGzGF6kL8xZTZ3gh
/NnVAFtA96eaqTM5s9nAWelFY2WJtpevLGnQrlpIRDwbOJ5QYcYoRrUYB6jnfTbVor3LUe0tYWQy
P92PVRV1L+Ws+eyW4O2x5Ryj1hoVYF9lSzxyX8M+ZmFD1VXd9tauiBPgft51mHI8JtYtaHaAP1pl
+s/VTwhMHYt5uQVbhR6JZY0W3YgC7Pn12BJ/KIQuoOF4s9u60HhObMelU19cNZYvh9zkeG9ljAhf
WJga3Xi6vbYtzDIt0kt7tpGWDEWOzrLP6QNcH8dMLF5nEMPAY/sh/SaEnmn6k8xUa13ssh5fyr4+
XZX70Y7pF1z9+p7olVtRkJSCE/j7hZ97tyGcnkXugo2zqcnQ7ldwCbcmFCgJ+ojOOPsdr/XW1vp7
cmfEC2u6vfxxODxNANyb+y3Fao77TLGo3CwxXqMIDkuKesftYn005nKv1Ah+3g/rFAUML/MLWpUu
lweYAh2+bMxQKWljyGYwR1KYnzKaOUb9Av+RyE3mOu7ozWlWeVWmyt49d3tI+nIXi8Ovd565znBB
L1O5Ef36LyUFXxku/tPdVCpeGQXsDOEzeEN9DRhRG6SKB/pFGlrfKA0bUKUnOg34TqOJ0dX/YDGo
oXF6mk730FY5QT7fuGOAJES5yyZbebc1wh8SIZm37TX9xXu/TvCjobL5wyHZ3hwDrJ1QgaJ6MMWu
q1gQ8gqQmy8YiFrdGfIu3nqVJNiYWKWKfD5xV6EIosMC3Pz5+IcGRCUCTUj8zH3YkBFiMbbpaMBE
AZUjiR43v3jnaQVvqyTKgjbdfsfVwPy/Sj+CR+JiWYTQCGk0o6H8zBsPS+1R5on9/9IJswIIB/Up
+KbTrgAbuJ0SnnEab3CnCWda257+dg8F01LlsQ87bf03iHn7BzOVVR5TRc5vEoO7q1bknow0yxu7
Ut6I65BJFTZ7DmbNT/IAA1TataDe179XJ8t9hc7Ju+jhaSJS+WtaFeteiOTep33x9jhmOzEjbVM8
QbV/r2DZOY1UJGZIhyiTBaWYZTtnxxXYoJqiDxF5Xk3t6q0N/tjvhrr+ET/e+Y3sXFdtemTTYMoH
IyhGWtkVq50moJiVPMkYuUZbOrAmQkm6iLTUWZxiHV2eTZEp8v4/46VZu0YGk4z/GyGZyIFCMQ2+
qyyuxeDwUHqQtkv/X/jQhpfBskq4cVr2WJa5rUsjE6At4Z6oMj7+T6x/tu5/H/o1e9AuutEPe1hq
b3Wsl+Kx5+7KkJVqFgL/JpWfVrNa2g/LHWko13AKxsigIiHHDH+6gtNSx5WTKu1y/69Qcl9beDNN
6WvNlKjAe4Rde3EDr2CpkZHV/Crsox5dsSrvd6czK3V9akZNbgXsYgCtQkIj0/4ZfRGtdLAvm52q
jAEmwVo4lDL/YmEr4mQyYDr8dbF2RqPnYCXVkFF6IVO8MuMIsECdUkqSOp8wjaV+aQL3CWD0AXWn
uyS2mOn/3C2ORLixZ9eNhOe3manu7xoA6u3ZwtGyzOax0H1hyQUTZTMvrNNPA8i6MHjAwt5bD27I
oVYB7I4NqtXdJ2h5F8eMx8hBlzTInm/clkqatSumn4pYhOc7jGdG5YcUsN7XQXOLYgGPlOGel4dK
0EKBWojEre8pyLG3wwD373X0WRzVJb2ez6TIl21NTkkuybwcdHVhqo/GswRUWpEZt5QY7Jz0y6C0
9m/SmfiyGK4JQmQ3BDHUsEZQuj3BbOZn1tY1nXlT82YZhPDloUL8RJoJdEl9KTwTcQVRyKqBOOMo
xXUz6IUM8rxIdQyE3T87yNiiS1m8E5FGSrltRSZLxOxk0Vw8NFgm16qQg4toOAPIXbIhxCGE+hHm
AKctWBfgDnWxqqx/1degbyQ0WxVx+0EgFVNM8FWKkJuiuA3/4w0UKfP8xKraDANXaSqFOmnussqJ
KkI0jNwDl1yUx1IKi+dCN5+JSXboueAe45CiSbzhI5VKqJqYNRK5VUxCkg4jdstB+uAqUFXbgENL
z1KVsgSinB0STxuYKW0z3Zq/THZ372vxbvoeS6x3Lxd7AYLd5K8u8TRhVFsvLXT2/E9gRQqwriD7
9sT2tuO+irRIbv01OUmyG2ojB0FdjwHTaYwHPMWNDeh9L0N2MMa2WGujXA7S7oJIywhYgCI8m8dJ
ibahX9p/LNeqQO+IIcVNaXgdvjnz378zqZSAo00bFbazm/CLgKeRIIzuEpmD/WwjUzfAnW2MpgGL
gaLBrEHyzoO/PjoXk6nzQcMyK06j2GEfysZZqSK5wa9JdmsQIxEIItk76b9zRpaUHX4U1TG4Njii
EX4m+fO/SXMMZODCFynUM4QlCLVKDRpJriCOxjQWF5McT5PNJT3Uo6gWRFUCL9u8uw/Aq8jTFmDc
3XhXmDisup0ZsxWBnVENsD06KgkejQvGcufk8gi1fhCgy6zbpbrMMu7eH+SBDDAEHltGRP4JDVrJ
H6GuhhL+ZRpzwnkePoXitWkUSxnxZQFJZao/MHLAh0cWX42DlEE8vRrlwd3t5YgNIuwH6dN5V763
Thvqllc/kES35GgjLw/6VemmYqs9KE5mUMs4q4W0yT+FSsiGSc7pSaxjjkdtuY2YWxBeKD2hOv5I
EpriVH74zPtgj0F2kvOd2tKrusR5YYsZpXbnfTIt2nlPTFcAvEMJQl9dgYA2Je0l2zgqaeODtmKX
+ejnAB0iV5JLGYzTmagn5jdHzxdxTILAGMTxnq1kY7eAz+Vn/s6d3vTe04UfmBTeUOneJVWmxpwE
XYbVEQpTMC8f/aSG/y3lG45gxDVuFCwgO54yNPeddSRx0iuVZuUyDjZ+KhL96IyGgfObdjAQUhb7
5YCEJfg5YDsIP+Q8KcJhri94sCUFArnvwi+j8Xn8WkNJZxD/Z2CcbRmd4AwaEIoYVuWmc8LegyEM
U8Zyi1SepatGR1zQ7J5d2Jc7QjCf7sMu85TFle3zTIje4vhxQrm37J4mQgDFY6OWrFR9W0Ryh/H7
6MIGnlU4pdDFWvUAAUm1/F191xee4pRrzvvShhioObSuWnFVECXGH7AYspDFuFN0DcH6wMe5a4RF
26WRryzLuHNk/PpEaOdRcYto7YznvsaBif63ve9kMyDFJhgBPmQOJa8FDFWZ7W19Vzxgt1DL1ZTb
TymuaMpNr/0Ji9hAk40eH30/lVdqAkX8zobsZJQd/HLUi5Nvc9wfLJXfZ7KrJ8s3Rdiu1mUNjVgL
w+rVi+zd8VSS40Sw4I7jtLcxLoF3u/3gywbKnfrua/cUdFlJAm/2XJ6f1Pp1E3UXQs1OrakmkcHm
PB75f8+Lw5e/GfK6cAgs1UlRLlbli57p3tklSvqSOfoDK4woboA8Hrg3M7gES/q7M03WJgRuK/om
XiFvVHcxERwMk2heVtz5D1zOPn0aE+x1cgm2SH0Ds77Bs+AjqEfG/BxZxFnFcr3gIXmjoEaE4fnZ
0rk7P/4Y3km4xAQWbD15cfrl5T3rq4SOYT7zlXgZm2pveiOAUl/VEZVe3oW2UfYzqaTjPssfA/5u
0hvNHQ/EHnsWwYYNQ0qKscZ8foyY1uiKk2Sicm07o21sjT5VzjQa6Ehqf1jTBYrvVxtAc9H+jnqX
o0mzQws7F/n/zMWfbBHS0wM43B+GjitJl5qpYQmNsYQxvgoF7QRytf0VUsaqgr66Q0FPhnNBrUMt
a/yXUocljZwfJwhurofgnmeZHcao7tEAUstviM3xvDAIgPnBM0TyQrNnscrn/dX/0irPxQrHfNzm
barMJeemNx8jjCQ2fa/MBghfh0tfNF8yMsHhlidTGDeT1nzZbFqaWaDMDi2NFAjliIXM4AtYdoMo
nApq6gAvlafTMF6PCvERhJFFB40ZYojhiJ6CaGuTi0JoH7I1RhmIUKutaMgDScFQPXsBZsmGv4s1
QhYC4TW3Lrl2d1Uas52pvjwEc+qtdq9fvh2uXN6XACCD55hQyDIkF1JgiLnT7T5EvLpU11Ee7BIN
SpfkY+mOjCrradOA44sEaAadIqoPnX5isyunZ/BAn6aNheuwOJyeHX0Bo+TsTMnu03G3lFijBFk0
ukgIxpSX82PBPsNS7naHzmqT41FTvUyUCbTGzIol3i515qm+Zr+jqhRw1xa2MsbNbzSahbrUuCyu
t5E/hBRWrjNHNOrmwqyKZXGmzFiFpQtdr81Hgw58yhIzc4VI0iN1kl1LrP9IYRTScXmJKJsmqo2/
3AEYvsaCZjMOCXtUNi8jnNdlgigl9y9GF0ECQHW+KfywezZWDd2o7cJNsWRwToVe5iCITVq/T1kL
W0WCi9ZAMPjBnBkpsyMOJquzvN9sWcIoW47tJqjxrqxicJnlIuL0zjk6XrgSXH/tkIJRd2jDiZKO
2KaaFJlqbodCMB/j+Op5XYL7WHFWaVUWoFV2QQL08nkegZpOn2XW1a3qzfeEGsXUmvFLVvhDdLwi
+3KbHAPdOEUZRDMJKx8soO1BpzdcJGPL54aB3JJcNqoTmPhlwyS8UUM0aZEzJXR7tAe9C/JALbra
Wv8E+4dJdO8fwc09ANXqO/x7/cPNFvco6ssISyGQkLHbFwMsf0EbM7vRlQ2h9+uhIizhKbkJP/lx
f3LtK4z/XDsKNQWe24FJHBb4IO2qMUORJA916/VThR/MEWV+s+DXEM+jOnHbxAbi9neuvAOe0TQB
/YIjVl0scsQsfDe9Q9tJRNE8AvZJDyTT20pCAYLj9mEFQICjE6Jo631XtoYau/G46g80CY9e68Pg
6AA7W9U3PkJPXW1ruDE7Vpyd83bDlDmsAgJxpiPFgyIfPPRTeTOLTKYY9UI7XtrNWPFg0mIIMgiG
BgJymFrT3HLbjFpvPz+RFBy1n9zZ1sEC7pN85QXsic/jvOB6mouY9Y3Jrz2qGd80AgSV17z6zSs8
BxpCCK0PZhrv9jRTGpO82JhY2vibUn/6+gSdHFhlgyIHbpI3g2U3TYfyLzgu0FLbfr1ti5Hxjzsv
Ct9QsQ1njAzIxT58JCAy+jpniWnHSSqzzV6M+EL4Dn8oJSVtA8+TkAF6gMzRt8UZaOUjsQylmRrR
waTK5O6899rsdn8hL3No7AUBStVywEO3wyeb1zHYb7SZ32j2rtj1fZfc6xBT/zSSAMrgKSYY/cub
fWGNx8kRql1Ui4g7JNyRxc2bmvYU2KuVJeB5BeRYOyBKjTuX/MsN7QyZ5TtpyvUf67V9NvHhW/yR
ia8eIj+pgWNsjd/D5lFjxi9bvLyTk0kcPndKApTsa037DYZp35vi2WGcI9aXbCJWHSUJtPtULMAu
qOyVErPk+eSh983YZoon+oyAcrvrFjgCf09Do/S/yaZYXMgwADHCPGCqyNcCvo8EMa85iJG7Uu/n
Pklzu8LgRuBO7Q5zGTgmy6aO7U4JpCXdUDmTLOjtPTg+LS3px59dvMZj2VPbWg+29H370vElcr9Z
BwXQN+oo68m+jKh9PfcGR0vN3OQKwScdfEoTfZ/+OZmJCex/K8cOMqFxss2XpFymVY29JAnozlF4
ILJjBBlRYZcagqWm1VgjKX46TxC2RXsEDQKp032Bx3JYeEYqwE+ad5Xq4EycOkIUsPs20wXPq2jl
+M/QKMxXswf18LAcxy6fZ54Vt1F+KV/Ag5wEcvMev1qriV1lUijx4bcy7h+P8wz5vfLzCbS+N2AP
HJfCpGbCl1Jrw+yBkjGdcUzjcvo0xyrsvgjR3Wldcsv80rPSMFFLLHInJYcwx/ZSJpv1w4xcsI6A
kxlG7PyJLXUFVcvzU/afsu+eMExqjLV8STgPLjgo8fL1icqq9Olu96DVNC033OLxP/tPW3xvgqSR
spv2QFgKu/z1T4Yy/DPb3y2AK6HQvQ4W9y4sIkoQdJvpfkTtASsoG69o8d7rY/Sb7NbaPx17yps+
KHM5cJyTcxUHkjBI8Lg4+hACIHvyBBKdtKhWwpkAahEjP8lH3/b/r+sEw0AwwXHoBK88myIi6UQj
2uD+9/oCLGyY+4RqEvV2EFUFT9pYtB3FdbUARwcd1QWP+aYxpUIx8nMveACN+4OUrr4iKY79WMRi
Tn5N55Eu7rDAxU0VGZhllVJx1PSxHh/+UqJnMiNekOwPwcLUM7omDNBtHjw04IFxUpeKYCt3x57x
VXZb2lghDaZRa1uZhwrHwdXPmmU4ssM3riAneuB6IawXd/bFurMdbhe5pfhYoRifCvX91wtDo3e/
Jr7XhKZLrvQORN7SxniRoqgxC1eAV7O6C+5uaPxySIXBhNX/c7iFEbPs6n6ueqY8PUAUQYwQfTCj
JEE+K6QO8v8m7/jU8a7Nd8CqaNF/Rqw9FoxQKNAKX1d0IspyFcXl43s7KKf6TwPSAgZOSnun8AAn
LBpAoqoZGgNOaaCVt9t018eHnPtd3gOTsqyej4wDy6bqpNKhv5DdxqKG8T7EjzYQoWiILj7IOYEF
vUSj6+UlkMe2cbmqLtOpqHm08bI1KO3lkyOzXpBniPzH7SFLU420Qj4KYbflvP/Q4u9T7C5allKj
i40lBg/2Kvj1HWwwI32xDrUrLK4RmQ+JOzItyR8ioiHkTDfbfzcasWmQpHD4GELrQnQkXmI9GFkY
3Ww0Z6iJT0Qet8MBrfqZUISf+7EFs3FT85T5Kdc5d6Y61t34aShRgXxL73t9BJU5dVNa/IyWPRKw
vzKPLVFUvwUTqh90njO5fGqstoVE5vSP7CKOb1NLKjjND2U7v0B0SWrdfu2b/0feZdmsm8FJMaAa
9j6uUavYqf3xGk0WKimD74Sk8b/O9G2zxsj70zYu0i8nMVTNg6p56tAws3uVYI80rVLElxjJtYAA
rdRo2JpATiVcb61Xs8djS19QsYA69p+L1JPFz89LRXFhcOdiIR49X6wMNzkga4kKNpQkmwLetTgk
qjwtzyB18s/U6llbcPxQQv3q8Nd+D5em/YaE+qvs995HoEKUoIuZNvulFQ4qQgZX9EYTGD1WbW4j
rQ6olFM20cROvP0pM5y8B23m5RZTfzs1fMpHX4xFEox0gti16INyvD3VCZ0ZeCDFkE0wy9YhPIhk
Wd/9gsgfiXm7zGB+c8hp7LhunNJm3vFwjOUPfhkY3mJ/zcqMMEucDougdMHutkey370lJxPuzzWp
cjxsjNFZ+fOGoT2w1ulxuvJmvJcEDsqZkoeK1OvFgkO12f0HXi9QgfPIz1ndTHxWCneBd1culXSi
uPJjtPw40qxJTu5Szmvh0CAfi0UORMxd5ZNchwTVo15YZJOumHtO1/N3Za4HXqU7Nsra/xoah8xo
DMNG4ikqyFNFacZd/ceWRqMuDQ7lGd4tRh/5FVCufRkhfywZzbbLf1QE3r3ncpfPbvq4z+wqy/8o
j/1IqYaDzQWdAj5fm9E3g4v2OrmIgHVX7euDqQ2BKCSxBXwuPEcf4HALBSutTmq6pdvWIqII959o
sOEB5cykoFhPxrkq0LySrLYedfSqDBl3simNpcqlSV0T78ZkIMR3ZX3WSJ/pCA1HiIEKY5dFNgrl
RFGFv0k7JrrllxyU5DhtfuCz/N+v2fsC8yiCugDV/dB4P4ahKAPeFg3h67g+dX+HkAT3Kc1MYzlP
Ie/awnGbe29q/Z17O8WY+X5WD5oK++7WSuu4kntzVivohhCet13eXJ3OFr1C9kDTQfWvlaPc1mxg
s/8uHB9ijNXMyCpKMmgDWmNWd2Gf5H3ElVhjB8k7GuEoKyc2zjsQOnLoT9MXm9wr6ZK/+qtLHaEv
k9FpDYGQBpyVAbhzK7JLahaIEytzBsAR/K6gk+mt8KSx1uxFxZGpj84npPXc1RnleGLka78tLIsP
CCp/4HDgYXYb2mjxLaXPkpxmVImzBDcchNhtNee4Mlsig3hw6uL30dezhBABjIX1HFB94RmxcZrk
OVf1sLzXbHKpxu+kdRY423ud8ApryYBCgyD/vW1lZj0v3zU43wc1zKfU7tEF75GJ93mqdv7CcoNe
kVVeLS2/UkWXTNTu0cac8Y643oxCsgu30HDLiIb+kt27seBCD2oHAKrR+b+5KH7NYBQz+HrG3tR6
oVxZdGAN8imZGb6qYjOYovdbfGJK4ZzAv54cEN/KXKfaAgP50oWErzmkZ1d5TA2f1ykO2Bn4YvDq
kI+PtllHU9QFwLBr7nmFt/EcCzWE1xQC/ZszF7ZrQgzQBaiwjRS7aWkLyRA8cWQPyTbOm+L22K8K
TDdykcCjBceBQgAftWnT9KDuLwx4F1PDj/8OwmrfQN9wrVU1SPsPjdcyOsF8zdRWvbMv5jRjMii5
9ZrepsDmvDgOju2gl9YXEZ99EOdOuopNAmPt8ctEa8dtyVUTRIY9NyhV8WwVmRj5ZbUUOqSCYvBt
Z0Mv/98HSQao3e/oiQKxAEEnHvMzgtyvURu4/M5hVvjxkEI3zz0G5RYWbBWmPoEU02uV+RDVedBE
RBPL8TGJoC+yAPAoFA/hdcqXZKXZXdWbC/HxcrwaskjPvSDDzxYLeKXXteLiix217s935wnVDRS4
gXoQzM/KGCX7+kmxxgXHYxCIKERYVHv6HW7eOVTvpJdddu1aj1awMbwUq2iSVq/9vtVY6WwRD+r5
9K/gLCGyZl7qLFPNKYWyTht3jJSnhGW1Sx5JfEBZiLg7ZH5l6ZGK7vzmOT/+XCokVpnL30iXBoO+
H1MCSbkeB6WYmv1bKj1ET3oWBfdkdS78yzbcOOF6yk7euptjeSygX6mIkMLEzUmE9yxuoASHlsp1
o5q9Z/doMpcQIS+AMe+X7T1eiqodt0Px1Udztl4CbwO3GZDKy2YLT6RE8aJvgCC9G2bW1C4I5sbK
aPL7i1FjSN5MLzzCQ1b2pwlxG6+UP1eA6QBiLToqfJ5n+9UU2XT+g/ojofp3CEYNLQBKv9MIlpx8
CF8156Xkfyv1bKdhS0QBUfqZQuJJBhYNjs5grNkZrJOsL3Cxr5YUa/aWZGKr3EB04IzEwDtuW3Yx
Y9ZSwGbnjSfuHQ7Z1786245H4EVjVceirC61VUAs9vwf+DheJjUtD5mDyO+6wRnMOEjcgW39W8yU
MYwJb+VEza/1k1Nn3mS+O2Fv+vV1VKXONkYUVwS/WVpmJqSz1J/qyaH1RqVXWsbJNXmzbLZSkUPK
bqKtpWb75sfk9EN132ir+itWUJY91NNNU1mcp4VJm9yq44g5dw6Mv6zJJ4uKpyYf5bEkfhUHTwI6
Rt8btWik7cwKs+bleGuLQpg6djMHKc/NszH2w6qXRmilZLKFWYhfqAORIlCYqjCRDzD8qtCqizSl
aQFRPiAbPMOMpyY6T5qGFa1G3jgUpe6KJEp7QOBH3fUNj70ZsNdF9CLDMhVTtSCgk/njUbE2J1V6
RGlnQTEEqo4bn3SiMFp2+jMrJh4f4EnF0XRnhycqI+qbueAqlMY5YWtFcpWopEIno3nAY4+YJEfw
FD47do+nuphdV5ik2Zpdy/a12oZCqq3C+vcRh9tP4sPz8wgIP5kAbbXHmZF7i3Oc8NhZ3kaxob98
smM2LnbX/vP/XQ41JJ6IJavbiRv7Y9LFjop+F+cXHihAa3TFNlELvYLPZoXynzZT1rDa3Qy4v2Kw
MxJkhr20mxyPNJJ+hyTMrhzChT+QOUcdQGv7F6GZc2JTTvPiLdRDsHTLjK1qiS8eX1JFJUdJ+vXQ
MpbufuxKMNN9s4/ZuuaxyZkUMJKvF+cpcvWtfhIJzgitDOA1OnJWiEPc3BzQnfvM1gWEIi76W8gT
D1qpbVLRiy8KvppLJhNGhQEOK5mnpZQPyPw0w8OtwLUyV+WHTh053cN+NBWCTj51M3k+nnmUkMQl
ZJ5p1DD3eaw7oBsHaS6ar6HPE/kcQ1svjNJMb8VxdQjXnwULxmEHh5PJtxjtMzFvL0liFkdYTeRl
LqbWp97a9ua9JQKpcDPbJPjLjJXKuwG/DPaExV08LlUflXlF4xBsB3HQv4mEdOHWqOZVFXnY+SdN
vbRQEiIpPbDJddHld0deryR1FO+zC1F9dXVRhZNAczPwUL7Qm0qP2jT72pyX3VGIyj29Lqq7FB/0
GjBjwSdNcKifPtcTHCyoV5wgn8RTsGFB9bcpb6SCc4zWsdxppMTh2my1kLM7ckOevi71Se7pIyBI
lISyoCHjsjOcFeNae7I2iBEHb222z4EH8/8Y3E1EuEVTlq5IRIqYse+srTUkBMaLOdHKn4sMDW7G
8z35efLt++rUVxva3SwBO29hX/D99pSQ0LyTgTuf4e0l5nX9kmI2oNhVdunbvaCbMSC6ETs+vdA7
W90M4EEW1kH3ZJEt0DmFeIGqMQO5GNIiELawyR1wwA/3FHHPo1T72yUOWb8oPTheUOy432b9jmyb
3cPQxOyvt/67gVudL0JeBFXMjpzG9qy7czXcDsVWXmcYvpR7zcCuY7Yr2oZzQEp0ugMd1qtZqdwj
LXwG+w2FV3w1emrkw/j7velzmUvnU1j1WQVETL/G0EvEvd/UdGGBA4TXshSX485hRqjFp4UUi1d7
ORjwlFVIWL3haE71FH3VEYGYKMdSYbKLweu2onwSTmK47oRWXKtjk+7O4iGawpYfRCMmgbQ+7XFB
aL/FvzgLvEk2l4qrtODXzAwHYReIYc7UgNbRYaBMOFAnm8j3aCuTOc/xNjfTFfpFypxyDR1GFfFP
H3+7DSx1fE6S3ji5DJTWItHiq0x+e8Roh5w7IZhXPjZNBHMurm37jFgcbbiFeiuup6tq6DYOkRc+
GIVaLckZwZtsA8VGcjQxZp405x0jR7uQJ+gtSObsbrQRP3yhzSH1yi741+3tOLdA2LcmnkNIplZr
d5GCBYbMHbn2Xv8uBM5phs+GKgHWZ373cynMFbMrbz35UrJoPep/ChY24D9za6xtCqQM+5Odh3HM
R5LTyP91XDuanGa1ZZa2SEK1GZhsJUSQecaG5aq5H9UtX8JxVsagiwR4HzsE2ysoJsYFBozN1Eva
5geLacUaz65WaFFm+kwGYwk5V1+c/5bFOBimBX+xlZb7wFvk5SLiF5xBzorozpCdFFohYNfe8IpC
DLc/cR4D2HLyUU26I3T1btUBZqpQnsY/VDq3VlOwXUBHzc9leSRj9EhO4yc5ZPlX8F8UiM67hn0Q
WyeEv0dFxpwnXoBpYARYtqY4oibLCdthybYh0VhW3WL6e3REcVpoSbYVoAZhYRWyedXTpRLY7ho5
fZu0MVwNel/MEdCJaKIqCwReyev6c5REkIIGXvFZF8mZ1hKdtdBDFE6Glmdc2fQsMKc255bmyAFO
29HEeFJCxUBbhSi+teDygYfcuSHBmgkSa7ohYFcgbZX/+nYxQKEG3JceegNopfxPcX/SllHJGH4W
fGiNzQAOebY2DvWPGf6vmLpuqUHTOu39xUHJHEzcbRiLGI3fOqn+JdG7Sic0p6PFC/gcRccv5SM9
TS+dySZA1LIWJmPERzre7yS+5DcyOUb12WJkUxRz/3YA+SV/7EgykA59Z5KvLGi+eweMY5tz8Vea
6/LuqpZh2Q32fEwebmztRmjWwV9VhaFBRbaSAzdIqY/jHcllhN7jSWQALvuK+xth1WD3+5SJ33ae
1hl8ODFKJxTZptGa6Mt0GbO/BhFFUe20KtpecpcQpQTQhMYN58YLdJUU6n/iCPCFSgES4yNif94N
q3O6mqDhlMeFkYWHx3SVSSLlgeBd+Q9C4Q2ERpmP7i224v3U6SpK95zVArmBNDauYcoXGK1EAk7E
gB8qSFRv3Id7u/i+wsk0hfNWjDd7ltTcpkZUqgwOxnmlB8Dp6s9pV8rBKcqwL5cuOkA6hoZJ65wg
AiFvnUTP3+eATvNVYysHiXsNZ+q4HY8jRhyfr+iEZsZsV79RKurFbUvpP32Msmi1tuG9st3zwGwJ
bWTc+vL0o8KquYmTXb/f9qCxiSXp1xCf+QfxD4tRxbuNMx/sLu/uRxnWXn4nDs9GInKSipAdKTGh
bl3OMQLu/ajjrxLiUv0CmUH9uVV619+vVNM1ptcoogKErAghDJwAnrZMcVLXsN5YzoNPZCIUfk4F
ApDGbWFf0JUHNkYrns4pfM77aN+iESOHlo4wnwrQUyxLn4+SbHkjBPeysnHfJ7bOOarZnZonYcv1
z+J2nIst74AL/BoBfRMS7naZf6tfLdbq99mEJjUSx0NembJEObpI4VMbAI5NkWTi8T6o2WxTPCVs
9+rZ/DLn5rVPMwqlmx3lmuM5G0r586yXBv60cNreow/oFJUX1eCBEWuYksRQhN/ENKXIa0C/O43U
HyQnAchkz7aLNkOWfA/6HlhnfCzuKHUw8jxzpy1pNo/JoqwNHssnh5+iEpdBgeYtvwYJPwysWiil
AY/Dk8aolZZmSPN4Oo9z0tt2s/APY3SjDy7BJgpfJiy1GhPTjbCoG9bxcTcbi2wBEriC0DQAZRew
+7WbE9OegWRrLOUAx5cqteJpbngM2wXpmkXVuRkgl+OXpHH2Kpzw9tpoVMgKAFOwsATXq3DBNDHP
tHzQWpE013gow2X7knH0yo0ER4UKeH4WzcNp+9D0bnNYFoDdzO5l8BQbKq3lBy/Gc2QIeoQCYKie
SqZAtZBfZpK/Y/usiaGAXRiPgdNIX+GzDTLxXyaNJaDbrFdLGWqYxWaZhg+8JawSMwDDPRpm6++5
GJ1UahXoELK2Ge42oUAeLQy7YZiia22MueXozXfvfVxPK0YEcQzeKkKjSdL8O9JZ2H9Fy4TjKdiY
7yHRhh5TIrg7ziNdVsFwL/mfYYtFT06RdsYn4mKichgLsZJtC8CxlMp++I7ZcU/N+aYa/gbwu4dz
84rI5AMvKwVEH4rpHczY8r7Eyru/z2+9FvN0pesBGNfk1+phyxkK0UdGTEjlFiVOocrWquPaiizD
wtW/HL2o6nJUbTwiStAbtB2Z9HY0sBTEN8T2YULioNoK57f/bFoXIdcsedbN+E1Zgggf7i8YvzzY
cVjpINRHiKnsa5oXJyiimNYX2JKp2ILszBblwGuGFNV1YP5nC40XHDhIhpEhL4sCqWnfiUNV6elC
Ky/teeaIPpM+ePGfDBEkp95aKw+7twpknR8jVq62D0zjr6dJf5c+57nyNEnDtWqUDFo+fbILlfh2
ZrnVEGu/rdpvwxE3ZQ4ltPOtkPkRf1vr+Q7I0VfzglXsXZv8IZB3+hFD8Kx9vAg1P9zZIkN1cbLm
NAPPJ0P1bNHMQiYCc9vXTLErrPPxPJGOQLmVB6xvuyQ5Lc/o8I7vkrjix8y/e3vCXarN+KjodfxH
3W+KcuVj21w4ML+rih1DhpibUdXboBGMvxhAo/yLVYcYdPtnoKAMaDtDGGzrh7r/ouaEYDG5naoY
iq6qQAqNbCjIocy7v9x9VpIkxGkVBvwQ8nEdkw7+59QjngMydl3wexe7YlhNYIyr63Ck4WwUClZH
ozMGfrAL8WBwKVZ8Jqoi2OJWHhCGZAYTNqbgMEXiCC4XensPSlvKx5Mx9yyRxKHQb+7IWgjK7/Vr
DdbdZsEWgX+9/6/CPwnehNvbnocZ0M+bN4BFpLSPttn46BS8x2sHLWiLIgV8ntsBfx4L6Tmjg3oW
JFuUJAryPm0taTR6z6CRuHGf4irHpIovja5Az1CuInlROTwqaIZ2l/X8cLKe85kTgHj/EnJUuMf/
WcjYeGLZjS3S7/m5CH5DaE0c7P3maYTfHCahz3PufqfhzVgzyKl9oMNcvLWlGzISuxeMceSpK1oh
x33F5BnfZSK2M+ZodlobsB7jGDD1zxzJhjlTEUNxKRlsYMNsTkXoejyHAPDzVApp2Y7dOXErIXF/
MXHc8lR/HWUOcD8pFzo9bHfyyEsn65aOP0RQUVpho3ldDq5sgOyz2e+hCr8POB3fbGQBQluEXFEk
DtXYoryJ21uZfm90qdZBG1AWTA3tzBb7mKj5vxVh7f1rtcZJDvaqTzjULP6psNAxTJZAPL3RQAu2
OF8I0uyXWcD104HMV04hW/1cDmS4a86e4byrW9RocJ66oAOuLmJvZWtEytu9KkotP4Z9JBDkaHMF
nQaJRsq2ZnBiI3vUq0LLK5o4P6WHUipcGTRhykw+03CwSurnAo69cHnyvmH2+nOiMa+8hDR8vtHB
nAtVb4gax0cydUzFnYwbZ1ivGdyc5MWH6U1MpvOSXvWnaCicxH688zEgatms1DyQcUbBlgjfyknh
HzmZd4oOQ5x4ThdFGdHKN3I3z7yDHI55P0Mv1uHdI/aF6f0fZLMZt/ZKdzME7zlGqLCaNceRHTom
IXMSquy6SiCI+xB9uCVnUICQPSl8TtuyJW/4kpP40z7uW75B1Bwhr/jiQ0jbzxbckm/NJQKmv4wC
evir8cHL9CdSQqwHDuwjaPAmDs52cSI3lQVQayZyuHGVi0b62UZRVCH/QEEiqX1+qOAj1bLnJjIy
OIiXRO+CgV8R8gu6nc0FqlZFHO5AMYrg3W0Gq6futyCDDi5PFnM3LZNtZk+nWpU9eBSBMkioKLml
fkQj/ZqQPOEmUd+cKCNbSaeGKzUcuQVPg2d109E+9yyABxHhEeTPBb3ht7G703dFdWqfKSPOuvdZ
rEdKVf7NWVnbCHlYrH2ncu/tjm/YLX+PDC1m/VqFctAUMcsf1sNz/hR7dwM1UdKKPGrPWj51NmCO
yKSbzYZc0Ls7byBtfj2qkB5swaPMZEBR5pjZzBcK+0nFkMH/XA5dJqomTAZDFV8mYh/39nbZ/sBB
OaPeQtcDvx6A5x2upxQsoB+1kZv/YOiYcZsC0AUKh2W0v8b3CJgaAPvQ/D57RMT6DO1R0659a8kT
NuI5i2Ks8DM5FVST43qwk64m8BKTU9ID4DPKjLZQVUDA9yJr+LE6QgGw0mDi4yr+zvuPJZdFKpap
xc868Wmbc6D0yqrkFKFcx59J/9oLQ5338EazyxcamhF0czZv8qsc4lTMOZIEXdfEFYRpChbS5akR
4kufUpPcdurqqZu4OMQ360QmimKM7ycuQG93x1Mo90ZlJF279/WhcBcXjDBKVrSCAGWYnwAyk+Iy
fX9J2Db9ZF2ltKRW7l9yBCY/L4TFYw472HIjM57Df5pzjxIo9XF9IBrNBti+1H4+qD2jjHjOe6UO
tW3wXn7f+UBUCc/stoKW5fDyaYf2EUc+xHtGK0/v4ZV805y1C8lAGMfzTfk7+8O7VFMyOs4Djc8C
lNNthgnRXMVEw44CqPGaTqBgNT9YS/o040FKyFH856z4F1loaJHsmU9WeA3pA0X72wOBM1nYEEF6
2DcnHtFsI9zos9eUOGvhsvdqBVfL9g1Ls41+nkF0XdSMWAqZQOopd0qHk5i4nicGb+dGqokzC9oK
B4EBGJxAzkawZJs/nZWy+1POAPWhhTKRzpNiyKmi1qX/l8o506eJ7R8BBzZMo+b+Qg7hH2pThLjJ
gNgWapP4jbSbYONiRUmy/NZmF/RJtRPP70iL4HUL63lnUC9wOBHMnnxsinkDaBYLrwHCtdw7Fk8b
nUSLF54oVNx2Q/quxjarJ/s8FNIfP3Aod4mO67DTecj5Nym1XWpAz5ATuxTrScjEllcC5qrOCrgt
8HV8hnwtIzAR7bC7819pJeCYSGNzDwnQCrcMVwr7AEZW5qk3MT0pcwF7SqKmXPigphV/mLAfNvOd
4dUlWlepTAaM+7KsrT0wqAWTRBLorFW+78+Pm/FrrNKF/Ycfwb7MgzCwsEbdpR0kmQRpT+Txi8h8
IOTqE8oovSZX66eJd0VdtzBmd2HPiKJ4bcs/gYxwcQeovenfdmulYx5ye+vE/Wr8JmwgApg3kR0V
GL/qWlSx1MSSwDVIbZ456ZfLKoMk8aSMZzqysiC9UAnwdRl622R+wPFKf34KfAy/skCNj7fuHLIK
I069QH14Oq1FPkDG6lNsiwrEZX8yNTu48TdA6t7XfYheA8eBgAuUTRZabnDiI547qw1yxwV+j5Sv
uk8SGgoGbQPcH4YEqk3pcyo3Ott6UIoxs8geRNH31xvqHEmS78e9v7f8tOGsndEDpaa1lp7rGefW
lqugDwJaipCZGMS8HDkceYNbLOmz84TYfkxGcuR1eAR0oHDQ2TvNb6UYV16kQtystcqMXSoI/1yL
eZhLzheL+Y9qGiOp/+hUMXtEM1Y3WxS6Nphwk84j7DCy9HJUSN8VipIsecj0uWsWwdGMre8XzWqO
sABDAhARjnWB3+Lcl+jiqsy8F7Jd60iKqgJSeEGjWelHD5tMPoJy1212UYktmJ/RPRgjCWVdtWQs
Xuz13aVtvS9xkG9hy3LUUrFtA5m8rRDc38fDETnO8kdqwKmcuVN7Xj/QlFRJAqnGNRnT0enzWRpA
IXjScZITYCbI7TbdG3h9wT5eqVLlQ4vMxuxa5jyTZ6W+0XUrOf2d4aerK+QKeFs3xz7gS5MuXJYa
kC2d4vMkpc1WAuwvf2buZ7owhauRoOcZjPPGJ6drepEikYEJN3QkGKgmsilxQqNuDBkQxXAj2i5F
lJO/DwgYiCeMla7IUYQPx4tyk6tzKaCwugwOPA0iRknS+6pI7VtcWKpZUBc4EdgRHsWbhfKlpRuI
TiZ4r7EBdZk5x8POEsboOMCaoGHwUwuqOoTuwY3NL/5Vgyu7lIH/W2GeECLkJvjYKNu0oM1t9aqD
FE5wy0d1pRhEPusCflGnGFdY3NNXPva01kcs39bapgFfL2I/GCb7zfl97UlfMoVss6TAA/QnM/nj
OORTQln4l250jN3BY93Qi2xYCCrNtgXg2OHxJRRQGCyu7nuFEBVrRBB2ia86UwAy6+9yK9lIL0iH
bUUhJQS49QGwl6xUBpeiJbU93p/ffIFlJMHf9Hee7PFuHRtKAl0SwLzlQutvUpiFSBB4oq/Ev0xA
n7aZfYicdUNobc0Khdif3tM+3UDp2n5SNFN5P43A4kGFAxuFOv+gEIJ5N2gCUZHGYN3qk8Md3ljk
ssD6hEh1x/WbSuFrsMWRi7HNfMyFUQMP0HImFrHz5i5HJJy7PxPoS1tpZQ/ukiYacBwdHYCZWe0X
WwtwC8Y5ZbJ6ScyyVWKn32dh2jFb4zn6IWp/6atK6H9KtMbs07vS+TludfNy1BXzurvt8elAJSx8
40VYjfmF6RqBX4G5JzBfXVjDtPY+/Je6cJMiByWPXyoUP1A6tOnbmh22uz+yVCUcnUpW1cQ8LWPK
T5GlcvBa4mESZjylf3S4yS3X3bxKXivFFFjKnO1sIgWUyFF0B7bb8BG73yvE3qC+k4YXlw/lVQXs
5hI+s394UV+mH+XU4vD/sG8FTjnME5NvlSIbP8pxI8KM7IMVZ6VQARLepJkNwy6/FBKWk9304ZpK
L2PHz5zS2eG771lpvOi+iZUDL1xp0uI22BSE0Be+ncAmX/cMMtfsIAgW5IDvm106G6lJ7emq5K9t
7DRznw7VbdDUnMMoTFjtdxBaFNywJQ8w9P1Sy8Z1hvxEFOHBVOjdYRmnugeVxQlD6w1SJk6Faby5
i6usVWp/O4G6tdhxcsp8MsjLo4iH9KDockDjvIg1sKMIwpxWyafAg9tTUsC2dhwOUe/5Xungs8d9
YLnOYkuET3XhHPrPRIFmzlDION+STX31TutRZ4W9BoXNQKG5rDMVovOCn2dPGr0P8qPZlso3kXq4
4Jf5tzu7qc8V5Ga5vvxbsAb8SNQVA88tO0jaIpvAcQsYN6bC68klwEPAtLWfANaw4CmVShsWJBKT
+Lic3KNYtMLU6x471ODdQbvNKJ+hlFsXvsspATLerAA6GNNQ8upIoWM7PVyv9haB8m5sdTTxx7Ul
WKH2mLlEp5vEUT+o8hMXm9a0TMxnRbuwr0ZdPLm7v50+7TlQwKSF8BzDj+POUIzAtQsiNJ0Q+G6o
kZM/4dcqVArPZ356oclxy3SkGsKUV3BKIYWrWgC9hsm3V+PbftHqFwe1frpQfurYrwvLLLSjFFJT
nRb8Av1iHP9xE4X8Kx/6DSu/4j4f7S8JHEYtPSL88SO4RiQZajdd7b40RK4wdkpEMchoRu9JsDaO
beZ/s3kKDHCeI6uOJemS1FToxX8cEdo90M2orx1P3QjMsiw+R9fqZiBudRJTUplFUeKDZQfeNtYF
1a0ickkO1JUkqK4vJkL6isI8HVHdKsJw5lOpz4aLhCO2UNLCRPeU0SJM00f76NEzaF4uYw4zh2Dz
dzIFHf5Lw3wgcxQNSX4394iM+tutptyRdvGjmQXMxNyrJKHangeHQS4QBp0jtO+yjGv8W2mE1Vct
z6VrdISc8Z4Dgb/IzTaD8tXq0ohj9C5LTIieJzl/Pm17IxlpVXQRvpp3Z9jTWbwHBOH5SQbj17WJ
Z94UgeOjaE0538bSzqwkBN7zmcenFtxcCdUB1IcUgkxjNn1/hSJWZbt+L01ke5eZDtNyyxae/BQz
AsBGOhU1QpDH7+RJx31fhWp9JKvaXlYYXCXKOWsiJ0isYnMy8N3m4OHHToqTd+C3Pv+XWFidQ+Ki
08p8gYMjMB8+bPXWfw27YWjto4F5fMLhtVDbN3G0xxjDqrIZpzGHbbnzuHzqaa96rW+KimpVm5Dq
cMF8QeeZMfl0fOTb7QnkpiSwLf+hI3H9cYgObHAz2p6imXSKx4UVsmvwoLdcn0AhWvQ8uT4mvE7M
vBzEMBUJJoQf92L1WohQRpc3dLWkSDecgPBbmtGGhCClH2i4xq7p6UIp2qsD9EiXIdyA9XkjZNGA
hnyIAY6AxBcWzt/ICWwmxBatHDKQSfA0A80y7/ORIvvPKPLH/RElb8KiIBcZhHlvPehgua0CMtVp
4782Z/UksIsQ+dLD0NTWcG/XCCttOhHR6HHoQ9l/WxbSKSoj8GsRVh0hKo5bE41sIyGwlSRwJZB9
dwUKuWFecbJqgmRiJwzKvpKY1veUwuqnDpSg+JdEUJSAJGpPVf3NRilNOMxGyZ924ApEr/P/+8qv
iedh6+O5BTYLmgGpkHp0MsDTy/CHXy/H7tBYPtQIgxd7H5CT7NO6kF1RNqTLBEgoryKb47jQ4lKS
66/24Ar4yu8kZHFa6UcT19wS3ax93dzG0WRkFUgiPu/GhXhFhzvt2Ahjr2Z+tWJozLmIjiBk5nuv
sqPdmTfe1aw6QyNxHynCIYm8BN0fQ/vx6SXL8+Jq9DvdHYVKx5ibM9FIw8dy79yajeQ9XumpR9G5
igEM5Ma5lrHDJbj7a1XouyWFgUpR+mRySNCVdCjJoA5hqzly7FJ/cbweKAmv/W4yZCOj67nGK7MI
n8d04u0c+QsGh9wwvPkPjUzRcvlWFC0QRURG6LFnvjTIv+3moL1HTOj7MOGlNwXHiMs+/hGGxVX9
Hg5xqysPiBeE0aZ5mhNUggF5SSeLl7pPXIjOWlcQTH701AhetktA9zLZuXorg4b5meB2+mCTsN2R
LOEuZUEYHJUSdNu/RK5tfOhhztmC8T91pQdWcrLdKX6nx8/LWG2a51ejZhkRjwOgM6/j634Ke07O
0YplykTxfWTmkg9yKkkHUWdWqmVKzGHmcGIel2ocUXQ+LhNNxdpApyBxcNssZwQnZedyTPva9iSM
5J26KvKHy0+GrbKC+uR3aZNPCo8iOmfGQZEo/xxvimwwNMnFQW0/rfTOEu52Wt6QnFvzR0i65APC
pBg7HGvQ+4CrhFtGlh2A/wkBRe27OtmffgbsdIQkU96KQXQVri+j8o2a2m0BxxiKp7e+6BjVk4pm
QjDhseCtdYYfMFneVkl4Tvnzjxn4e/IqAICO1EvbbswCiD6L8oQUVMAsXKkYFNMjULCnpk8jjaMh
MtvtH/9Ubp98POXyScV84rFyFtFM6dziO35MAEfH1R4NN1uvfkUADwWW6Tt4xbo8RW+lAQCxiWEc
6byXkvSGsuxUdu61PvYoBiTCNPZSB7HuKnbLTWebRUUfSvPDTC/8k1vCYWCTvXslTFHCGFXA1QlY
YK/OkPlap/8hmnF2camhPbcPDiMXuwH55tUsTKmad0ns5PhIb/Te5QmYIBPY9oaVOC3DyYFgbm6f
MJtkWODKX2kC2FJtiWUiOKjBZch781vUk5mEApU1K720f0oeqK8ScnHbYgKTKTjxJvSSV/FZjcqB
I5td2QuNUFeYhHJ7Gz/gltHhT6hw/nldZM64+w009yNh6BkDSLHatobpI3lDG3SJcew2rjtjaOSF
wYIkGumFg53ZD043UpKYQQ0mlZncInrHk4/xzanw+CSpKwE8UvDf8gSJ5vw7rQMOkE/cZKAWP2Qq
cGXV0x5NYr8UKNDSZ2DeeSZU75GctISO8Ur2uQMBvtmJLnU4qmGZlLzKP7nx0ZFIvWxVfYMY+OWb
JGRGDfLeXrHMbnTUgm1X11euRby9FBOof/DuPr6ZbhbnLkgFbzDfkRiQGUti40PHEJf6TeFY5zMS
9oV87Mz5VVdvQaMkOORL9+XeGGi43Dc6NQ8NqGt/+vTzFCh7/nJFlkkp0i5Sj4IPl0a5RmYRLfOq
47xT1RD10mmawgbno7OWrxhYD6Ob7FX3CgFd937G5ZES9zvHq65Faj9JyfSXRbTZ5xa6eekUnAtR
8eD2KWOuD6zpqUGME0DtOQkuN457x0dMBvfzsU2qLPvXYdvBTUaovzi2JEbK3YhuB49Q/uopAsaY
nekSTGXHunI0aQcLJ6pbkqWcPVsqfc8pKIId99G9I+MMbp2wsu9X2oKdTjZ5rxm/JMfHX0b45EIZ
kKmoYAf9ozUleIJe59JZyFmCDFhz+AcWtGEVTz1xqgCyG7XD8DOkpLYAwb1Ge+e0n2AWusuFkfFT
xj/hO/PfCKphvyCpd1qm+UzfdlkefaEuuw2zTUkJKxcgQ9CnPUv9Mkmudv6NnAgIr5Z6wBtTB/3q
Ne+KivUzV6IEK0k30HlKWjlyj+uUG0xfQhno8bUZnx5aTT45hu7D4iWchXepSMQ7WIyDBSscGcnm
feQ2K64QD+4AIhM8XZwsRsV3fyXkbI3ZHGnpDLs7UCxb8JGQs4G/Iz2v7rWCIEWbN0I+uu+GjBdm
IBHBWRNaoKIDStmb47dzhQ7iDUaWZbJ60QbJ4H884G8A1h2m/vy8B4+VnjwLg7c8RmwLxzF9AzLz
i+Lo+EAIoe6RgWCJd8wr7vRSakoY+G+7qCzCBjramR13yEKIdJphz/wabEwsR5z2iZMnUSmNwoqk
HnBGJl5XMTMAHzvW/RvSpcdB1+rejKM1dIEJ0GMa51KPzLrK+/Ql+3P+ri1nl9qWAVzJETn4R7k1
AGwjbm6ddZuyUxVn/Ez5yChfX5OtUBq7+nNDokpowlPH496YsZiAsNkdU/n3ZhG2w8QzB4w277YL
jFe5tOcEaztElqOBZJtGgYveLzbbZG3H2KNL4nmBPUxwX/wdbXq2b62jX7ds12yVFnG2Zqcu1z68
D2RWC4MuqbFNmhM/xhSh9krPshF/4aEgmbZSW5Jv4KX/5M1T8x7CLBsn8nBSF3BPmxP4dTziEEv4
zcucGv1xGXWQBYShfRbY2UdLVAJd2PSItJ6wVpxB3n0t1H4QWlxL22G1dyY+pNqCIPYtFYTNgr5m
htAsrwm1mnsiuuFKx4GyXuSQOxNuOI86a9RnKCL1V6gALQtoXdgdnu5m5MKWwG5Sw7prw+9Cc1sT
W/bpweLmEZaBu6zFkhBEWIaRRDG2kRmS9Ij+fPEwxg==
`protect end_protected
