`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QM99PriFLrXtWj/tN0IsiXkm6Pgk3NhaS8nu4q+xYRs+lAuRj/dzQIEfFG2ho26711DjgHyMLsVB
GMIu7ojWaw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
csMBiJqFUhphGpJ8C0CZ3WP/fqe1Hk6QOrXNPqKtCjGAFdr6aTMU71aqAjleT8Q+0GJouQDZfUya
YnVCNapax4rPHxgQXvv7KdJlvurWyfZBMKy7h2cGSORTsIj8+5iV5jRR1MxaSknq0htfAAcGlYkC
UUsmg1cV3uHcijEHhXM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MpzgZQFDWcz5e/05dIQRYNQFbaNkTg//OxCQTZSroaQnfjLP5MuhzZL2mw25UtNrVL6c6Fr3+3Cg
hMd1lNiZsOi+Q5M3vJ0PCC6RRYb0G0aLKCKJhmImpW/mqcTJ5tkkz1CADc+iDvh410xIq1im0T7x
GBgDBJXSg5/zGwE/T98oNEl+pdQ8LPBqCXoMMcrrf9FgcQuPAPVVbL4uaW/hVd/KFWHGOPq9AybV
Fs/dYEUKCDXdi9FMy08vb4RbhbCxbOYeldEYuSG0NVuFO0ryFS3i2D42lmV5yf6fyuXUNKaQ2Yo8
lU0jWWv+8lZ+DVms0yF4aHkzhlLP9kj3JlLTHQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iDYlJURwKtDJOxS5pOVPSCxWkFEd+fZh/8Hl9Ol+K4T803X2Ztxnym+Z8W0HA3g5rCPCXc0gs2uH
rKTv0QY0S6rpw0oIM/z5McDu6VE62skZ2kme2PhVB0hqCpl0mTETz9xQ+MBzpzFCoSLNdkXrGznl
6YAptg5vsnAxOSnsXMqdyCy+2Eq5I+pGD4olf7sXdd2+C+6WeHgzZA0gwoPIoc5Hr2Y/QugDaNCO
8/qXr8UycIetJza+NSyPuH0OKIIkUjId3aVL5QrfeCYdSvyRy7pdmy2mGHRdNH0Gl/UikdUrG8On
eo8fXTE8N4JgLfofHv9FonPd9jEvJq3z7tJLZA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nALZRx1QnssyitHsTvpOhRXooEsllOceqk//PFkk1PkaDTtYKIJ2gomGCUxI9+vQnijvRlDgN61m
j7Si2FRrjkTMPeHLfHAAKdhys8SWQe5R4OBBm/GCfhX5i3xuasuX5EXnaWpgTKcMT/7qrBwHbNbw
POu22NCZN/XVMpdmG6MXG1enfQVcrmKt2yZVED3sO4UXxY0IlDiBxpL+YZQz4+oP1D0kGvxyYh5Q
zJl8Q+CSVmNSFf1qZajyOJgBwbbDJef6iaIJv9MeTdSRZLPHL6Eqlpn24qAKxEVYhRyyxzHieofU
VU8ry5F9gdcsV1sW9k/62iTNgjL6juSAG6mKCA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SWFYREqxRUZgeQsKSTLlG5+9n0zm+QdW9Fmyeqoumqqv11Q8QG5hAAnrnbAtn1sbXVGazWoFqxNk
DZzylr2MIdgL8NZl6sUyNpx0UCUg6KIOP4a/23rnfsp4Hn+2tmVDKSN1I7P/G0LE4HvPPUUm6Rs3
6NYO1zb29dX++DIQ9us=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dSqxWddcY8J+x+htmB/Q+MObpfG8H+bpNQ+0BGovkFGf6QaVfyGUnVnzqWqESuJkhku5wvfV9wI/
QB/YLTRReKyTZaxtbPvehIo4MNBQQHLp2p8b1Gsx++GWmpi65v0Eoias9irriitVXC+PJjasEoEH
rRKcUxMbCmEQCk/FqaM7rlNYlRQAz4NIsm85EnKOEtFl9CpmxO3Xc3TTU3sKcPxz4X3Tr5pC507Y
BA7LIl/TfZmLK5x/fz9tTYi9nR/+rorZnx7ZPEDGhxKAOHIuH61nM1f3fGAwTpMfkhwa0BLli9lJ
lltzVHcpCiQijR7SaK3mTIpKZPY/AENYtX3kkg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
srGcJ4ygSfnfyvxgSCdRUxA6EL4w5qzMjEuP+WGrA7EtcV/p4sK65LTpacK3FsavIhHcK4enS8Pt
KfNIk58s0PrkrXXESZua7CSUh6M/38w4KEoiXaBf9zf9mBua8k+yPPrRa4P363QgN3g3m54kZkIB
3jnN9mStV5B9iALCUPLx6OdkoLLN+EYy7eGjYvOd0NNMxPUge7q4QeNAQuAZP4SRNxe3iSE9EawI
JrOn0/FhdhRnDz3IhlMiq3OVTe0O7aketBaaIthYq+93aDuQTPEP1+q3c6o9rJu7gjquvHbEv5wI
IeBSfaAkF1Hn8vD55M2or9AYC06aqWKqspGmuA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74240)
`protect data_block
CO4TE6aL9QE5LJ4Uh2i8yIfpWUjandNsyAyj+bmdkcCYOClU3flZR9UfUg14DDJHX5JMxJShqmja
gM8NcSbdSnN14S+8XibzjiRh9PzX972/K1QxHP06Uggfnj4iNwUhmEX9Y/I2CYaLY5MbqHocE2xS
umH48MeactHz382AffsLljIR0zjb2fg8DLT4D79u5d0TTvLR7tQtLaknRrA/XDIQ6f+Y3fTAD1KW
/o9Q9T6h8jjUawKMc3JtybAPCwc9+5NlxImTHPkJTAYtVqkASrN/Qb0qX30FO0MhfEwTO+7b45Ya
63BxOzILKGK/vCNLfiUV2H2dV7mTLqSUUoknwGOJO42SYucLOQ/5FjInvqbrjJTygSXDKfUbIlh0
Gz/Y32yRK6StRFEC/lFCkM881Gsx/KSESpKxpqsFp/vrKbxDv/T+3pMEd2VEZ5thSkn7KolggVfY
IOnviDw3GB0Q2UcBADAXXg+GkhBagiJvYb82MXdfaN23htSSpeG/HwHgeuwJgOhIXUEUcpWZ2abY
QXYhG+U7wI656dZcwqFJpy/K3KWH+/e+6JvZqLMzLJMbpvLL/mjFQikYYo/hqFlB1uFF6w42LT+E
R26kBMD5gN/yPTicTn5WmJ2SjlbQTid+JGXyEFslncBaEHUb7qKEO8EMVjUn6H0vyNfj6s8txsl5
lHpf1tgYxumLbosVDv5os5sJGudratO4q5YNMFXU4jMSa2xDHHeNKMpD7Qfm9a3bBH1mILqD3ags
tdF0fEJhlR8x2gf5iS6pdS8xWQRjKsyA2zguzCdUxLf021H68drlCy+eeTonSoHjNYyT9tydxOOS
7ODirOiw47eZ6xZV55cWq5w5s4VXjv8cRV3N2UbuhzTdClofiHY2N6cQQlwLn1byd8OqiKm/p5mT
sli5cDWYldYWmsbznrclHTPTNnKtlKT9PWOFSNEkcMWZN917TH/+nhqy2HKh5wJFggIlGUARx1nM
yV7yUo5/IwQb3GJHNiiHJ52QoUrSyaW44pxHWoRpknshkFFtzl8CbvnSBVAo91ZY01EIWZ7WJ6On
2m2Fsfa8eWdAA+YaVSFJhFbWOfMEOoYUvH7dtYmljTmnIH672lLskf1x+VZqIzkGVzGrst23lna0
GqeItXKUcbiK1BaRw7tDZhRnntFVhhRsZCPrsUO9m++0QQBAyA5CVX1k7MgiXnDMNqh2HkBECNJz
IkBXh6JoLL3BWARl200TPaESQgK6xe0cgrQRVaXIjsojjxOhKwMvJIIG+pBvYEOF/J2Kg2U9aldV
K+gqeOiDuU3cOXkf26IibS66a+GPV1pKIluTEeeRkUgLVhuDWaWMxEgiOzUHIrCOIdTch7Vq0xJE
PFfRpmQ4Mt5JJg03PKkwGJv7xSNYEUtJXqm54bD2ccr2305Tg4tCbOd71VMwxjmSdTLYoQUYhgHQ
WMll/SMZ7AdSlVtydZQmMRppLqHL00mRyRPWfNvkp0cbBYp9vLQInUX3hlV+AGgsBjRPOHjgSJzk
FHfYTJ+ydKhuBRGuOKHuPKSjpX+nKZ+btDURC24vm8EvKobxIn0bT0jRHHFsjg2G/2c2hd41XzrC
ph3o2k1KopLwotgNvC12KLDKtc51xiZWWEQkZA81hum3FZ2u5obphmnolm/rZRnxNekx9MUvxG+R
o9jNi5ntuXvpTdag/sYm7aP7apIWaP4ybYmBLyUF2G5S+41tjCP1UN1ZKtxfInCWGanJU7Zmfxfz
tkg0cKjRpq1YU/l11u5PE3c37BjWOkqkE2KUWwqYsgjjJmRZyWutqLUGlVJl2jwN7lsT8NpleEzk
27KGBfuteKL4xbS2KZL8WEWq3cw/YLHfIQYFOYuRALiaINYTQhyAnGBTFEbZ9QdZwt3mtPrrgRZN
YtuYx3NzHyDYSneVXsVv3S48eWtNUR5vt+nQTGyOysw4rr7y/DSIt6XI79qdTHckhYc3wakDy6cV
cNRQR2w9rbwXaP+ypHd1O8EVOX11+nlTvot49ioFK2V16Ub8RsE5kY3j4lIi1qcqlKW587u5sr2l
eWjVF6SSd7hvosGXQ5wa+d42/XgjOuCc/diV1DHL4l/iHxyJYAv0HfVx7jICL8BKtYlJuINAQmdt
k+DUivcQJ2c2usp+xOHaGZbbNmJUhDJ0WhDMY12fhr6eO+gNdQz5aiSyeBtmLLm7TZ9t3WkWbzQb
cIeYDwIyapvbXEpuWk4TRYvffGDH0rjBdANwdU/DOITHBcii1wDebAf6AHPTwzybEhpGdeOrTxJ/
e6Og7G6QtllemaRdlTBM6dac23ZmwVGzXj9hzgiyHwvAshOl1/2qz62KGTVmBdR1f7qcca3+xXak
Keaf7WLJpR/SJmLwdfa6s/sXh2V68eOLqHaZh6Cl4hBYlCwplttbetnm5pS+IbrZNsuOJiJ8+UNK
YA9KzDslXqJl7qMmhG6guZKuQMqNtPI/XrmrMB16o+Fa1fsGAnyagylWUtz2cW82lYdMMxpC6Thh
wLjKiE7AH49q9SyNCjBoCldoYQeqAveqheAq6ZvtLwmPTp5I8pAYyA4zskoIYs5dALKjC2Qusfbi
l8tGXh5SPkE9A1aMM1BVejQk1yI1CUQ2XN50tA78UE5lsbqtDahy3fGXCvdOGmDvalroUC/Rh+P2
kbwGk2xAwdNG/Nu7s3DvnMQW6wkrDblMqRQzyhwkKiBNRExiax/hYlmkP9ZqCQx6f1Nq9266bGMJ
GtLZQUhRnvLeeC0hOiWtWPp0VGrgRYbXi/6fQkugc8d+BsiJXFuZUeWR4c7+ICBl4IMYb4yORyKa
PiIY0pwEQS1U7OrtiOpdkeryOYxwTCnQiDecXD2mYZlF71PfZkXPxHA9xbsy8GxE2IGvlrFNcLuY
IV+n7qQrdsH5QbMG6CAKgtu8+9uM/sAX4sPohgkfYZMfwki+GyHrWtWdh5Ik3wJ/oT90UOHkvxBR
VG05krd8wIk+l5qmhknc6q2pS7iddRmAfVonQac8GKRo5bcqOIYFt0TKablpC5nj2RVMz2c9Y5RS
hbk4LwC1XoxMV5BNE/i7HPFYFcCpmCBzjpTAPQbZearmwgMItSeOhegGrsL5OxwqMZFQVpH8Ng8T
M03HYqxT/c/SC+PrZt985VTxoLPOfBqdiorFBa7if+w0FODGLkeLNMXpnk4kfWjCVY2b322SYyyT
1bv0HmQquCuw8e7G0j3rmkOn++F+2CPd3H8foNiFyEzXcFF1N7kkyRzxFUKJdXiO72dm+KPqmZWR
bFmqaX1ooTBT2u5PxcmbylH72AHp57cQ0014pFmfBjxJsG7PIF+8co+9YIdVbQUOz2BtkgAKqEQi
3E1Fk8Iz56VsbYFXkCFwmie/cD6/HhiOKFe5cq6oC2L0F4Dbz/m3goqmGStuVYLTAtFM+YSi25db
eUR8kul14tg0zAswgHt6/Cn7rXEW7I8f62Q2H+DAAiql7YAgzLCJf3vKX98UoZBKfSkcqpFHCon+
lkQ6DpvbU90RETgd7/9VY+omG+oRoKIMPgqGO3RmedAJ47NlA3UfeYFWbuDJQGo/l5rKh4MkP8k8
ncVM57/kLrlx+GpNfSuhU1krhUf1BU51ADhVlR+RpKb60wgMFrRZcXiNAJwyBstKIFUu/snF6Axy
cko3VZspbfo3QQpzsSPtJOZpI72dJUS4GwOKxuOu5i5aIxPnAaEkeJwu8KH+edlogQbh72ZMTrls
QJfVOQO8fo0ShgOnEBl0nt82wnuUSOCSc3SEdmEWX0MOQ6+9z2GT/+KocZkwJ/iN6YXV3WRfC8KL
bPS1fjT1I+mcJmm/r61Ez6D9Y34K46PKWKXv7dqrMMJNiLQCvpoT4AItI5KBibm3oSx359lk12Vj
9/gIFxODIHG++kO40k2af6TC2ayyz5SiaoYxzut2S3qv5xiaHoS2x6NVBl2uS411bfnNoZcb9gH8
slhM0vjdjp/k5IJFSJYaA8dt/slQw/CdBEcMQeOhipZWRRfHnTYdUqQDGxeTimnR1mmQWdM36+62
+4Hcqq1c1NZEby9uwcZUXwk+ZVCaaDH9epRXBfrD6giZEXEyy3TOkFnXMptZAGAGD2Rq0nhqAeB9
xD5HaXmSCiqmNDhegV1iak8lNDKnVFT2pSD1arfuCWNHZlB70nJ33ZgGqnIRR++vEPHpmUa8n3cT
6VxQ4yOmn0GHhS4i6E7reRRXCA5MNAWgejqmfQJFZ2e3vLkYVXy08hqFYPgmHiM3njIn/Pdxe+Em
BXiBQ4Wgb6dIm9qfiWv3+emEptWtcgH0HJvn61getxpHhyG+gJWqZmX8G2sKsIKR1Id47UhOfWuy
k3py9kEIwtcgJF0wDne+HSgrRxjC0VZcY9+QvhTfDiqindHk0Jw0SyIwQOUZxYe6IpR/MO2o8uSG
TOOHtYSmfisOKpMpteVR9g4q8RqIvmys+W87nQUYjLVu6/D4Ot5t2GUvjwcjK/QWLyF+lxrhi3yp
YUGQ9mBSMc/WbWztPJIvZZtZ3jd3nfebVX1mTdhuxtX+5CeTQcRc0mNwnVCJR5ea/ggYWt3otW8i
R8bX3BRZqJPB4KVVVdhqRu+wXgzWbPTKb3mfiO/VFTqHwXZqD3gmv2q+b3y9sGuHAwmzVh9BiALD
Ym3ZuO7WOlFsxm1EHGPDBP/+rJoYFT5KO4qURevhh4vrRs4Pxa6FaOWoWfBLtOLkBxFtJPhr9U5K
XvFNBhgSrQmEbbGujWZcJadsd7/i9xGRbE0hnPGl4q+XuurxO/IJdornZjaccay0Z6pqmCit2aBn
rOAlcrDKIov3ey9CC1Ws88kZMWxcso2QaT19vvhpIiqSaZ0pGQJFgKFRZmr+ZZkDgzb675Vhf5E5
O0qjgLX064WoBMwGkhYF1V/YW5fyn21VRm0APBA5GR1IGl+k2hDy4IcPP7wBjZGBM3BOv3dZjeHR
WLdYoUdKGsfcXzGUzufbPHEaY6UCqKlTTVkBhiUQNPHASWUjaY1nRr9M/cLcIB5RaiQk0A45cbVI
F+frwWGNP4gstS4lxtyv6NthVJAUugFjRWxqGe7xMgXUilwb2fHaNs+0Wk6Mw1CLCYHv9HlbDi/V
ENDI5eCiCdWzb2yzfE8LS/xbBj5c0E9o+5BAeciRTIQH/UsUFZVazjuAjRo0BjN30OK85juR33r5
J6Iv5bsUvE8kX4am6bijAJfHDi2ZDeQMeMXHf7OvPmS5YWJVjpxJgIFyFx0YcEoDtoyijNqClro4
1tzITP0YA43qdNH/UpnGdMnsX5/jXSeLNCN2/amRJSDpR5gXf+7+ag/Q4hWmsrEkotR37ucwfGGp
bfOYRwErUTktjuBERNV9z39V3XIUiDuNPfZ7QrobPB+KvIplViq8XVQOE/TvnbE7gpaIieme6w9v
LQCjkf6acUzoHR3YXjWNLQZUOJH9HMnmctfqJnw4A8GcBP7WLh+bzr7Sw4ubYaWPWeWwxvzlGphk
vw/Pr7G6zRdZlWkEM6yopeuVnaizbTR4fJBsJSgCxQXbe38Kk3E5ReXCSMXASapHLdSEanD+4wIx
Jpcl6k0nak+ZvRy9uhjSmgH5jFR4VaNIQF9tJl6rBsIcXZM9v4LHH1GO1BZ+n6II3PYbDKPpzzZg
0JoZfG+q531tHk+Wx9q+CHovEEV+mtV3bN2Voze+Al7iqbL2EFbQSnzXh4dqrTTCi8p5p9ZGSS7y
r7tPpt72PJVxKTPjMFYmN+AViV8rJiLvOGavUKN/tleW3zmZrPqXUiq9RQTn0KIInkDOLkvv7AMP
3OqfUQX+da31px7whWi7nnvjQPmI8re3iaECHWvHYLHgV4RophWPwghQkZzEzcaqE6tTyNb99T8h
iTzsJIK89+sKlkJwHWnyKxdbhvqqU4iiJUa4o4BacTvHtRdVQgmV9IhiJ26vC8KwPLUdzRsff41d
yB5PXf84N1DKW9drC+fbEAMAkB9ZlBwI1QrCJAerfqa0v46psICOdsFK6tIQoS77IBEXY56lif8s
Iz0AsifVb+hc24FCrTRcvb8B+J5nvDqabZUp+VC/z0qPUqmC9p8HwTKHqD6Tmp7TpR1Jy7UGRl85
LMlOSVBTu6sYmWYGSPmXoxh65YLQPuh52vJ8WowCu5Zgnwjcp4oUXcfVBqchO8QTxlz4hA2LPhN6
Dt6G+rVM20yOU0UFTYF2AvSKy54tS+cy4UBu8wKuJBss/Nbi0ZWu6mPbBOUVnNIMcHDru1/ob4qc
cmXr5Z8proQTY6gavfiurk6KeEc+gcKC2cPsEwZ5G3TCyW3H0N7bCrSUwA+NwURi8Z295ZKcs5wA
DrpOdqIKlZdj/zjTBYGDZXy1PS47hJGwCpk2qGE/usjOupsZ9qJb5qIU+Q3Y32Llb67nHhSYxV+2
xxvWeeuM6xjmH8PrQFOIBgXb4lyKaYuhA/V23tmBuSx3o1u19BxDnKJTv01tVhEz5mHi6gpsh8St
VqneDtcMX8LvTdXJLdcn2P+7s1sQqPZbMLINvDZJcaHKtzEupOK59B7y1wLLzJUzvfN1EO7Fk7iJ
e4Twy2MOZmxJWbcTT3fAtlEfU2ZP46OHPTSgvodNqDxxFTXwLn5KHuw1yEYDlwTa9FdwByACZ7Or
7TdRIsXj98xglbS4/x4gY5uiv2xBbdP3Edpukv+r/L/kE5CfbD94MvpvxMrVsEOaCsrYbn9TNR2o
zY95w/HQl+lX4K/aBrxT3VTHlF0kH2k1MK5Zvr5ixF/mfQmGuzyTbqN/N7TZgMTHLJBsrYMFz+SV
qV+GmUrqFL5vdEG+vS3fMvMSdZJrIQINmxrx732Z7x3EbXFlzkuUviU7AjnRQDy5rCgeIJxEXRMU
pRZsnteo27ITWO5aA6b1KNG7umFs5nOP2/n8bcKJEjuALpo7W5QY3AyWh8PExjF33jXOolctDgVN
J47rQYZ2NWyTCwwt5Hj98bZgzmpS3xi+rsBeYIPZ3UO9PgNQpdTRWtfT5fIYKrPqwH0VNLXdcpwZ
pjxFRFKZSjX78roajxZ5r1c9dnQGaBJoniYutPZAJiwbaxMOFbo4frPijKsDhlWc/i26/qJMYkaL
GlzFcFdIyVcO5x9FI7mxskiT3KIzznPoePcsLSht69JniCocPRXTo8OztGe5FXtrHvgMNcq5sCjP
22PmTmeNI08I9WTWDSJA+bGkHXoIibPd0M+MEkWd2H0km+bO8VyNFUK3YItZrCzBxvzrIQnCzy5P
Pl/Wt14I+iD92jVjC6XgeFs3Pa28LDzLFc3oMvNZIEbdIYLlIUiLovjukt6acxJjuao86PN9UUa1
TCOHgoEhegHcYdTpuhKVzlbzHGcWjD1Y1Wmx3tqhQtfGgQ7xDCXJ6DFOdN4kFmdDqwHQ0qzUpKy+
RWoiaQPb+9NimdKTAO8qOL43vowzl4gQPU/7PKZZZ6u06VhQAmKs6XomWVD+zUA6dS95qTAkmbAL
Zn2DbZ1vg/yTd8SyW/EyYrXnDl0No6vLj2GPnFRkHUuLq7FXVFOpiplESMHryTaZiY1lQ8IGar0G
PwC4BfkUZsb57+jV/JqZ30xKAbOF53uQDKEc31R28I6goEGfNPbRK1Lmyt1ObxUsO4um5oChz7k0
0e1gFhOzPr2dLwI6HvuIDRFOBIVv6eX8ZDipfzLyWCQdavtfNcWUabhT3fSi3iKsF5sN9qV8J/po
ldTTnzqjOMoTy7s4Iy0+rL0+JYWJF/VIb4wfPrEXFIViuM8zjvzLDfVwhH5J0V4p4KjLY3UkoxBo
XPmwWwBegNFxX7uBKfQ+y09oJxkF2xmjCloOYNtOJ6jtkfELr+9Jw0hsAPvUVzjdVSjpiKgT6uyj
nypCe+6Y7cCH30DuQ5wVkad5E3Prj0GuKccSnAcHZqUBCP8ug8hO/DtSPS37ra11AMn5vI/y2XOR
+LfAQqUF/JgQ+xn7im0piWzceZ66v12ZcHHglhwjyLjr+Joeljea22wIFxqKZNh15OhnzeSOWunu
/26YzlS+KkUalx3377t4XYiMnsD40diX68Hr0dYc5uE8GeOrb4pRPWcrGHc9kUNQwBzeZvbTAGFm
jLElMrEYv9RDL8vqOXL35a4m2hX8hdkqkWG5yIo/hwcxgjKq9z7KjG7g8wXRYKgC/fbTWZ2Xkj5f
HABy5SfzxhkiKu71+EufoPfnzmg9swXhiK2/7hQ5DtvWtvVtOebxk2O6PlA2JDXrkErpBI5spNKc
eNx39RaW5A1ULkd4vQX6u3kxE1SV+hIp1IdGNSMCMxDZhsQtXxFQ4yPoL6mLQAM2b1qUFYchYJOh
NF/RTUmzWOmXnbBq1XheBLPO9AEi7/IH2No/pSsA0QtEsprtjHeyEombqRx0jcE+FHEEkT/W9pki
T+ZWG/NNZO/xIfDIbujoP1dwoxB2jzDzCfz1hhY/uFQ+lvYyeTSkbPwLUHWAleLsWeiauIbchOu1
q08yNol2KcWcVqGDTwYSErkYZJ6mX7Ud27lSDYrcBhLB0abYMQbUfbLjJr1k1C23m9+mOunilsuT
+XdMHm4AuG26dpkQDC0UsuEy8I3+QDxlTPQEz5utxvXZEe4ITUAFTE2ASCArtfGp34gF26gEgHl2
LPu53rv4lbIoGH2MY1SivfWp7lCYxAercKC5Fst6ikr5ZKZb9GfOtqtovEDTJfkk+wthlk4DgXn+
IXNcxt4UnuzTjouicxsZeku8rCe+sCR4chGbkOWihMXboqSqzvWkqCpr8QsMauxJ4zi8yeSo6sKK
wgdLg/Nze8qmu0ZUHGhxQy/BH8vtf3W+lOkXCYvOLVXPF7uHTxdXMsU3FpeJAw904dk1rrySaC4X
uwJgtkHkFVSKmNiG1V3LkRQ8X+JyhDwrroRYIZW+B8oz9cn/v92aXWvuWfHl+N2bzY1HxHImTzLX
cPsdjR0+EI0LPmiXDH4aZMnrTj0RzlSMgrc1EOCFgsxnMC1LSkY1rOtDBYYFXZZsincBTQCnQbmK
8bmtj52agoQGzP/j3TJVIUHefVw3W57ZV2HDUGNtN3sf7VnZpbxUK56q7iF9/Q15NMa4n05Cve0Q
tePVeBGyR6KuWFhkH3cxQ12njkmIr7/0ggS4v7zQLvS4gu74340PI+M0wm/mjE4iKPEEaiPAId1P
EHB8MRuVaAEQaepogB82diF5bEkMARHhBSeKAL/lt+k7yyHIyUZAPzohdmfngevVjQjGZ8rXanQp
OaetXHRTU8INIG5fxCy5o5NKJNsZXHAS76yrO98bU1j+poS6iJT2YfLebrcK2AdK+9F56y8ZiLmv
I2ThlFRrURQ7Gc5jsBQqSKe2gmqglMtgn2KFXTeCNxaPgTR7gWsDRkxz6d2Iz3G+TS+RfZTuvE70
a4TBTwMcH/OrNTAMdA5aXjOXdLkUnLh58GY++QmrEOvkmctIchgJ3JrIsy4Cl8djEVqtND7eBDR+
DbiwoJYt3pSzV5FGFR/Tbr0L6b24lQ7bTYffADRlfWjL5iFUXcNyKR7jJAaYJWHBHDin2qnCi98Q
3MKPzGMitrL17WUjegLW7IkeGfPQq+mqMxatg2gCEy/QAA4CwnUEqED8FM/k44fzM3CbG4sO71wZ
wv93VYJ7o0yMRTuTIjT1GSCuV43IG/v7ZdzlxuQWI0UpcfSX6xA3OWQcWuTvVCQe42hhdC1jWbB0
6mpxO1+uQgyiJjL5HKH6tfKhyh7nVlb9VbrfGZhTh1p540I82WgCxqkGR8mrt9aFJAh3Jl3t3YkJ
nguHz2i0+PhXzsAfF4tvjlsZSffLzwESVEsQS+GMnkOmz8D8f9+Ty4HeXOGHeYX4EFKYOTTGePok
PNuSRlXVSNMLzRPtagu7m5pzriHlkWwqxBNzlxm0ONQqPL8PgoDgwqE/nkQcvcKIDAvfA/2ZYCLm
ufbA4mPqkgMgkukgIX+MOICm4ggZGrEtDVvLI0i+c6rULI08ZDeWUZOOs0nRWMeCjPg7hEpWfpsy
n+GgvmbZwrfqS2T0enG9ppsQgBTyh92e31kRJmRTQzDT6BgJmLBLcOn6P0DlbffF/eTQERBRG5qb
VeBgMCf8IyaegUXAO9mW/juuFFN3ZzR5ZYMA/UWqTWAWi8HHDoQCRBG99E3KzBaO+AoAq4hPzYnK
+cb8y1IwYNqDQyhMCFh0EetqQXp4DJRzPrQVA4RWd/+/G1lcIdioHs56aj8uEgqLd5S3WSVHBZDz
3GQZMKAXKlA+8opuFnUU6wGlREBJc52Q1hHgnUmvJ7pdKmu+fpyBEFgSN4MmgsbzDhb4Ynb0L70X
d5+2U1tEbEoxwAZAB5wDs11ui1Oz/ZG/Vjd+oJzcpHBU49LWYlQaFisosNmG+NAma3r8OunXGhU+
NwHKOh0ANfa4df//6+uFYN4eLaL1kFhXkfRiBsKEOywwZOUa4txGIESTMNClqevYe6WhCpEcTQaX
aJ3qSok05kkQ7UacQiwGqUUzCOpWVJK5OuTxJWr6+ufULSLN/8Ytl+QKRj1MEvPxDlPTSz25CF5a
OzypG+plaAG0OWyj9hZoww/cOQXLvFQMcicl+NujD9V5W+0jPP0KQhG0o4k1IcEUFYQ2JTWMgqVA
ysfx8tpOSoo02Q8axKplR/fpQPznej5TPQ7UzQqdIbEVuHXFBn6cLJjh7LXdPH9yrMd67RHhx4FH
vsNjpsHgmI8r007JBuojMCdpW3YNmO4HMkQnvxZR/hbWvPtuHhdandvsHXsNB+OOX/BXmBhJw8jH
fN0JRyldnaIzKU1HEQTBuBVj7vjdhEAkxV1WoUb31vptyN0OxGigv610Mb8J/oHFF9mQlcQsh+/p
AJMmC2lJDi20NpXs7qdUgZUdTlHfUnmS8UB5h3j9LxDJr9EdeDSXc9DyxC0R+gcFIoX0rUlhTM9Q
VdUUbsEs1IywESY72k08Qfh1IvlkFiWkbE0iyiOy9mTIY3d+fuvWTnKPTeY7n4rooqgg8qjfJ4RP
nx6yQUZFIiLA7ibkmQDfcWSDfWEmP8WWTBzPQOAi4UquMeqcgppUA1zXi7TezRxK3v4VuQqnk7BN
SOmb46DGD7DvJ2Gvy8w9+H9dNwCvwOnmSRog9heFKaOB/6RZuGkAMVKFH6ptfVNAVy2SKuDDeaWc
0rSga+TWU4rm4RG4R/zPabIEHtRqiATwVDt+a7GK6xCFEQlosH3RnxnT43nALSWGMcm8GPpF3bZy
/fZbuTKFWhxosLjakrKaOYjuGVcgyAa1enGM6PegBBYwAXWFbGnxf1mSTit7HXwnR4GgFMWrjqmJ
gNDNvVCf56AyPQq7kmGGi7M6kxNzqITIpNH6H8guIa1x4GsC8+dvi3AKRffOi/ndPtcLhgy9p2Qz
CDse3tTD4GxCf8S/v4YnCoKYk0xe3saceJUtv2xd2yH7l0XYfRsk/Q8l0Z4x0cNz0/1Tve0Nwo90
RnPc7ZdMQKb9hsTYop6JdMFEh6GfXhOnWjXwV7VuY3kuVqrwFxkYsy5HWpcAU41f1tkNMAe0zhnJ
zC/dtB8DT6uHTjO/goOWziO3sv0k7H1iCtRS6XLxh73eYOted6wSiajvwe6DY2xSW/cQNfqBljDa
AxMD/cjcut9DM9bJIIGpIf2otc417Rc1iDerKj5vqPvb+DUT64M0XF+msz54owc5iQ2ohWhg8EoK
vm6UjZCVnvj4gSy112VkV2JLvbPqoVhgnKAJKRMIZoea0lUjoBf2xWvjANBbOUxiQcElmPYuwM7X
wove8WTIRGuhgJRkG/jCV+Z2fYhlfvWjZVUQZvwJV/NoKNg78UCit0i+e9uIXiOGPMWE+kiSUxBZ
iyceVrYcSKnygfkiuYGWTJdFfowIn9GIWC2lDriRJl3jwoMS8P0YyjLH5a+ymBpOtYBuJvnlEKdD
qPM1cbA9KyvPRWt4X8i5fLC6F0Kf4d7o5MydgpxZWAGVN153aXvsKfXSEIfsdOkx1p90xhr0oq0u
ReWKZfC9caWvL0a3eLo4CigijglaDY+2mLHbJYOsBrrNoHTt+mKYaAiqasRQyUv/w906WCPhxT9d
oJfOzWzGhWUsmslIgjIA4xr4Ot5R5i/JP7NrBEW1N8RR8KzdYnb3SzYeHz594VMaKa0hxV7XXwVZ
Tx7RdTa+IWLBvuU8oU/9A5FRZUMSStRfxqtw8YITbjDHS+wFnoadCqPzY4EhUsUWT180eorfsUzZ
Umnpmwt8VRdpPTyOw5Sij4yZL6+AmV+iZ8zjc7XTEpYIxXPtiWUCql07uVTATcuO40tqc/OwZbFB
+0FAx997IzHhpGRFnJCUeFz4yCfcWzlALOWenyDRmmzoifwUHdoWrdfwk7f3bquyA0+q0KPrxEk5
XoU4NhzB2cr3KcK/7/vdfl68lvIPjIE8Z59OMimIrkurJjlYeNrXZTc1nbni7tCqkrJFggSot7KS
4Ei27PI/JbqwWjbnGNn0hyFwVBLPjfEE8NZK9BlwF9JAlCUNAe3AoEMP7Cv46/sMpWPvaRrp01bW
EE1Bi73ysEORBkSgMD9a1x4xdy/FESkw5ZZe07UPakCoY7uhPAYoAaeMlfdutfYXSsDCDi99zk/w
oy6Ax3kosC8D4E74OS/Du4KZmWNCy3HaY8sH8xUYXwbrNCcSBXq1hZ155YkbeZnx5ZzvksCGqKp4
60QDWFXquysZ7mxxYx/Mp14N/FB51ymToUHZUHcQ1OkivbJy6OpPiVCdYksGYBCJEBFX8mmp2orl
8SUrAzE8VYXOng2PkwMuaKw8BKTrSbctmNIJ/swgkp00E17qtWXsgt99GFJ9f71wpS8Bm1PiwZMU
FOYRA9rW5DQu31Qe3ZB7DrsIMeiwgsVLkTDYaqLO04iVMzE5CjmU+7pws8px6mUZJbu6CyxWL8Vz
SFs4KcHGPXcGAGYg44DSY4crtzUsdaLiIsmVoWW1329Lkp96yMWYnweoI7NIcXmhN3xxFTi6LMmc
tKILG3I4F9a21/XrxVI/CzHf4KQbBlNgHLChiajRtie4Ar4DAyywC8VHdHb/Ftv/B6CXcLI8dgS4
MRaTXohAGRcvk93ckBxHS0BPMbXlh02mYQmtPB2cXIclhMANyuA75rMDTuXFkBdbbOLcXeiLzE8R
08HcoZBvS90tZ3jsvwLMKNZgBL9y9au8nHsOAzmpg3c6FR/obbbEPPHuVA44rYLeGI3ZxM3Jkwvk
p6jucDklyFLKZHI17bS1hQ8BUYYFfYj2J/6WuT2zyFltdhuwofWFgloExJf8MaV67kOs6I3BSwkM
7AKbK1Ealz82XhmiZqyVUfqDCtqRw/FZVsJHwbx/aHx9SHU0ebvY2WIpSqSPV8F/ZLHUxT3YHDrd
UUAuLnGiTlULQK362Kfx+j6kn6GudRjvnHOWN0+ni+P9YkvcjRJh0xXT8vESmPorxlJUPAM4VRbg
q/nowwoye1wkeuBgpLZp+S+U/MbQi+1m6cHqrKJjHu8xXl4tI9kX4BY1tVpvre1ouWyFdwDDQSM/
/oSP9iiwKlUEY7aPODEdJidPC/xskonB+gBOfD0NLEn9PMpU2tUw5l7DeRQom3PQ4ggjwbMmwjw6
ByZt6Lp5KeUJtAKpZSTtoNEO3KIfWjmZQNJOZ5rql4Sbp7gP44YDlZFQxsXrJLDy7ZP91lKhuXcu
Tzp0xgKzo7R27YOKQ4vln8o6Mnf9qeopMF7pNxXF/xiOfq0VaasBZpPjixbrwDIenmc4exe4Fhfc
F+iFsoemeq/JZGK89oSOU3VectheXex6wxxDIDY1k/SWPwKGbJwn1JhFD7xZdVc/070u6I1C3RZ9
KQ8UBz36Cngtasgcalg989dtgutZ3Cl5XCaEs5BKOaznYj8M6ul7LM1LDpIs5XJN6MVNhDZ/sHqn
2GmTErRtY+lOotPGA8JQ78HGAnI881+y/ZVyimfpX1gnlNNXgVql0CtCbjHeHddzOZEda506DXP1
auHyptyvOn/cDI1GO+ij2n8bfbVRCPMqndZWcJpokh+v0XadhqaeBajK9pWk3nXOc74lUchSVxQl
b0X9EE7aOpd/2QYwaNUh+BLO626E7hNVhKXR1SgrWCa4V3zcm3/1APFYifiFv1k4nak1WbCO9OSr
M1jkB+idsby95mZWhrvbgu1kWY7QqnjmJOsifwR3RfC1YOwttryL8iAz2QgmyQHcUc0rKubg0Bx+
Rrelzc6v5VWFh49/xv3zbdyb123wCfpODBv92hCLAw344jVmMPydapFnI793BL07pKd/886PsKeH
1AcLI2xC1Rcz8g608HPr6aTKUO6/TGTrhH5wjIoc+wYeVaE0E4DMay8ZOTne5JABbBg2hyoITyIb
AwCOemVp5ccq8P0fftlU6PRlBNjlu75L9Mkq/cAln4INJwsaGXXxRcqvFMn7jDPln1iCXPbiwHPB
vPm24Szwb8UWYue0RAxih+FIR8HcIigr6T3NaNPJL/cD8/4mFKhL+Ytda5UnRepGw4ZJSupFy4C+
Hd9BEtSqIHrniHvlOaSV5xT89S2d2IrepeZM8EIGxC+aNNzL06BZ6B1IX5zYswkpP+kRjP2VYlek
j8YbSQV4y9kqVj27AzfCTL0HQSkeITxtUOo/XZQvGcqMBx7Nf3+Fd/tuinaRJMkRyW18z9IXtx0F
69BPzTzuY8ZMkJ3QI+prryElLro8yGKaWPGwZ8yDUjzJ4sZDvcbWqmZQC07/AwL/LLFNxPmJKpeb
a7PjW8qZwMLytRMJ9rSYJh/+HtgKsqWBErEtQmvm7uCzT+GLxhx4Xk4wv9yISVidiqi6N1ANt79c
oyVp7Al5QVzRZXQPpojB3KbLckG/YAIjW4tZhUxblqET5e45gEs+hTQFQzjGypOwhY32kMWvpLX5
dprzNyiIKc/XSWuhcWGRXOblukYB2sudNxumy6GO+CyyWhtcHC+u8jDlljzklt3hZsfd7FG0UwCU
Z5DBe5Z65GQKkdmR9lvL9C2pDvhwUFR0AiKYzvTpS+ktHDQzLari4YU9IF9TiPq32xpcfpWMhk4f
BsaVWLKJuYvAbG7SwHeMERjUygfU7fkxm7RiU2MQ0kO42AgdSWmOUyesBAiBGcL6dnWYLOPeV3F3
CNlAoPh15mrlDHBmvi3PeuZyrkHBBvHQgtkB8vfSayXLCcKPN4a3NHPcykJwbirXudP9gNDOqfUG
k0rPoWlgvCxBAygaAGK931WuxZUBMHTmTb0ixc3N1Flgt7eo8urhZK+oh/2TE5b3ZqZahYkE/mEu
bRTnSUzxZ2NsT8ByMS2JwfjFhVEVquoO1zgbqVH6imUQWIZV5Bq18DCne+ydN6ttoTCVkAPXOGpT
WJz15LCchkbvkdr2JHFZNar1oxpih7F0z4PaK69LbB4ZYlrAuXUmmRIbeZpQlcOxjVya4Iyda+7i
YAxw17mQaJ6W8C9+M2NbjvP0fB9dkh6LbLTS5y8Rf4XIhqRLvXTQpLMdaVhnffPAIQfculjEcD5A
fcSUR5MsozMuHUeqVb7SRY64kzzgtGLqbbdm8ZEc0Im1dT8jC/3SmCyRP50Aq/sziBvCZ03AE2ij
WWGCC6T/IiTZRw2yw7kC6NTvCDycR9LW5OI6i/dMnrak7GijEQrlpTElaOlwl/bZgrFPqGpG/6Mm
CHxAl/Kji/+kHfSddEBFXXyhlV46inBucYlTIQSCuB6BtO8UyAcopwUgtZgXSD4y0VGjiTzxUB1/
UfgiNck5eUJAxoMWvM7NumMVQACk5897q1ujPXk5qcoBhlFzSd25S3tZ9vCUR2HopdJHkDHGK9q+
YIRlQpBbYKP+dj+bw59bsUHkJd/zo8vfpunHWdirHmCspQvMOvJTUyCRPczVkQJ4YleMdTLL46wh
I8cISwCUfhn3j55QD3tMM4c9EhdeZOsCHiKYQNPvfFXy44utmMJUEBlAOPLKWsVMVQGgc58SVxcG
xJyOiUwHOI0GlJ4JjCaEOjIW65SXh1mYHX+wUv4DwRs60wlXCu3hgUDnhXHcpUPnXH0GOdyvPbPW
dBBEYcJ39i4Wy7TvOW8CHppRrrs7OGxPnSI5TpSllzzH1SVkYXB7kWdSSbsfStlzL3lxLqhA/z0t
JrybfK2xEtt6SboOHsC0JSOVm22JE3IlgiZqLH7QXns6a4pQepPnx2+R+WgUVniXM2cWwHa0n/t6
nMI7ACGeANPwW7Kmz3zTS4/bX0tmifmkiq8Cu7gjqg7FUGQJ1w5I2eEpOvNi9CaiCl4soueTA4Th
5QeASoSZ5xabG3I5uCPLidPSvZ/xIX3BjJdtvhozlTOjn5W36+v/vo8hyleJDHJq0pYtS23hqLoW
4/iSlbGr3jwP/IZDUzZ5tyt6XRys3EkSNgf9mPx2bTYdxPl6T8DT5ye8+5kLUHgmzdd3gi36Or1m
lAv+cfiPgAmAH27SrTmpiVEayErQ77Zwsc0KxxmPinU0AfVfWyd0tACPKMauXBwwY37LCKj1lcZB
RqHNnI8HXyeiwF19Vh5tLJAnaF7F/El8vgxrXC8kueOLRHwj73TFw716KZ9gnDI7OzQXWv+dQ/tm
VOsSnB0dFTkkOpEwaC+02SHqTpmZoFNxD5gJKmNpY/5L2B4EmAyLZUvzyqZkhICJB48/TcSQggO/
JCI8r0fs29g3BLE9HCgPQeH7QQ8hoxKLmxiFoc5RK/1wwVlAV5m5en6HJYlmaDgmPv3dTx3sn8js
wil9tMj/753hhalnSG6yHTzoupRfFF/w3/iGCyHntllFUFb6BKOgPtzDvglKYseBvq14OANmbFg8
VSpwvjEpUfLuX2yJY3REZvTmt+kd43MzA+9GVDM00MbwDRatPvhkqG9pwjeSjIQgBfUC38giPpbF
aUObFsPTO74Q1gCvCAv14p4EAGPihWXaKiWCwS6y9m3I0DbYTujD9eoMwdD9QhKMxyOZ/cOOPeN1
cBAvWOjJGQqvIIVPEqdANoi6w++6guslGIJFxBaiFUutjXHtgCWBQoFu3shpkbEk86LXiNSKLL9g
65bU8TIwmnnTKZY9x2uZNoGdc6rPoVEDw9VA1SFLv+UumIMECSRi0CbD0zmDlfTwPMz6fwaAFRcJ
hnZ986eQKIBPRmal7q4T68uJpW7rCRrrGjwkGJrdU97AN8O+oJI8BruRoPrXLQT+VV8uFS2X8v+i
yhHGzN8qmLC7eLIOhF0BOunjmJlj2j2veTbI3ZEmJhkE8iy6XHVtWIFPo8Xydlw2SCBI6nhRRsq1
FbLlXnpWkfiA65l/kCOZsGPj5n4w5b55c7+U2ocr5gKg9+Iq0qO4z2uK70dJKCnXceVvX5rHJRwK
Cjjn+bW/aXq86n2suaNJR3owN3V4kzbvGipVkSF9nvFOdYfE9fzREBo72UlIZq9fSYM8ggx4Eaku
IhUiKOs23KiePM+8ZDXSGyTTLeIIPz6AXaGXziI/DBHDRmKVjEwXkAxY+dp3pF9xPWR+QOax+n+z
L6rKx9Rdzo4Z25H9As3eTqier8ssbNMqVW6QlCPphSaCU7cjbdxGkOSyo2KQxM9cZKqhkCh6VVAk
fR8TXZF9+cdENaWQ01blZR+MWYsicH4F8fNtnlgb1SN9xgGcanQ1paLHPg3zl8qC14aWRbPgfYDb
g6AmhIUa04uw0nN7nn4J6CXxHqj6D2pOnB+TBQQeP0o6RkxpUIpxU1sLw8Yp5I5kdy3tozZB97iF
Dd3YwZeQh6idyw5PkGbkD5RDJcqrQLwymxIxIMwXj0uZ6/Z8d+ygenDVUsuPqpb6L9CBw81lrYYu
J9wMbpnRLoDZN7dVyexIRglAeFoUU9Fjen4cx0UZ6b75X3RU9qBf3G2FoC1BiVB4PmJ6xF2MRqX1
iBL7fC5oX9nb16oWzE5SvlSEJ6v/FSTPjwDHL+4govdyYlIOMfI/esGueZkhxICHTt+mrlOIC1+K
UM1UQls366Gp/55aEjC7BJw41hXbPFK2LNZsj4oZ+zJOhl8vAyBa5xVZzIn/aXDES+6drB5Cdmj7
94gGYmC4w6V+cu8nN0x6JcDGFzNmwlMLZND1ghAf9ztDQCBg+OeNB7yvHnPVYed+9eV+Q7tLSrMV
b8I3OH0M6WTCAvGEhxklo32XUT3GQ6A3Trkvg8wIIckAdNelFStMJ2aaawu7+LfGWXtKeEMFLixi
yDXiQ0XfR3mjVzOTlc5wHcn1mwzETsYzCe746qUoPlwTMO8IUR9g/T2E0wOddSE7N+B3l4ryt1sG
ba6iauFZAzvAEjSfCbWV1PxH0u0MrScvfbygWAXzwRRxT74LoH6UBx+o4t+oqpn/jEA/zsfybJq5
eE7YFv2DhjOKbvcCZaeeQXwRNDNnuyzPHQh/045hnFEzMOEONVHJth/phvOKsvsdEXmaZmZWgkiV
YCdEON3EaSQSXh+/TWsa0Kc41qk+WZtD2VBn6UvOAPO/Q8Y+HAvKYj/H172nMqbJ6KNPorXR805x
m+ybCeMAW6NKCTWcLsHQr3W7JePTxbrK0TGEnPK3WnsqcyvI/TXVHqIw4GXz0galFkRB9OKPsOwL
VynhocTkRRhLzME6gDzkDnXrJQ6JaY6Estgj3sDaaI7xvswr/OYBPsM746kkWJGbw3dHz/1XpPR7
FdLgTSx8/OnejT8Dbr1a7T4/Tgz0r5ekoMH6nKeTq+0v6vJ3bR5KH6AuY8jHL1EZW8qvjLcwtXbf
uTdQDLIyLhJkPSGkr0PQhMXsOV4ZuqTweNkhooWZVUvpbNOfET0I6gFJgyZGQ6IKo3l85FhOOQrE
r0NZqw9akZeEhU+gRLsoXq0bY00jMh7wLAlVba7qRZNXzennksfKejqY7wSlQQApV+Il5csD8doI
gSX6qHxYFvXGZ384dyZV4M7igAfr3qvkhsnuDxOtiJNG1AsLZ/PO6WNPjB8RYs5XTFzxU1gsgBJi
gQz1YOnj4p/LR2opPfENTf6yeTfrGAh9b8SQzHLUjWzSs7W/8HzKPfEq8yS+gbH2bRn/py1S0pja
wT8KBlM2TV2R3E5YP1ataQWeDNNuHweNCI/m14bzM26Sg24sanI6Hmr8d5AGRc4f/C+mo4Cbf3qW
6qThxB0IwL6GoyORZoEfzihyLnL7lJ6q4U4OuXk2/yJ8WJVljoBxzo0kDZqqVJZ9MuX/oQLv9S3y
ltA86MIWD2V9Qv5NAuLcRXtfwrxElixMh2sYLXwgqe2KhrYGVblCYNGdjd6hePzAlNhwDaJmirpt
p2uRytD3uRADy6Cji9eultvKLaz0mMBBBUokI00qMNU9OM/velEWBHxFlfgAWYRxBNFBNDi0UXNQ
LAUmq36haNjodx9Ii9RoAyTkVd8v1UyAzqBtB8rTc3BrmNeCTQLuY6zAdTO9klfMOUaPncvzGgey
1KwO05veuOAepBG2/YePU3lgYzRjvbCPzf/KHDdFUbR/ETRtC++Z3kQ/gegDE1fbEA1b7GO0x9oo
MYbGsYByyvvzMURdxndLlLH++XuGuJZlzC/dK1O8hJbQ/yJ9jjhZYvYU4FdxHYsryeo744cMCn13
V+k+wN0as8pO6xEJbmbRWIXgEMOO+tN5O3E+LBt77eFgljvWUzeLCZiFHF8u3CunYuXnPwXzlkJe
EKj1X/1fsJ/gsfXTDbgnZSH8Eiy++B3mLWSIfskULDLSYKurraZCmra8VDNNtR9L99xpega5H+gA
Q5kP2oq3a1SL10aVEL7xKPcen6KTu0l/guTY1wBMzIoQOD4ngAvmysepb4Thaw0GQBRhJWYMs9rt
Bs/SnYb6qQ4ir8ov7DKC/5syuEgJokGzbVgJUjRqItrlqhzZuc+NfYyl/wYl8crAhs2LAHakT4hy
M3dEGELj0sl51gDYRp2PEjV6W84UGGD/Ux53NolC7o8ndgQLp0g/POFPAwbG8ZlHHzGMBa0wuke8
gtfiLB72KxHxldEJKm8Es/FoN2CWh9fBMCbmna4BAlTyAWxKQzVsAKdTL8vMsh3Iw10QzN6aBvWS
3Uhef3XBYwDMA1rQXHlgMO1YK+QDiADYAqDPp03cryaH3HW9nso3QfExAXXMvW0ArpdeFJ6qkEr8
0rl6XErKibEWhLG+H8Wx4zHhNq3238MkjOmWjqUkMhekAUyBd1BSePSUqZIOVuvXRM1sdnZHOxA8
LZNtLz6Tu6rJu6XFhNCaclHfd1UMG9p1qrUmF4V1KcOCzMCETEJDvkLTtDdSJFQktQm0Qi9IBYqG
bakDbozGije6ahRLryQPzn5SPqLW7s/xUJzjfT79dHNN0mF6dSZT+MlRHRdYJkc/9wahic00SZDt
+DDHHGEVlGInStGefe70cvUarNN11cUN4c2hRjJZjGNB2tw2AGOPfBcAe4Fb6KBNnoTxpj6TJpwt
5Qn4lOxxpcsPqRBDf6vfHfqmBAGv8N6qwbkzJJS5dzPGLIadj2143YT7NWnHn5QUIFlkG4sd6HHS
7j+kqBdDegATQG857PphC0S4jzE0GnxAhu74TDnSG+IWq9P6jhFB0mmh8HhAfjaYTDD+3M6f/82M
YiYckNw6/2cv66Mm3xodD40XaUuPh+JX84/ZJIAv6YmvT4Q2bKThch7v5Nw6A31CvHD0ZTcdHbMk
eaT+RkFF+89Bnf0HoCZxl5Na5EATZfTFUIdmh/Tnr7xBg++QrQojT3KJoC4p5lGNicY7IBV+grUH
4hT8DJpxF8JByKpNvzoFvp9vLtAuCnszynhCtowItXPfU8q7QwhpkR+ZizCpS80RSG/psLiDmTpT
hy7m2XzPO78pMZFJC+VXs9a5K+ju3DzIEOUeOPjA05Xd8tUYfMgmFScOXYvcu8jPZCNhs695exLS
8wd4hlJt1MU8vYf3gWWf118tYb0B1VWYxqF2yYvCNSRX0j/dpPbwBlpeftbSjHY1zESKlXOGZBSF
Gm0FdsSQQtsgQgMkc1X/YtJKPNSyTZP9KaDyFNgMHGpG+TII5/ncW8+T1/JLl/4XT31SQvEntiSm
7aKOjOrQJvDnkVEiCjoH+e/CdOvUINIylcrWxRkmLMDjetOQ0d6FI42+e6SOjwyBJYSOx09XXRFL
M0NhAe7PDHDW5bsEARkiH8lNXQet9Jd27A3L4NHSRqwfHdpAbJxmgyD3+hN/g+bPHpb5ySrvIH7O
92fUmiF39Q+9rx5CMX8orBym39KX2xCfOFku47em2AsUEZnQe9B4mEG0m/lMDMVWpvhvwnbxSWQp
cyN/toBkclAJDZ4QDETK+j9k3g5XKlshSO7KUbqPgl/OaR7jAadDT4JX/b9d3/r3+p84FkmIWtPq
0MWfT+3wyjNzMFpd90L4OAP4T1BfdKi119P+LY4+p95ldIxlUTl3CCQg7WtN68zOyA3Dl39TEnY2
cqRi5YnSWxltM/Kgh1geiNoxM4lS0EV1tMoU155iYYlFiYCUw9tfILq1ur8QOZtYgHUGGjXSwwSk
pXdZacZX4Rgg+Um1rIprGQdjdeyqdIuQVVI2z389F43w8FCnah85uXH4bXj3MZrOOTAwVKYFv2ut
Nsq6RW3hC2DzXSER8DMn+d89Vn95d3ReyLfPnZ6vrtUXhNe6JeoeJJTr5CYyxcY6wD4+4v+KOsxB
9b+OLv6WJSaUQkEe9m2HMIE3vXworPXzQmF/pDh/PaD3dNln6DaD3q4xKkOZ24LA8R25BouKvSOG
BNXD9SRjxbQsYqfRJnIb6hpHiAMEPtlm/VKTMU4vnzeTAWW50J0oHz4RdJ59OuWWxDyWRMS/OMZR
dyftt40Pib+A4x2LYpeGBAlVaZPDorqq0VNUcVTBsN56IrOIycXyWsjfa0yQvdijkSYCDk5eMayD
u8X/n6xjGvKQTCyPPztU4kyclD6iKGHlbSdHsiitcGtD8VMd1u29LikvY6NXCshhOUxCY95UZ5yd
ptPUdAbTAFaKk734RXygt1m7CW//pbRufbUxpEeuNwL6gWvAAhdrd16abtT3oJH3XNw6bOfWFNYp
qjDV7mazEblH8L9sgndA4orGCJXyrnqw4+A5enf9ez/pct8t+4zbsCTh9pBQ8dGGct4zmvLRZkpi
T1fgxQ9vUiwAAajQukynN+FaVxbYM7qyxjO1C7DchGtVvPHVYyZOdjbWOeHJ87iHM1A5GxYPGvdv
l6QnVMeKZbjbcyzyQGpt92anUjeC8jNdmrEDDAhzRA4oDRD5HGNvtiJCIorhmIsgV3c3EZPov3LN
gEXNrJQG1olKyqEI3Q3WRCeyCqa3bUZyakwgLCkQZ1hmRoDNSdnD2NcuKrSBF7bod54v1fhwRGag
TXn94To5NmdlZCcJS1L4qgWHTpO7UFSCyEXxdN8ot/9asD3U2WiPuvnnkO/T9KSC0d8G+aOf4b16
fWK6JNQ5NXXzK/58P7MhmAVeY7HHmjwChBJrj+NTvQlYKWG7LqjCimAzeX6LLfdizwn/33ghNcUu
IWW2khuRMaHHWEYC8+7JS0/W96tkUmLuiPowNq8f48rrUa/LdsnNNEl5Df8tmAbt0z7j4En9yHka
tjyZ460I2Sue36r0zcBSEMlLQEKCTccOUn4LKvvrL7oRCZPeSSD0YRztumkiR3wNaN8Fy8ptai18
7Xbd29ScabyDW1xrOK+wsIVWhP7RtlShrfItp4ZveR1A9rWbLKu9DkaYrv55YiuQzDWdNN631AoF
PSiKSUPIoIRA1Wc7ZgJxIXZnZS+ULOmluhQlJHFJaDOZ0/GX1R005Nzz4HJEet6n8KPEKQMaZd+z
tNXK/LB3jT4cmBOsXxGNjsv9rISWGAZf9mffk9lt1bBZhSMXve8X88/dpS3u7znv3nWsC02vMFY9
eJRrT2NoUgkcyuWYKIOxUKrOpatpgffyBqGlbfr2JDRemvOsob3dr0KrPAYlH4xtTR0U6Mv+WxOb
9ltewhHdwWxvEH1xz8Iwq2BtYxvmjgXao9abmDCcenz6mHPALIYakSPGfJ0+8/To/7xzwd5cuNrg
Q1WGu82ObaGRQ9z6iqjVnzTkubLpZIpO31Qcp6RwWqcOSw32u8cA9nJR0L/8Q+vW23g5l7lcRRqT
TnXpJ0xO7JLsu7W7/oCYfYVCnWSQ/HHU+Ou9mxRo3tg6yPkqRXWOCRk/gG/lSqiF9JN+4L9AvLz2
qhYv469XiIKQ8oBV/3NpubK0N2A0EA3/ctNJHSrGs7d9S4jEjb5YjT1L0kUrxjhOGo6DsULwBOSo
TA2oFv5Dyy7UYuvDPqj9tr/++TLAGfO0pIlsiOw0N5WelLAIWaoLhBKeJMQEOx4IP2jkrJ0Sg8iY
9dKVYxV8d2vJfs4mzu3gSL2QNsgZ2CDfuGeE84XOv0nS1Ci3QKjni5Cfpo2iQbw6QDp5g9QwZqzk
E+Avh74i3A9kpIOpewaIt2z0jE+WFZ2F7qAIcfIyBSNCCGBD95qKOxeYn4v0/cFvky0pYVZqGLqK
sBWQHoLvgtReMrEg40wRa9cU7DmFozaOIwwstNFkanZCCpZ5kIdOK4pUpMYewd8TOy1GZo0250hL
ErFUMp+rIWEsMUZq+T8axTAPQy4CUm9m6BLjouYZ1ZUycC2hQ6B2nD9RnEp+Afp9wsdQPtNVrMqs
mzDhLj0d7CSzykRJMgPhDKgNpMizIt77d1JifmJJv/9Q9siK4MPF+s5BiRY4kGD+uLxnSiA6y4yQ
0HRbtSHWx4tCUmnBM/Mx2acY1sv72PTuOljvF/5QmL0n6yE65TLzzBw5KizBNEYR0LBS9U9RS0W9
ye/vfxzR5Y43aNla1RNupximtkeY67DNCcjb/sEAaYs/QdM7jTNSS0/zLnP7hrNA448gMTQ/gHeA
o8ZFlNMVDf6IZqlRhYQTw9+ttT/zOxZ04P4HTJyUP8I0sxIhmHRb3llZvZG4zFS0em0rbHQbnkKh
WK5Gzz2qvteL6jVpWaNukJiib4PRx+qk5IrRnnUr0uz5bqAAmlZJPdGe3gXZA0U2Lt3h+czGchmn
wHoKDBjVwxUZ1Sshp5FyRN9APXBxQGcUpgCEr0HPLG6uCuD5iDdZ1Kc6Ha7Zh2lSiB4CRRngWNwf
n9HSsgv5zd7nZb957LASVFxo3vc4WlNLWBi5x07wX0SuWj8hCMEoeWoCNCEOh1gn2ozliOUKOGSt
3QbKSon7y6gX04/WItH7PJGDqT1QsEg8EFuwIvlcGcwpm2Q5jzqAhBLbCPvPBkdj8pSg7lYTmVty
PNvt7XeVuQTKlSeHfb/7GCkhcXGa8UkgWWdI6SD2Njw2D03oP6nzDuxibPIBuppNTMo2rkdZEgOv
1pPgTfFBG6IkJ/zVTZ4J/pU31vxdTasHbX7pZFnHSwdOFiYCQ2Wz68WmO6HOvYka/tF4zKdhpSuK
6PuVfXJViTH84Orwc8P9yx68r6oimu3OAvucdndFgrp9g3OldLvq+EEDdgHbKmXHR7REa53Vc4ks
LGHwxzg9IqzgYDsVn3AvIVFcwFczpnkv8IVnbqKbBTfURstd6nbjkJiLsi4eLc0zNB8a/uUQ4Adz
N59DRbJMhLY7NC46nlso6n+ByN/XnI+acOrT1Qx5zo1frZ+SL0YSeVq1dSnSUjwiwIa4Ll/RLcba
oMwSYUtybxFPV3aEIzUciXpZ8YhKyuvlpaezMfQLv7l6cUqANiCxMGMk8ArnEVRgtgALCXkcmv7K
tV+CyWAvpQzF68qb47lTaToDJaXwkfDxWpwm5d40zjQTMOBzaTPGQSRcsPvU1Go3yB55Jsu5bokD
MTDX4j4jgyFTS+mIRLoiz3GDrW7lrKsZclHXdhpExMrtYBYmYZTTIvmPoalEZJbo3Qbt56/vAllT
xs+n7kE/b/BQgKEy25VaYd/IRMh3QRcG8E2GLyqz1Rb49vdCA998J+u9qtfEYey853dIhakVoGq8
Cu6QI5PgDHl0q85CPkHbZe3PdRKemW/NYtqXQxiqPsQxQfX90x0ZDluMb5LCxBuRSPmANB2L0q7D
t+IiL7GGuPQQZhB49nNIlrKrWnBQpOdb91h5wekdkXaGxGq9H8QyPOfy6N16/Lhf55JYeIpW46MW
HjV8bbdO5SI2IdyvjSK2GV4A7VhIOxoGHDZJLkT2zLnhtdevZI4G9u0wXDrLSk+FqFtIswj71riL
z85go39IjL0qWjPsZpAm++2r1eTuKx7uUruiBMjHTZEA5oT2Tm7GWpOqjb0UesHWr8aZI48/FFPO
KOnmPtekY8BRke/uFu8DFcar0LMvhBZ4HxhcUaCtfTgrg3bwaNvvnlBydwo1fgs7PAnsqtG8oGDe
ynkMzVLd1toKHbSQOZwsSsTiC6Si/b31petvWPr4f5tH8e6S7X9UjxuH/hSY2QJ6i5Bzg/Ku3fXR
r89zDSXecxv64dnGJ4nA0l4fkkbGcm9+1bXQNvllTliXiNdMnpYQcnjaw885S0uYxpivq6Ct69Pe
9/pxtThwkTlkSMc4adciY9vRQL0+emksVQUB6UCq46eMfcVYC4AnH4x+lRxL5w9kveJ6DbM4So75
Flc0c/RSpAbbd6aK6wtTqRYElN24EQ3xyIggTrjfyoszsLq73txDCdGx3bpIZfiC+FUPkAeYzXuQ
d0GnMbCji2g5CdipWrqJXe4ybA93AusUTSd//a/32MlOaOJdDG6MaOdoYawuaaFxLLfhhGlflQwl
H9CMhfqmin4nZtJilVHPfCWddmDrv9zJmgLbi5jFw6peUrQtzNq7RUzuBJ/0KTL4Mu2pRGkPx8ag
rQDOUqpDyylYGvromdxrQybd9i3I3gGXiiZd2o4IB8yjjjkYdu6i94yRr1Y4FbsK7m1Zzgyqzq1b
ciQbIO6bCHU7a62vnFbe2bY+Rhjda56ImbeBj3lbXm3RXx/s5rxzy1AAkNv+NrHo+K7sUCRq1ZDd
JAeR6Ruhrz398MkCrl0KLsQNHrxGyGC+p6fSOO5ded0fyXFsdiHs4QaQ0MeW3A+7Ec/H6mGtyunh
8qmpcukr36nqYS8SZLFb5F/7W/EK3qKXl+umPDJ0IpjFsHIQpzTLFP878tAxvnCcBjrGXMKyS2qr
In5FZXuVPGvvd4G2Fxm0HtMMdO4a2l3zMIHn9Zb39Ot3fX/Zlj/2UVC0qO7KJ1VU3rAvP7V/MdJu
bVyotRAHLtQG5wB7++HRa51ouWEJlxv4tgKsjbiZHY5brvwqs0HMFmlK3Dj7jJPqclZn1cSuagHx
AzP+t7a+vtTTUK8lp8Rnil2QVrGxVeOyHHJj7Gkv2NWLnYfWz4fSGwm+2Mp3ft4+oYsO5muHhYWo
oz4LBlh2XNaCAC4WVYguI1o3tGUDRUPuzpqtchKqsCLy4CKAm1SSV9i44dIHqG1eCkka965OtiFH
nFseV9d5esE8p7XzitHSjV4AWYSmYoXudgRi+bWOMoIm2PmDLJiicy4F5k8cDMMPEmiiHiM00Nry
iVFxeCSValpuzb+XqSRxMer15uaiypyJ+EiFDnsTz74xvkqDQGldIqn9ATXIfMM2EizyZwha19nZ
Ar9Npfo2LWMsKAc3WsNVGiynMoS+wNMJQ7QcI2X5MbvBYZ7fTHPoOX81QCBZv8W1u3I+JLcbcMTM
c73sCTNdZBNYoBLDrWT7a0KywtN7XUTr/odv8IVx77WHg4glAAJtyJcIbmqB+2NVBK7s6Z4/pwUj
ms/RSex7xPy2wiuW41Pobh4N4a+KJWyFgwjcQ/xP6QWtGS7x2QRCWx8Re+0nbB+Age4fkukb/JI+
ckOL9JEEMUTx4K72s2vUCN6bB1snkVAFUcVzNHJu6mBZ53okydamGlZ0k+4mjpn8UItQsTsKua9H
KrfKm3EYllcvYrgFv5TpfNZ3hvxEui0s5duCn998aP42Q/JsqrDHCwWqqsDGxtfTGCOShoG4yIoE
FsU5Q0COLUuitq806uQjDQqGNxZqJYrughu0zbOVc0vZct/e5CFgF7H5jgtuNTSUeJ7K1lCkpPc6
pnzNBHuabwn5F45FRY4jRK3ig/LvZJWWKAXtWBE0UtLi9+BTxHA6JWUXR7iArXYw53QvjwrnAyZ6
Ym+jI+hK4VoQo7ZIDpACD4bLMK0q2FGODYPwDRdm93cMPNRFSueNISBkP/0xsA7w/S+1d3EXj6ab
1gH1gb5WtilwlChGZKKjM1ZnDctlqDNx+EOVpzFLth6tHtUMTH6pjHPEsn0COHfXQlFsGa1pUzp2
BXqZVAzi2w6P12A46HTAxQQIg3epMyOZtd6FNZ0lcO4KBVC4LGliN/IUMH+dLhFv2RAAkAnLnvyA
K6YTFYWrkePUR8/i/g61/bgubJkeKHk2mIlKpYdW6EJTTnfxIfMXgmnaEq7xgM24CnGmfWFuy+Yz
Si4hCX+gTbsgRRf9EB9IwXD/mAHeKr3kHOJ89ZVmm85iSpgYbEJ2E0SjwVqWGyVHK+k2w5SCsikJ
eBoiVmz/+r6E/CeM5czVUCqBla7iTnYEdesdvRf+6C8l1MRN3AWMJiGY0dT2ofgMsg1wZEHQaRGK
5/qqvkXcO+oU4415HwmrfyryaYQyst+jdvYdSU7+IdqHW30R9aZMny7FNkLlQ6hb1yPtwnoKhqzg
deI6CBBVhwuodILr7v6BCWNEIVAnSLqEzBd/D897imUWyk77ErLieS7YgqIev8V9SDYBY4oCHmHZ
xtZHXjY+dH4/JSR29ecgOAdLxrhlOdLDRyjSzZlCUS8/C1g8kngKsByHVlfFswgjntQmgCdFk5nh
5/4nFQzdq9Un3HehRLyia7ZOJfKmB0PQNMPdJ3L8ofwCmo+oY9l/YigsX1S2f0cSo8gKCN9aUJ82
ZxeXnFlazUYjdeSSGIZkjtYjVZdI4I/WLGmbMwT/kdbO4qKFhwP0vYpOW6FWi2AUeWN+lWinV4Jb
eGd7BFg/dQqHlUlxvLMmrF/c07i2QfaBnYoubAMZ7TXLWMr6J5S0f1VgFY793Vh/fAqpRxE6+gue
ITfD+1v9dP6FTgmAd1qTvkPZoQ+ZuZq3b6fEtq0izXblii9SkWwjagZSj1rWKjlU2j/FZcXPOkTu
E5V2CaAOldLgMyr9VDsheFcc0b04fGGcIGKmU6QIvpBrFyACeJHPuEOpF14PcD+K8xYN98a7TR/J
eINmTos8dmGInImlYcOtMNDDzRbUaGmvuwsXbR5DrBMEocrPNGhAVKjrLKCjZkQ+AKLV112Oz5J6
ui9prdBRX9M6h0BA1N2yX545vJTnGwp4WDHNwduD1sdY/N1UWoMRU7EsKvBkYYwXenv+9jSOBtZj
IHNFxJOUQhfPP0TKy+u336/ynMcULoFP/gblFEI72E6PKTT9/JiaORdmip2isOuwhNb6p+58ZM47
hdw9+BjaPMeNsA6OvGVgRaj8QQu0Nc2y+xHhvD0xvCCdPETgdhHM4oGc+MntyEd71CG53pED3xoI
mSvHaDMcNaPlGegZvIxAHbBQqikg34jzjvsfheVhrlBCopIRHRniZnluOEzpzD/KK9FsEQSuPJKK
/zFVdo+gO8MRHUS/03gPr/Pl9J0QNfZAHRAfIoKb9hzmlTYZyfBgHS67KzGrd5+cG7NIkCiFE92/
2RPm2VgRsTro1S4wZWw464J/+u3P+yxroIYeEGpch5PB0VQaCdSSY3y90vzuJov63zEgSSWvBzse
GyNA523AmADi+DRfhJj1P3ITTEUFvi1I+sn0wVGACNpNHCLa1L1udwn9c7ZmYPmJgvFwmvTK+JuN
Hp4YpeQCuTAi39P9VQVYCyRL9xNIQA84DQw4l1XxH0sG8MLgTdyjwapeXTDQ3Me+ZeHHCwAuDRpI
x29Psjx97f1V+bVi4FWWxzrhOxKZJ+w0vGJE14n0MDGRA6SMdMyPAatHaCNtiAtpYTWVn9LtlcyL
svsEVx9jrWOtZnxmnh4G68IJOM3mfzNuZZHhxoyTMnmXzSoUQkFRbCq94hUX3hMZcaBI9VAWiZj0
SicwIK04oiKuduIw08oVJwvdyygykGz8k9iMvddSjoRkEQyeLKkZ/Hcilexyv1AfLIo2NhQQihqi
0tSDZ4KWxtZqhE7+m6K/pjs9/D+T4FuyulbEt9ZZaG3QqDa7b0y8UIvSXp3RPa61f036Uh6MRtbv
MsmWqbbHSuMei3xXRj0BEDn7F5gkb2+Z3xT13rl+KHNZCfXMtxmYVzctnXuFSN9q2kd8kEvhuvFp
KvMjpxV2Zh7b8RU1mnTS2tdqx9UoDtAuPz44cckZ8vxWKtt3Yp1UisfZKL3duAb4bUXnjYHcQN02
wmJdGs/URXxXb4a+KLKF65NEYVt06xdkdzE8ZYbrSwZcg9cqLKei5CEKPZl1jtMoIRVURAelH9TE
9OuO7ZCywZ0FLmI0uEziRrSt1ApZP15tYNuOLV7SiCEAw1mvJEB6ZRMdxh2E70eKMVzufG5/W341
oO3goJifs4zo5fhDrtAnM/kcvqW7VlEEieUEXjFOoPX1FHrM69zfLY83sg0L++8TMNHa5sRWQkb3
JoU3qr9AUD9Mpjl5FDEwG666+WjDm6Jrbc0w0OGC1PUFUXxoJiK5Gqk7mw2dfUE51iDFk+d9hf8v
LRP4IoowKOs4dhh1Hi5J1aJ6drGwNObA9Lm/v0FaDe+o6alTg1RNuxOSjaV6GGoCxCoqAE2+KVYp
nbwsQzugnj5GggFN5/93Vf9IRS8FUw5GDDP3JbwTztkyrDoSvml4pNHPdZlAomxACygPRaf1tR9p
K5qF4dg7MF3x9zUx2zXvj732JzsvreX06oy/d80ow97UF3kAEgaaGoi0CiPpvQQhkyjmf3qaF4uH
mkN+zCeMhPPJXKu/MXCs5sVC2RKjSSI/dAO15+7tSsIHRXOPrjTjuU5MhIUenRPosgwiikkmWdN/
sMfRk1CcaqUvY8ZfVBWxbAxlRNWx+QuCUcxRIVlevYhAQgAHCNKK8qeUgKpFpYMxSpd0YIrzXX7x
SBvkyRwjiILvEOxZC0f2mYSPnPJaDzXt3Py9m+2++9gt8fuY3LopQmKHbutfXZYUbN9nXDjCFCec
ENmD5tZFKHL/QN3q8iTPsjj++A/h89r7yYWq999awMCzO7n9/vSB85pyZw5Y23EdOn5CDth+xmUy
R407qogok4nq4+LpHNo+SBrxYjA+V9bUB7nA0bBxWPoWCLAz98w60xSY1ASCwttd+FsIXq3w0JbD
Nbk8U3m/VYQGO8bV4FM7WPoReW2qjBQcnEV0IwwXmAh5pYm/8BJfieXFHdH/Gfs2Oi09KIgDnVmv
iY3zQIev0xqEYBfCM3/VlRgrY7jIXcpkbxxLQMu6B99QTc6I6eyfIs5z3ioGm8RJTviLmmKY+//Y
CrXm2WzUKj09z/pR1bTC+BROOX7cIhmE2Fy6HvlPCSWdstCQVObK57j2SX4heW57NZynmEvuCasq
+k8i/D0DUy/kDi1hNuJhOyVs4V1ShJEurPcgDFYlcAag3hZ50HLg2NE0gIqtt4ospexM7Gjxv+AN
hFIE5O98NcP+Rm3S7V3u3gK0l7HOeT27RQ/sh3vgA+EGNj4JePtaLbhunQo88brzC12WNViTDSyw
TGkXH04u4wdktWWWYnwORIpKzjuJCPpZ6mlsQAZJ//270/00BXuB9L6jsX1mpyofRUL+SCZRfj+B
S2kZBM2gyBdgzFk0tiyQRnjkfPBVPGkyam7TsmHRsc+DNGQ+ei+nngGvWdoU/3hP1rGVmNybIFOB
czPreTRM4MuDx0MGhOsgNSHv9XVc68NhBbfXZUZIlep4Fd/MuHHyJZk9/vlWiafhhIxhCsWfamMU
BvbXxNbHimQ5N27Eyd+pl73yOX2a4V9ERAnoNvEz12sstmI3TARpKzIHAYtnnI5q2uiyWR3mmpXX
HLMCRQ8kY0o7cR3yaCc54qkhs3Cq7PvgYU3/mM5JsPUhyeDnDwABQjJAqoMQFtzdvqNlDkalwDNP
OxaJmwCXgZWMZinbtNTsVumtaF1YNGC5rnyRBWCkhfXOkN+OrSy88k+KmQ9UkycrXE1B+/tm5ZZC
mAhE+Zpiig6D4a9nqJpXLn1erPmfKFhGzKnMLKyAkEg92g+fdXp0J21vTyrJYRbTSXCXn6FRIj26
NCLPzje8i3qOGtFP4/eA3Pi0SV8f+JAyalz/VMGdXMxgjvbFPfN17o2HR8i8buvGk5QQZodqxoca
RSZt7A8O2wO4HSlbuCGs4JAcbyS7ejj5BMYXcmLsx31buWAFmMYGviQY0piAXBL3gBBjAEPhzGsX
uDqSTUaF2xjxQbuP8Czz5kzqJ4VVx2/7S0rfC9mxky6k2ctsVytnziEDZmy6niuNRatbVgBgZNIu
RYUucq6geoADZVfPRShqcaV/JR0/RAIXYeDJ3nkFhkEL0ECoJ7t7cRfVPfJbByPNX9NHmQzvO9zz
9PwJw03X5ZlvdKLmFm9+mjy+8BK4eJ5aIQ3Smhd8EE9eU9yPy4UVJhon5wIyOlfvKvQp+mcW5X2H
KoHF0V1AJEjru035SW6iYahGHfEdOFAMVC/AGFa3uDrStBA3f1JruniBwASoPYq7nRfkp+AfNRIz
zaJL7kpWEcPX4VImCBDVJjNQIlc6n4TE8V1evvK3nbMxfe6p43jeuYN3w8VZKJefKze9lSJrXIBv
VKPiybQuqn3/TCBsT/OVZJuT8KQvcAL4PE9Uw16EfRXpJr0k/dfjX7u0xDhWNF4HfnvK68o2iQKh
BUoYktRVbK7HfeuPTTESuMGj7ns3Ic3SE1nmWOZmt9GWQWKWUCQVmGf9mj4nhmSYuzMWYtltLecf
lRySohtO95hkzGGdg7dccQ19aHINrFRr+s+EcJwEH0ftlUPy/Fu/dZGDqcntHX/fsQIIscQxZUsv
8ZHcpaucoiPKZZ/vHDg8KtC/Z+VafTc5WMNX0RPLgTxKCT93qTfaBGn/ZGQd3VCxQ0gAHbftUUtn
2W1H4UtENzujTia/GfIYu+eD10J8gqY+rZl8BsPcSSl4uBSdjQ/CJkn52awspy50myyvHsK7IDbG
nSUVra/2sagCWu3byOUjC+LpK4ZEAaRA3Sprpjk7ZlIKCFpd6ZyYYhPQD8EgrQWp31TcGbI1bM/V
fxNYoJkZ+DDOcKKohg7ALl+/pvnil3kPWdA9VOIrgvVS3w0TdM86zxxnT9bRvLHQBOGo5dPeHRS/
L4cNb1sQLhsj0Zw9T12DS9j0gyd5lL0z9qDc2S0OgQEgv4r85/JHA58grqtUdhRKAKhdblxGdqTy
a4Is2gzMwu6o1CuGjmvt8zjc/D3hIlUyDvAtIzST6qaz6QD8K63RcmysYP4vlzDJbTPDiP2459jY
v8U3si5fewa6oMQlI9DvSHgA22rXiXTHQKey9aHxjNZS4lIJOEdATYTeay6VT+c3SqA6E6l3hN+n
LBrnzn/YU3mWLLwJLjLhdcxwKQs/l1dgSS6k6TG0zdsNFFGMcgI9+nFHfFfZXKUbbKf6Gtc1NKhx
O8hlBr/IW71BLqmDjNi+uD5dld/wbevMyvTNQ7NW9OpM8GTEnAd452IzfyUadsA258wF7gucsStr
COC3iIFJyO0AGpyLL+UpZ1G77PoXbKaj2WnEObjbeVE1ZOdmRi/buExgKUR1xuL4cHEu+YGvY5u3
SB52eo4cB/xbFdXUuZVb7y7ihIjN1D7a/gllFdVnndBCmKERVRF+WS3k82hq27boNv6st9A9MHmz
vgHyJAUsT6+YNhpqit9xVb8DXlbeZhUqm3aiAy3Y20U7JehlDls4F3T1b8RGZ6aKFPOIaCZAJ4Is
FpqeHVfKhffulPik7zLZoBZ3KEREuMuJTaFw2mFOU8GYU7O+WMR7MPot9itkJF6VRT+6vPVpwcZx
kh4A4KkK5eOn/uFa+Vn+jK/dnMIJ9VVi7E94t10RNONLxiA7mHDJJdfdLiGj+1Rt2kYZCE0knEQC
Fm497TwUGRzzYuz1B1UacVYufe2LbH+HQpYDz693DIWwO/QvrdfUA2PEm3e6rqhk00b8zWdoQrLt
t+ubsO4zSkYvVRgG7T3wOevLT0iX7fG4atqslXIyUlghmZaxdln1eQR2yTNnpVRBwqVTQ22NyCtb
XPFiOQWY1JQqwkivYbC2uCcdMZD7h5tTL7n5rb6HRzId8uc0+muarXECyrW35t7vspZZxns2wNHT
WaftPONjbbH/WAuoGkzfifhYhoQqTdpimCaajvMSjC30MeoVA/0wwdHgOX5ZF8hxL14W25L8uDhg
U30vXsp9gRZEhdGdRPhWZ4Y92yG20q3v3FJSbjsBnN7pnVoYhm2i3n6DO7/ml4G/4Aod+GRqVDzy
ltW7i9n7pvgi88u4lffimug2XkVOUJHlZTHiEDt1uDJSNfwoDht0O+3bVSGsJCj6ZrnMMeu7ijq2
ZI2TAf5j9TlK7ti0QFKzOOvJAEkDC4wWryY+y2Tt1dPCQkUZkQvrus81141qTD+WHG625cdPU7Be
uOyQezC3SyuVoM0Y4vQ2zY1FDIsvEOCPvPDSFSY96iDQ15AF/zfFnycTTdIeKd+PhrKj105ki6+/
YfZPWDacrA3MvTyKrKEwBBNFrE8tattRXMCpovz47fmpwyWFcLIyAn/U4sb4t+dyBvyKG7HTwURy
cIuV036q1WfLQaTIuaLUivK2ktrLpSQsZ0CjdjjFe61VlVw36Ez2WMvsI9YM0OEmpAEOQ2Tn0HBC
TNu5sZmn3IkPpdCIPajMV6SqFxy1qMSq80XqTkbTKMTvl1ABirMDxCjIfUAgB6TY/EDWA/amkgB/
cv7tpFf8Xoksv+iHwW/vdic77OxFYjpHup8zh9GRvha1/aXiRmRr6xjhpZwetmBhh2l44kTshio5
xm1UaJ/DOKKf451o27LyIxRQt2oew6ydo7gp6hRmDfdMnFSeeUHKIHflQLQua6ZXTGgyoML7gQZh
4++fr45+sDOzIFI/FbzxIJNLqhwt1V5Og33m7D25rdBnCufQcvZ9jgJUcm21UsEbPDAEYakkZFd/
wh2gyJFClWmRjT4f9qggR1/S024m+WEZfe2xkW+Ff1TwqOa4KJxGAhRsWxu489tFSGHv4orziWpU
euEz62sceP2IdSaOgy/A80Lqwp3qNjiFuJ/USc566q2mb4rDln63tdJkemRCOygxY9gS/epJBKJM
zY0t9PiRENGeAE+AQiPUQjRa20xvxELowzP0qmuha6MhJzlCmyBFEYxIEf0I17dqQkS6ASkb90yT
1/hKJMo/GlGrLqafu31Z2uKNtyE49yWhSxHTnfWQp06sEXWiMt1qBf+snpYhMtb6djVdMdheJUR1
J3mOjn5w51LoaNIEgBh65Wm3URyVZJBvNggqRkaHdyt9AN/dqkaZNsvNz7AAgvQ38eKeZku4Dfcy
bOVKHL8UIwA5CbTygxdwga9KpUfGFFg7Dh9l8Tt4i3C7iS8cLw4d+HiDwW26wltqxX0q2/2AMdr0
K1xl5AVxKYeXtmsfOevHuiw42+q0cLeXSiDQ3h4hbGvnGdFfbdoSuuwE1kk+jCpyYv775kAiq3iP
JuDXa6ZmNdDFxVKCR2tqyZWN/rU1Uz0mP2M4Iki3sxbw0LSEjuuC3lpUYw1NsXU1epRdV0dBOxcd
r3Mf5xQ2YXLUZqN/b/LtWWPM06F741YpaaYEl07D0octRdl3Gu1CuevbeLf2TzL1wn3FvFu8Gb8K
NYYJH1aqlhycQBwM7KCAr7Q7qmhTwWAwjL9BZnVnwUyfztQW+pmAaQe+NZlTGZBwKX0BqK2E8ZlW
W79O+YBakEjsoPlEBtivZPeIyws40Cu+TzaqtLj3ZHS7jZG6+JPkb63MWyhb9OIh3/QVVycX4r3A
FSOPSKS0Mff/3ijESB7VoT8zTgxEJ9jwCsyGD9LgqTFTolPetEWdpRRvyAN50AOyI0fchLmUxlic
oXhw4TLA5k7GBAwUkuKGbPYKevdI/z/LyU0a1zIzssmV/rbyFIj6VXzk9Y7kCq06wfYGnFl1svr6
lOdiQn9cV/jpE9MuELf7D96q8ytPDPABzHDpQoOcn45G/uOBTzDacNNZg+GxYu3kWJovspy7/X85
xnVCNIN9nVdzW8c3fvtlETb/7fFGugOsOl/xW7k7iSA8z0P/sqImvpDPKEdVg8R1kQqWJF9Dsx42
q7q3VJJBLl4HyS1mDGyF6TqL3RitrH7/yozcg7bCeEpcjiWMCYBl0M+5so5GoiCtffVpCH9U0Q91
lA4dMhRi8QAJaiMZ9v35V2WSOsBH+/5uI/C8GOCWONmt2u3TUGpUCsl0ZDlbOtWV1HcrmFcUHBqX
5ezAgb1FUObNwhksu+H1OGEi/NxUbAtP0OBmb60ZQAaEJq0pCLHWo7xifF28L0scrik5tbsEK6Js
UY1DF3I+X+Dr8mIJ7RD5Iie21L7ZnI7tT+lre177leGCIxkZDbwtDWLYOCo85m5zsMI3FCP/Tkx1
d3QVXP6Axv2MfJ6K+2p7NCF18z0TOZ9h14++4f5Fy6nuK8JQzt/XWI33098k2R9/BEG/5YXAR60u
3TUn68VLSJGZml2BSKBwvbG4xMp3LqRE3wubb0clraOXXn9bewDQ7Gwtk5/bLMhcimAp9tb0pGh0
XNvkvxdQ/aOeKjw0IuVaOgEnEQv5YMxgQL9dG2iOHmwCXMl6mtUuleMhViGMTpgKrovHzJCTIJN5
ZAXJOQrmPOLnq4wSJICfH9D/X+jICh/HtcetXvlqenlQ3gzTrH+6OgzkwEsBlNopOAX25xyhokbt
hf2gufbcJRBb1VewBl+5TjSn/YwWLw5SaPpWpX7N+ap/e7IS8jHqsvH62Z7JlYg4zoRMIr0P8T0C
2QjNzAL9u6+V0bwP501j8hQSSepbw/UF9mePbwaO0AxXSnhIN5x11gV9Nv3e3wLJM1mwnvkXlfuQ
0cycictpeOTY47BfLEXLaX5NOtmtBF3d8owqshrawATQQqs8MQ4L6fl4M6UOx9ZnZCwfmFyzjrgq
URH70B+UseBgmOxiuuy98sZoCZZwmvdB3dmmJOG6cFc32ifdtc7MrKVMsTbXYmBlByXFgpGYr7KP
n/YeeVG+P44jmuTtiitsBj/ZK/FqBx2wsSu+qdbSktThuLJsFcdEy2CcYeW7DEsITYqM/+4+LfTf
QqUsQEOw2dKn5Yfx5L1Ih5kxHsaty6uyZyI8g4rhOCd4awWUpMk/p1dV8XYc4wHs38M6FQVeuRlJ
RNj+qwQdMEX/EUJUA2zwkXREWCsVY5qvnyMhS9K09pZsOSgA3f5sMK1ef86LQ7CYYLdO62qszPfh
iRJoxU8dbJ4eB9r9zzo21iPZVRm78cfPHRQ1P7vVkdoDwpHYLoBtpgNLBGpN8QQkGZvJQTiVGBlo
NSwUXMi1e7roz07jbWRhQa2BzzJyfxThmWWb1VE1V8OUnzvE78WH74m1vrakIBcIa2Drnazk2kxx
UoVkYkXj0LfLjE7HUN9tcko8xEJMOs/ZeKQTw2Exwr++8FzMQfD1wh4asTGpq3wnRe35Qce0vThz
EQW6k8klHvH9HmT9jYzd+ABj3NTCW5V6b0Fai0TkP67LtZHihyKONQn3pwO23nRgsvINFBc9Bm+m
tVwDwysDEyn0BbqhPCmoFqJdnyt3RpO4GlESGTcEKVzpinlrT0N2e7tBZ6D/pn6kz3HExPEMKXNs
XyuGBJyZpooygBX4PToTlzHyZf0LX3iyRTlEK+yN81FqsHQVTNIlDSNrobimmCMxgvfyHN7cSSyb
HsZh1BM59FK/I2aiTwUhDf4DNxmIP1HSRzYitTVp2Z5ukoGVHyCU1QtUZY0NhJiNnC4wfJ4Zj2sw
M+JeGlOGeXaaGwcp1N5PuEeA47iZfPTSbaXKh9LIvf4I2TiiVmbxnCqPcVXMsCPYU2bKkPvmS5HV
8SC/ljjaQjWOCz6isSl3sxFDSAvVIvJFdIhs+yqMGuNjGHtBUdNBVhn3VMlzGr9IuCfC4wChbWYD
ZXL6LXtQ8AiPb6AHy2NlnmzAVQQeTP6n9vkHvcvIWT489X96Cv4sKuh0Bir/7CB8urE2zK2lyXc1
b+uyq3WULV/8cDq9UvrkGXp/2QgyEqeHM5+EgFnSuOjynPGQN5r45oqNyb8J948fa+lcGxtiizx/
Y+pE5h+gapbpNQBfhayuXJ4ltjdsijCouwEchfyD1B13DzECkMBV9zo7tzdMRHGFlSrCNR6+jAWQ
/hJeb9/wQMkCfYKV0FscQgoev3d2JFUFbHnWhw8vfA+/+L4W01tEawuTibXJz+ZUc6RZnSNV3gb0
e3njjy56fl5s2b663GtHeBUkg/PK/RScZTohIBMmT71VMA8sjMKQxyNV+IsWZx9MtHEo12Q7WGs7
LanIOftCwQ6XJ39C60OJ749Cesrz7loHtV2/V9M1VyeihyDGYAZ4vhQWNTN/kjbvLMlkqMHKxIUw
PxnsbXvxLt4VXw3zLIXdRPRqVF+tEPh+k/OAX0PZ7cvawOYBpThu2XSpKYZR+emmoCns+iex+sip
J0Z/f8OITuX8hB9yBTIODijLFErMpE/uFH5AhyjrnzuYms0cZ66CKujST6XLDP2hPtqhuZMRHy29
LmzGeX9MI+BgOFlkPxbCEBtvLpG+iuhlRpLzQyZhxHjeTpy0nvDYgztynvzb0vAKkzWhsffX0jrs
0XHunbDg8aIvaaj6cVco3Xbe5oQtbGRWKkfJ2sAZMzqtHHgxWoKGUcIgh7ntqHgOovUwTB8VqDHF
Pn0buFAGc9lXWG8OWfCQOQUhdn9W8mmN8xR9+gS0JO3FIR4ouaqr0r4dAFyzHGZmFBF6buSxjam0
D3Egj5d3z6+f4zqrNk5gQBJLlk/3riy1fRdwMJVvH8C2swlhejZXhXYIlo0g3zZwnlqEuDWk26Xd
zOaOtoub9YF0f/ZbUlVkq8RY24PEfF156q/idIfs7VWE+aj+U3ALh1uQ9GU4vFzZaRHxszaTaTsw
ORbiQnY67nfQZFzApKQv0wWWqiEFK3FCjZT6T95El0CyRgF06qncws6zEAK1KcB3mK2Nq28tRQFp
ZbF8+UboeMnj1teCjR8RF7jcjkijZJauCrEIgjDSbroeLtB1L+EIMslMINIRnnI6FeqBC9Jvo6/W
Mx95nn2o2OTzJiSAGzxf6I0ncqiqSL4/CQunppLd9a434TlCvzKaxSG9dXyMAxwRRcDy2NfY12X8
+tSZb9QcU3y3UkE+aME25SLP0DMCbm3tgQWGR17rSNERN1AWS/a+sJPWhnm7Vwg1dELW27GY93V9
BWqE6ai1nfgWlfzufTnRES0LWvKnI6kwnUj8uyy/0b8zSyXC01Ou3Jbc+JCjqB5jZwpV/wqpYqYG
EnSaQ+KkjUncgdy98PzFM6YTBs9+ic9g/vRr9XzDSpBSq1SuT462sQVnkjjVx6aE1IjpYFTzCo4u
uXYnFN3DLs7SSbPGGMBQG8v18wUWa8XpxJD8njTzjbjLZ1MNA5MW5wux685VBtelKhPzgS5BjiV7
9p4E+ZiI7DkZifG/AkGFzAAdqv9yhhN2SuqSIlrOvndHENXBs+/qj+M+puF/lk/3W9kXvpIwHCxI
H+xcC8ie1wRG7W2GLTEse79j2TxsaKakCUp0871PoC3iS4TJG2FyLIEOyIWfCLlsoHqyuxaTO40u
h0IAScC5tOBvQIwsOo9zN1H5u4aH6yGmUjhMIP++C3tIv0kIteZpjK+it0Qqh5UaY3SRRCJt4xQ2
FR3GLQ+L4vfQe0ZWdMsp/GvWxr+/JECYZ+Yzxdvoj0Lv/zeU6XQdVC4Xw3gJNjwcwBvTjOZTV2fr
91/q9b+vShNiYXmJupi/Yk2zkB0wft9fnbvuPgzuy7Es+ZmChcNSLrrnITlk0iMFAemM+vRsRhLv
iGk6Z9GmzkFlzql8b7DWLal7INaEIr19lrTp0b0y74oL7Lc04QPiRFkkZwbyFHaAeULgO2x710rO
ihBlpKfHxE7WYnFyi0NE87UHwC0XmtYVNaCR6Crk+eIDEDzSkHSz8f7PFqOSEDwbbct2n5kXudHr
1cEmzEefi0UNBS+Sl/xmX3BE5NpFquiJF7oEft7Tubo3Nz6p6yAPRGBpL3NVqQkiT761L8CERI5z
OKyXKbMSuQnU1KeGsfCBKiITGIAf4ijlIhSEJJVBwoWcRMWn93P3yPmeChQnC/FYr91EBNcRt6A1
9ZgTjiMmeUGkFCph4vZnUJJg2tn4MkuSHmKIFh68azPlAGjrudB9CPhtzQx909o39THGYoBmP3ZD
3pMwF+ZxKNjbezgbLSR47EZLj9nlroPvgobE6UNib7836uzRWPPBy0NZOiCATMIzjPfviKeQnKlY
E3iN/Fu+SZ9Wf8kR19KDUSV1407zxWIqsbyiQ9DOyIafd9IwAUa9APTnp1r7hJYudJXw8q3XdKqF
lLfdWu/iJAZ8mFoWr5zHvXOv6W7f05j7BflB2kQmyPP2c/w0w4R8d8Zp/lJ2KUiFOPogFm7FlRBf
iUw6KE4BRSqVEOo1pYTam9JpI8rOpCzHRY1KTx+OIAbOv3drbpKV7s70WXvQ7vFkYnBhYtnUXa+v
Jk+Tj+lHagPy1zQm19+Pc3V2Rx9lROqkt4mEXA+44+PgFNrEywP593BnOnHzONdX7itYmm9oK23+
GKZvsXBFbVn+9OrDgdmV+IBExz5BU/9WJrA5I/ArPK8pcAB16w1MlVkXTXhqw519NWjJJ6khIVY1
dqUxtwKWIZz+GN2lTVEZuttk7yIMbPDHhwOKBHZpn/szEgfPVBIoGs2rQ4tD0juoOz2w98RaIj4p
sI/TTsksSL66TwuEF8nclCT1mBifyv/cs3uJz2moX6UAnP7HhYd4wflJSV+4K4TsjT9XJIdQWcDZ
ZYZUKEhbwwyeoOOn/0P9KJa0uEKfyBo24OaM7u5VufWBeidN5yxWheP0riMtL2z9MyaMx2t7O+qI
WQyLNXhbs78nF61AjW08nVxak5CjZpSrC5GoJW05yj7LOftfw2vVUpjiV8N4iv3LF7NqcDQ+cqYx
5Lpj56rswHyv/WK60f3kLCv91M9prO5iuw0S/AhYPJjznPyNstaK4UUrOmz1iiSi9NwH+3/qSGIL
M1KkfQNgcMaVxEa2VxvChzasXngn73M0Iv8cnAG8Lgb8xlCs0LsdDtJracJoK/wmGQWNW86JPXK9
xH1UVTFOGhCAopGdLM7hnWp28Lj3821aXRgRx/ncUSB7ANNWfDiMZ8ZleTrtknIvle87XWFiWwa5
EfVmkzaDezSKUgn+xhDUHOPGm3sYDCNtI8yr4RYkhwRwTqxGmRKtEdi/+Hc0fngGRV9YpXNvwfDQ
lm/0EA1DxrOVPKDTjM32QbNaph09nYf9FkE9+87a5xf7gATrZBtaHwfoIcnMW5lNg7wogtazsDhE
q4Pe8n0mTAz6h1fuS65bumb9W29mLdM8tRJl4/5Re6QYmx5u53tKQTIZpPI+50h26k1HvQrEN9o9
qma/yDx0SBJr810jQqJbloTcexvg+i9rgDql9yF0XLMeSJOO3t8zaDR/w6xpTbvXcsUzvPDYVhbF
p0dzh2VAHsWVkrgZVHdfG6a1S9PtrHOp+7i9qNhRD3LJp8bUSs7Nul2+i52H3wcRKkneIQ1RgyB2
x5JkOKATZrANqMNzN5HdDIwycmBnCaFTuvftF//qSeGeiS81b4O5elTz7StAlMKSrqxXmuCaxdq1
/yZNYWvz+/pYVHvGkYzI8Tyfxjm39Hui7xf/mUDDh7JeI5rMA3x1+OTl7whzbLn9D9wtped6U1rO
F6EDCMLvDRHzQojD0QFtblGxESMbidabAvtUFIXj03oNVeausdCwiQUl3z+iC0d84Y1QkGCh7GhY
W1g7jkK6/rk+ECDVFL0xn1gJwQ0ToBBBYvk+akG0UnsHMwgk5KFYWz+bNQAbSg/iPlBJuQbfbfbY
AuwYdEqpIZ7s4RPaLn7NQ9QKGeKicD+pCh5i87sbOzzvMm2pqD1rEQU1RuA3a23R2JxhTkKkR46s
XN3F2k1zIIBo7WgClaje58/ebZqMxSw7TyvvoQW9TibtiiT8hEpmf6rog74Xn31qbPOKMXIBCp5F
UlGCcaivpNMFE0xt6YpFaDavhlxS0ZdT3d891Eef0DPoyl4uvmkjBzVYtuG5TMMaJ/5OECjYMWEC
4wHgeuYr5BlGOg+As52Gx8tAEW0RH+sdJC/njEZPV3NOsKtEdAWitSMZkQmvF8zEw0tlRYjXIkF7
Hp1Do+hQyu06cOSA7KPD29LYVgBtjzAWE0GpiZN0xPD8BFOfYrAAP0p2b0VdNarKp7sZcAgpkjYJ
cYfVgoNam8b0+7ejIxyMjhHztIyPgvV1wEzLhV+Acg5THez4xbD9mnRMfnuvoVDYN8E/tZTtdCLQ
Pdz0MhdriwlHMPjXYQyT4Ks1J0P2P6e+t7YNiNJ9rK8abacASOlYrYrPOeoPkrYxniCs6aK7LT5A
zvyRh9TyxdWyxGqaNStQxWnEp0dk9psCj+DPjBH37PuWZNc51p/YcYwViu4INuWn8w3nosllnqcx
YbWA3j3q2d6ye2ETOy86JcOyRNbMFblKd21c8n1dZMsDyQ5TvhPcwjzhmFildT4cSYbMqIsm1EH5
0KF+eN9tU5oIqZT9rXzu5pboeZtxkp6JipW7PWZ/Of5Agf2oDQAVsGGx+fu4BGoBDUQ2AdLpFOj3
8boRw40teat5XD/d3Goj6SlxjquNeUMnzm9qHOfCb2aQgvnwLq2otWaggUHlVdftd5LEdXNAIx3T
hv8hn7w33NUuQMhxvyvna2ZbB7+jgsZT9hXCIu5bGdptUonFXzx4cK5EEo407wAb7FUAFVYPtZKV
GZVwWZ1e1E9uAsqzKJoe7u6IAi7Aus5cFDKKjwZpSQpS9MEsSZleaM9xquIhBuOCwq7SRb/D/v6n
SwCNJuoZhY70h3vOxHE2hVryVQ5mvxHb3JAXlTTYg9qYEXmgqeIrb05zQR/v0dSSyzNVVoHykBSP
6HnHPUhDETQGFn/+0GSzXGXFtz36+ffqEq5DgEMRAJH6czL9/P/iQDMV7n68VpcfbsHgKJXMVf8W
iVKcNQXL+E5b4CF3gEiNfeHrn3yY/pnq6f61AK3giNtnCBmfztsFVKNlIicE32jti4eD71oglitJ
XBPRLU4/+Sq6/A2ehqaE1cqsqUyjRN+5pWq/MWvZnEya11niMY+Xilp+Em8TBydznsFuRCXy0tOd
rUd2JugpnfRaTzkfuVXwmVbzlLmk5xT13kkyLPnOaAQQtDQSDG2hlbA145AO2VniL8nNcIIQK4N+
sj45jRiR6i0uUaUhQLtXLTjtIqh/qBHfnijgjVmRfbE9zG3/K+39hiyf9haiTPLLYJJxWAbPkpXc
eya8KqOTscDa2lQNpCnB3wchDt3XvEb/6vYOz4dGNg8QJ/SG6f8kmSIaRx+5+oO05tw228R8LaEb
03TKoDQ5PJNwGashFlxDQClsV4xVYsu9rwehwTqdxz8K8haI9LbJnLr19bG1hKSzfRG3tbL3+kjm
e31o5AqGWKgEQQMWes16oi5ePS+iQjUGRwxzzfNx9sz6ImT0R4RoztviT6UfQDKlXAxhMib6PVuv
tX92633s2D+LbbfgI5b+X3wwwacKRx/GLS1ihCp2HyoadVMH3wMXm7T4xuiFU9oYxKcWJ4fkhig+
oYAIPAy8vWl3dQiXUHkMIu4wC4+FdbyqZRgeB1TfqUP5QYscrMjsIIkGjedNqCiarNjTbf+7x4iK
JZJPH3lb+cIsEwrtOxktLlTJ9H1Zffjq+hKpNxIkn79hZtnychStcJ00Oy0dr7HhQPYrj7zRbRLc
jGFK8zn5UOh7Lie/OtsalyWk8i97o5DFtsr2VHrPT0jbluSDoMpApdPuz+teyBNW9KtK68V8ZUSC
gLSrDkVBUQ8DXApmFGRWGr4bmcdmLNPEYY1ulT2aQyJVFD7lr0ttHVlRsRSGK8w4w74mwjAYFgLq
YH/kD5Kcy61DhQBWb0euLS6zi2jHZ7zZq9wjCOKTW94E5tyWNndJG5gZWAA5Ohk6aqGk3X99iA3y
pkeLMB8lKeFHfMWIaAykhPRopKzMup/flYUy9yAT3QtJJgGrJ/EH9BzV7ZiGKpgfPe6oIV9aAwH5
LEEYmgkEJ8gjPC5wIm8CPuwVEs/V1LMtNcaFDvKsG8ys/StUv2zRjzmO4BUsJ2GtgdfDQTnx2isW
TJU1iBaz7IRguJfyZK1GHnXs/ZWhsZr+hv4qTVkcXFQSHswa6Tir5T6PGYJQEP37MsGE0DIJhTcW
cg4O+++ckmcOZaB1VKKO00fL/MnOZ7tIwoB345qgZiwjqpBekGa40zdTAEiUq0PET/KJF7Fv43I1
RjgVA349euwxTy9U5Rn+sppygzNrqEIYqoRQxv32q/QCk1pniWl6DCxehfqepfpDMUJNM5Z4eC9k
kZLGJlJD4QnkVbrd3ZmgqL3UkvsuKN1E2KAiH1eYgDIDRjqOmwOgo4Ta/xvahXJrRCVK58mHYTIW
eD1sqqWTrM6zZxjKOmQbcrSfJdipdw2tmQJKhdUGiEecpQ4jVCmmkYJ8c57XAHZ3eX/8dGM3tIUR
O7loKpLD79WvOMvMBEW+8lusvPS6A1JubVIut7R16a2CbZ4YXBuIf9X3D2HyG+LnRflxTzMKtRcD
7pzFUl5HF6zwA6M36Fguogk2G7Y7Rh88CRDf1zxnMP5PzrGyA8OUSBk052VUPznc1+e6Zrg2kvLP
HIb345KlsStB5O0OEsmvAJD0Hi3bj5LmWT89XBJ95F7i7LKSgai/hFLeJuo2Q6om9NElQy36JDxC
9v2K7ZF2qTJzaqa9mrC/03LYmZkCVBxhQRHjIbmF5D+QZknD72HpYzvcfI++OwUB97dPEF6Vq0uT
+8ZguoGBD8XIRNgACbtOTogQz4EF3j66QvxqYfkBmIGYbNy0l5hZWvy+mrWhvO33wCjBgL9Dm1hQ
SChXuT6/uryvR1VX/BXzdU31s3Qyjps7gVM3qNbvig13rCKEDVAJasc4UGLgLH3HP3bfhgKjZyOo
zTFtgq079VhyKVQ2to6XiAZoULBOHV4PPPL6ame3GSyw4aMB3h1LHfPoKoH6Uh4+JRd6cJatHUX8
QwgypQmVfGyUjcg1cClnBEvIuA0uSp4LSLxmVN6i2aVTbNFRf+gXMIgjEjsc+S+dxWSRyFIwLoE/
jPuEVHcnFF+MGSYUG5mQUNOn74zUpo2uhWaQFcDTunaeiW90i4ohXJZhgSVJjrZxjYKr00h8h4H+
NLqVH1TsQScyxksys/c/ZSTYd8MImcKejp3ui61UgbKyo3b98YM+F4d9BNoI55Jip5EdAsDMOmXz
AIkHOn8m7uhHgDcXA66/NEC/LH4KyPltiB6ZzH15tHi0KQjFd+pujziYLX4QI6Tm0XzzeAQR67Ck
ycRyroeyj2cgCnLxYKKl2YkY51eUMjfrt1Z9O5xlSxKp7zN4360l88EmtZOZp/aiG97cgDjwuB4t
OM4ZO+2sisi6/RbqrkMjDDsK6MkhgrwLXO6E0FDX1tGKoTKSUL/l+FipNmysftpins3N0e2T34Up
xOTBj7h8VjlKKHVFRkFEKD0wIbuCEbtyeivvrTKRczA33GzbHTRGBiN2reBXIHLSNNptjZKca0I8
YsqvMOetmNSZ/7D0Zt43ZdxeKDN1wD4xo8vRFn30VhxvwURhTzjSa5g71gPMcbW+sfNZR9FAcGJg
GhU2MfPMrEoKDoqyDwOUDyu3V9kUaJyjfiXLukRzicFyRTthtwh0vi7lBZFqFN7GGLZFA+fOiF4E
Q7H8UaWRo+rN4RCoa0wpEiY1W7ezscgBnX8nk6s7a2y4l60KnXU3z7ojJ1QGROOdujNkriCb/fhp
e9Ytrk5DQfSMjW2Qum2UzRVFFYQQU18ynrFtRHvaasHj4YOgJL77d1TLCOAZwPQkRaWwZ3XHWu/g
WWFXzpOvMFqGZWHt+1JpScuXgRWWDbMOiF0jijkcO8ksAE3HL1TPrDstPWqg42pkadop0SIR3ieP
/8e6nzqUj6wG/Rb3h2boR3SLWYU+AAKDZ8NgLeaQGGoy4rHLjkCsnRn7uXR1GQOwHqoUZCnqvTzJ
R+9hG47bpw48MfQOwngZJYW9x/HBYZHpkUU/QnefG1YiYs3IMz44ZPCuzyGPxVKGTtHQ7Ybum0S4
SfJakMjDSTkDenVFEFHu+3fLx/8otPJJifOOHyYMCR9bpFsjVN9VAlaAQvFqktRZZCMdFF6TKxyt
jv8I9/I2uwxXXB3eXTd4l6Nfke17/UBMYVJu2645MfGlUpnCyGP2Z+8zvhH/hPaPv0s7xWStVQM7
5vlkLffO+Zj+L11gV1uMnYfSF3wo8qe5EAbaUyx8HhZabe+h3fQTeSMKshsCbNyVAHRL/IoEP96F
38hU0cN+acCYyL8r2UOblQuSES/qbgX8QIwmZifgjpq/asx0kyBcMOTgW++kUAfOrvKd/lD79g+L
yxGtmkgaa17JQjuKRCjmvPC18Qsskox9gvaeLWYBvq3iNJvf4QJtkbd4eAzw5+LrfiYoAwzpkkRy
8QvCjNidnq0XebOY/QcYVX78Vxk2nvXiIJDs3iH4wGQhMWTjEwqqG1Se3wv8dJ510NP8V3Rrexp7
iY/8PMK0Dz5wPZnmJ1FqvmLhMffIo3Ws8C1at00Cx4NVR9UOd9GM7PPaGAvJYaw+Zl4SZOLnouBT
KP6vAgwVxmhvCT5N1ICTXPErfTgQFDd7btee9RaL5frIuinmIw5KQH3Jb4HmfFfsdXIpNO9we9S7
QlG06Y4DnlZ0HHpAo7gNr8vTEKn7fj6j0JTNqmiFp3+pErU9EsOwIHsSsP0bkNw3GrpCERGXUE/r
+XfYZotFDuHnVq6w70zR9hmCUaw3099otGva81k8VIYD6yEuBMFhrCUvMwJjuFSJmJlYniNmY0wz
AaVo+ASozh0qNhqlB6ETBY1WMm9+wpIJe3fqV3dMqzohFBLCWV5kicBCTHZX2WOX0mFShAdvWDG5
9o7D4iXgXpiLTlMMBxh2Rgv/quft4rzop9g/Vz0W9XI8zyKfmfqu0W1Mzx/URr3dT3rLzFA1bbWv
Poll+Rre3ktR5t28S/cOfxEVn7fkqQA+ZtuTkKPkJOx3XtE80CJT0FeJaDXzNG5oNMht++gsFi+k
BG6z/A/hbGrLO5QplaMkGnGdCuOxKVSUt9L3lXKgMcX6TFgJUmaMw6xtFzvWi4gJmEUdT2OGgTte
b/PitZqylqqp7GdUqDGTyA/ugtvQAOFbShW6UTwApr1kJ7Kyy8Is6kuFK1DczQ/NRNLh3EJ8ecL9
a4AYrCnuYXxgsUemxJ042/K1Ztuag5kPdwZYjw53OyDRs4SFyF3HI43UlHo8+DBhQb0+V+JetNO2
0MCSrq2ketbWtKgCDXM0F+lXozL/xOzAx3DdrKLrSVA1Xa+HhP0mpSoyfqnYkTiNbEZbA1uKX/XH
KbwuiYqc/ZYtrt8jkqyUSNK5+78pqBTmpOwBHW0+zm+LWQ3aq0uB9dCpOMvssUZaSsuta+Z8XZ+9
xn37qErwvWKvDYqbBr0FKcu/YGfLrxxHS0LcLfR9qL9f26jvb45GcwQ86jnf4fzkq++UH7yi6h4Z
86jZwTK/SNJ4k+VCXndWeoRVQyLK0Jj3zWt7jNXh6csWX8oWHQfj43Px/AU09JEZ5hXOgkq3WQ8F
Hc10jX3+5QVMYXE6adUHybdIxtz9rJSp5MyRjk7oufv9R4F2iuf/y74OTiGCsIzoTStAo9dZn1b6
Nxj2sIz8toonYt0EmXtp/2W29oPaat90DRmGwhJfjNxhYG2SgNwY2lKLnjNqWpYZeiYpGcjLGnO5
rmrXt7vqPxRtuoBJs6vBsudYQaoYMOw2GoqVKpcJZAaQXNrHChSKDca36L82oWYRM5ATC28H+0vt
1QPUedbqgGbZpndTg1O3JdhtM9BPrVHdhp5JbvmyYsckahFBZM6PBYdqo6u+z1zxNAp5NEx3r+CW
weu2Aa6HeHacIeBzQDXSCgTZiIZ4I9mRrwrXyuuXvPv0p3aUD+qOV2fl7mkYnTXYDCr+EQQNpYpy
hQy/IUi2Wwo1aN1zSlt18s3KcP8HGW4O8NKodc/em8d3BmmTE5csmbBMQd4j/eRlVJj8QZgMyhEK
8drudnDSq6dzM6lOb6FZc54SQcnE9WkioGKNGYOVttGLWagv1nV/apfJoA3+Naz46/9N7KWr4fbx
iXrciGFB/Nt92nSjEpNTNT4eisXB2CAY9F0ow7qt4DibtcuWPXMLgYKT50aTnyafqWj4NMqgsLe9
4FmNzd91vly9XYeKkpviqrSNdDYU3zAEOXdQfjaZPIYh0zZo3YjqC95X+cfiYFrbXWo+mI63AOZO
5aye3DE53UwziZzUGGRys27UllGl6JAcCKGzbysx64NdBvK8Q1H6n9LSBvWye/FVxVkv3aCgh+3t
qpZiigq8hOgFtTDsUECeo4MC9iMyq7mHwxAMju8b5rJy9BDYE0Nx3D4jpO6Y48KVz3/T/c6HdjJJ
Eux5DOdElFB3d4UsGnm8Rytij5PdL4JETUb/+w1/ziQrrVSDtX1rhnls1aGR2cfSPK5h0v1pZ7Ak
opsrLmjy2o12Kj+ioJLXr5AP7u6PZ3HyfKQzQKjAjms8G4TZfeEOYnx9NPbfLUDp8r65wuUy00xb
HmU969VkKNRm5iSVMCAYOLxKD2ont4J3bB7XMB8Z+Y3X2vwHQO9xEKQ+3zn7uaWJ3qnFZGyHazOH
WJ3XReGb5w8qPeUgOle15hUh2jzEyQC1DZUHoCSBFhTYOJXrgMJkpdjpHBEi2DUY8EqxHQIiaAF0
80s6+/+UsUHlsd+9psk4cM6p0NvaiPRzoVYi9A5W6IOneue4cB+PZqyN0tAyolOMHvgb7krzph4I
3AsX2c5pcO0r0cYhKgm0izHXLQD5s/1iHm7ZlKEqW/6aWm40/f4HjVzNF0yihHL8EO6nl5rrkP9h
+A8mUdSFvICfxDiMOCh7/WyZeULVeVAz/2wJdMC4f9Kzrch+ym4ViRZWXdCwAhal6TN/sHNKxwwD
M17Zs4m7qvXLdaMkudn4P5EHHuUKOW7kJUkqqqvMgRvVpaq7YrldimZ5+bXUfrG1jzGFXTxi4D5N
KnOyx9wAWLhJTcPZPG5cpTHe25toCBlztHguIp0P8+QjRRu9VgiGczwvr/cMkwFWB3d8fA5d1zSu
lJB3gznNwCmRxETXp60Zw2pwcAUsbqSM0XT6hHNtaKMYCOjBvz091WHhXWj4SMxmWiPLLUkqBHcm
QjV9SkB53bF5VywbB1RmH+MqCgIdIsx3cgg2vzAzLR0VCIt59wuePAHlrraXJw0yskKr3TmRBMZj
TkWa62ETpfk9OLlddQUi4ZBRKJl/wzFXQS0Egxji8Ze7D6kEhYjQz1Bxg4rNVNpZOSq5YnHQE89q
GoID3IWiqKGZk7CziL58GoqrdmKfVUtKyzLk9hwW+IlprBOJHlfEkQy2WIFVNAzpes9ObsU/zMTU
z5Yg2bGcU4JQnwTbMTLTWtPCMWpyxv673+wxbFzKQpD+fyFI/gYPRD7KSLhu0ILj5KDmav3//zC5
u/ZaTNVqpUed5P+qwg5On0vHrTqtk1p4vwntR32JZwuKSA2vCLNflOMgI7Xua5uLPPxiavODBOwn
z5yZr5Y9U3DHXLrAyIXiSU0jymIO+Rqx/HCNLXl/2KYlLfekMPcaryU/LvI7+K4iGrNxLosg31cJ
l7UsG+2yGav9xw0oBU8jU4KesBvFXCdiV0Q9aDMzyaZmnCXbnS7Xsl/8i1DZjwFpsEwKRP1Fcwxb
j99Kab2AQf9jIPFkiIMRfEm5Ot2AW4Ulhfs0gL2Z8ZPFqliZ16kNs9K09lgylNn53zwtwU0RMmEk
CommnAzJ89HS/G/AELzHggU6QtDV6YZ1nbS24gH7FIEGQW6dt48l74Hlt34ag8ebjOl1j6/gkXnm
0J2oLU+E8z6YWyuseV1kWAIxW8/5ceFg31STaRz19Q64pz8BGVzUV16K8QaU1AicclnqNOgFh2HL
xJPu+IkCYSf3WHUBbHCCCJsOsV+xQm0ypXOKxaLcrNlfRmzfoE1YQsKy0+BTzt0JdoRnP3apGaMg
hsnmH1IU3sTTHD9R/Ap1+/9sLLic+Sb4oDJmWsL1JFq1AU1aWCZtWYsBhuLK4m1WryDqPwYEkMQN
+7c3jn+qX3F7qzD/fuLlClBLxpr1KH5lVD4imtA3SnX0TpW/ZlTJEKpvahnWaFBfUnqxl0m90axa
1qGOzyN6xxsbb76DairBGuAAI2L1iqTEzOWRlnP2zuDFElp9CBItdsLPLi589NG4B4v6NNsLsg1G
uF6fD5jC/G433rj+2nlzst2pBGuK7vhnA0Yr0puuWVgJ4yw42yoXOSiKMFifOvitGRov5ocJLPoO
Evd3Agn9TOZ1qNu69scnha38TObRSU1ylnXO5isj/ghUBZoZot557xuRDfAryxM2CfPa4Apxntq9
PRXFOQ2NKqtrLnp1gG+BjBJtvavLaXiUpeCRTJi2Q9PAmGgneVHWRV+Y/KkvMtVsSTNNRsX8sH7W
tZ4AUoT7UUlwmnvXADXBDTox81Q14wouM5uABEAu4+ETooRv8iMOaZbDN7XdnUIHjyTfr6tLda87
ZV48tvh3HGmQjrRH5s32sXS99y2OQrIARirjTNFzJ5ewZOEehPJCv4UnHtZrgkkZIXIUsXmfHipz
sbXEdYUlKoTOPIihXswJMDAKSMJpX2BLqaq6GFfpLZv1poDX+M+oSlmDA2dNXAjwm6rTdajoarzk
Xqm8wccIKs1s+JMgwiQRz3DhRrQoYMxeN1rvvZ0L7LskS5QQPSoE71eSl9wmjvXIDtbDeryLrYBx
CNdHw2NTVl8fKxPYmFuD2cL2Wa97fzDfFGaO/Z/oKr5gW0CIqxE9rrE1YfZniX/6YPLWD4LqK128
eQO8wLCMIX02mgWzQQtHOSJxkTwyVmGhEPLBuzBELJcMmJI66dmc6lHP+boFw/2J3dvYKpjwdsyv
Ef1S2Zbu/jLcNiBMwumnX6tSEodtT6ah1Zsqp+dzllVBjcj9y4yJTSigvmD+ojK5dTrnQRxudtKe
sNNWN/UQSJ6/6Rc94PJbsW5OguRK307wyhEmExmhv1KN1DO414p4Iy6tuJ1mN9DotCpWtTd0IzNa
JPdFPOokMeeibiaRh8hycRCUFoh1x33EpZo72zWoj43cPn63LLUkH0UjV7YG4gZ7ZbThij6lmk0X
13L1+2D6EwTMKGLBR/xNyQqJUj+Oef1SLmNNV3ysnGjA3VSlbrz6y3wdLI8KT96EimZOqjPm6xmA
X4eFU0521KFPlMSjDOf48AhUd14F6wBUxrFPDg360S5wxuvU4VdHyxJGrEKMR99PJhccLDuHHaKs
90AOuF29oV/+WyXVLLeGNDrvyewlwC5sPQVXCKt3SvkKRB9EXTZTT55X/Cvfn3Wmof9YHiH4T3GZ
sxut5zjF/BFb9Eyw77zG+E9/0khMfOIr8/1AY88pC0OSDteX1pN4inJVNDjv4cMzm/PoivcgR8tk
lJQnIIGaNB1vHfPEHhn42hfx4ye65W2B+rlZI0Wqd9AZh1F2nxrIZzUCqEiUd5IgD4vW3rIXj8R0
DOY4CTpDK+8MsPo+hh4vEQIeITJtxXPWr8eVeEInh3k/8/Iii83jD4vQ8sbxlYJUw2s1ulJzilB7
JW2TBPgFbFMxSZztfT2EF9qcDdwCrpvxE4S7GRVOyn03+s9Cnp25DazSCH4jdKRvd08Y0IO0FFvt
Vz0aXVTYEOPLFKfwmSXgH3oIH842lummkOHkVtPm+yuytwYcsvY6qryatKJm/oFUHAWeP83fTxvv
nNmUS+bZQjzeJVN52DvbDT8DrL6Lq8WbWv/BMsIydcUewFTzOhqnzkMi09OyTE5TDKIUZczU+TYC
kForTgt5R6j/R+j5dZs0eU4cAlpqcBtLC1OM+qnlM2dzEhfsU0aeVMJleYhG5EiyYRc3rz5NYgsM
m/G3CJx/Pa8KWNHi/bNoPxMThb5TRwXCnMXzOUHNUgjyBOIUXBNahedsOlkmHOqE8ajDYZkMWmHP
urh+Xc+AJ+FoMLL3wVF4r/RPQfKLH0FrYyNjQSyIIYguYk5oioSkduN07WMBTT3uo0dUt1xrLEEL
gzTEYd0oBpXyJVdXhs2Zomfb5FBMI+wViOCfkrg70KA6DxtHcrqqhuQLxz01Ysn4yFUQcsuV0ZSJ
Ey1oWpDUqsmraN36pWXRCawDnEpsgaXtGUmCbFfzkC8ChptT2UgfOLNXD5TEhZP8JVzK+kKqVYJ8
Cb4MR01y2Tw47vNNToo/04RZ7HkuzpfxnD5Wb8+RJW/LaEiEbwV5qdPH0x08vtABvQXmT2gCL6SN
EWtDhf9wehqUv2CgXYH+k4t5pdkGl7yjpjtEv+nuyNpxRWm4+RuhrIPn6TKV63DExQB3Yxu7Bja/
elTSL3YFnLYvj7ZkMGqVuUhUfy3hWKNhqdp+gMcghKmjhERfa5+wvYOXnrXa2lI7b6avE2qGaN1L
zwIOWAstEHuJzFParVQ3C8R6OoPh3ykr3XAcgL//UYgGQ4iGJSl1RQRqeGsPYXlONPxsOtK7XsAF
bGG0P+OX+V70heQjI5yhR7v7b2vKpllvsdp2/e1wwes81U2LPWrBn1PSctDEMhyyVODdNR5TkXxY
fITubTVkM4pNTbTzJKLS/SiBtEQG7QUR0MsYwOId65JxwQ3h0y2h6pYLv3gFFH4HN3QgnmDqNnpb
j7ICrEE8gREgFEDQZvg2XYVU2C0xeDUYuZT79E3imnSEdtZolmyQFGu8Rr9HvxDEQ/w0OCL0uq7s
zWIjHeONuHeFQ5NQ8WsDRY4mGOerZe4jFXDUOH+c4n8iKnr2XdSd87X2zl+AX9lOoWps2QcQL1YC
O895QekuyWI7dIdA1vgJ/43ff503Nrv9gjB48uCbk1ZnDwO7MeSnQrOEWMSvK2vTwWVoz8Pv02QQ
LVkHgVplTL8XeO+utZ8FIhzwpjI7tMhTfXQcx05WO8eU1aqvA7PdAkH56L5SPQ2RIu182HFaZJIz
AvSvI0cld4qtqo6oJ8Ui+Qx4Ca2DOLuR5sq0ZxGnpJhGnA8xkdE2Bsdwwzk1Qqerbk6IVoh4/JD+
sKx1q7bQda5Gt+HWZr6oI+Vol9+St+DxKHlAzj89OM9w10sVD1hxWCW4MHu9w26OLPg7PYsJn5Yy
o2+x2Y0OE8AsOPR/hR3GlT3MUAAYIXnmkp6Uw4wSZzCYyTXl5YdPpw7GGJnnECYtlRIjLMEavN/T
EBhpAuK7OninkIT+/Y7MkSCsAOQLfK69hVLz0R0ytK6Ui6q0wWRGcQpoK28smdQ91bS6GndD6j4v
BaHNfU8E1t7Z/QlPJiBOKzyJv58S4zOqyFIE38VI9Cm9cgTae0ZghDfTiS7ZZ1Mxa4vtkRrHbZx+
3YCuzW1hWQHJk5ZEWGU1BiugfxHJfYwTI0PesiOJ2rewn9gUMkhTe6TzCaaOiAUaqkOLKNwucicL
LaFm84C9WP7TRKh7F0KHdeRd6w3aNXpV5+SmU79Nme/rV1pvSAS5UI2JyLt+LleNCFaUi39PvALM
b4NgjbAj2PBm0moeMeeyAvFFxozRZlkERvN3jfusqL5ouw8KejcHwLeNq6dw5kISsJvVqtxBj9nz
ff7A1EK7hmN5brLgWDRHBjRTI+jHlirKjuHFod+kBiyQrvKl6Z2t/+mnv5GaMant//03r6MGonOo
MqKio+vIesqXySG7zYtPNRYDNVrQxTKGeXXw6/uyPktBqiJZGHVFqBcQzwYV/+YaZ63HAitMT75f
mAqJG4z0CgtWPkosvT3agR4NInzBYi0c8RbjGdlXHGppvLkrrNQK7S52ZJkomgLm9bByIpGZXc3J
FkbFxnHZWHC7oK5tmJ8FooYDvzXvbIxEC/3+u93K3iJ2hcAdcKdfp42CsQqKlzCRKlHaoHHJPJmF
C98RLZggKwUoptGL3wBC3L0NgiIDUo0KGetd/duBY+gN1ftaQKmgdG7cmycLdY0EWqTmZH5OrD/W
AvMBuzuSHtZ3BUc6tqlowNrgEMGZQr2BLWaqJFrkkq7o27vEvOVS8a1Ts5l7ZiEniA9HbdZDEtn9
3fpgMCDnKsK56x4IQI3UEZARQyo474dUP3TvYtnEaGBTwn9tkDpayXmVVzx1t78SkKZ1Ma/K+PJY
QRcgyAzqax5oNDPgErft8nXi/CwhMyK1nR2W3eNquFY0ohvYuNuvYZ2f5v2fkinOrG8Y/Dji6jAk
zJGrTteVuvEfsFlGXKVJsFi1l2FAzDXXHNmwytj69fu6NC/ejCsMbOwWRPq+5sJAbVoYqdWeJpHG
SiYB1ANWuVktkUNU81rL3smMUbUAVb4KtuXP1O0rkdAfYh8WdyFZzdGc+jNQcUaVnoi6Z6Nqlra4
8mX4qJzZpfboWmZAaj1KR4tv1wMD9KXsdN7YoRbVtespILmdGdN2xCxYu6SmJq1HadVbzD7fWhMX
0uX4+mnYuYS+cqWwL1VrJnLTpr6BSjCVbwAjDr+vG/mDh7CVmc9aJpWJuTmKmHfK+BF/FLsaXR0n
YboEiiTWd1dPnmGNIPR9v06ygT1OqqeatvffJXaP6Vd58qYtVNh9x3f3Z7ButMPlO+gt3Y4kX4U6
wX4RlshYxplI0rbSoxJegL4kZcYmKtrBWhdzppIf5dCy980es7OqbXk1A6fLzyGejH+EgKf/SmsC
sB/lB5ADzolgDfzi90yILYAjGWhSPqy7VW0CIOupJni5BFQ2yoxGPiLG2eoGx3LH8KUQ59jPIvff
CF3rQuL3cnuD1zUIIa5GJAmbQvRY8Md1dHyf9YBy8+nngEhUHXtU2cnAj8qhAN9C7sSRRV/NPt8s
fkUpDpSWPXDQ99pNFMbDwC9pKZUb84CoxVHqbOzF0to3frSTZYXNT7sUHt3JSctzhtce2ZH4xYTT
Vruk+ZjL1uAds+LTY4RUFp4C/x7LWQ50Hh2euT+KpaOIxkfXHaqLaVUM4y90uFCqyxaJcqvEe5JJ
do1iWgDJb7DU/5qWhv4uehOcetEdcRnR/lpaJifzskothHEjoPDIAZbVsmJcvRt+IgClhKPkdKdf
VSdQIQvZ5B2F8FqE4oJQivusWFhUWsr0CbmIfXZq/kb59DwVg1C7mxhXKfKUtGtTVxoJgFrN2xHE
nrDJQhnYxO6Io6cbbcuBHzMDxcf75F/+4gqt8OMNqofqBXS1v8cUuA25hNNf6cxHMCdjvqYV08am
+Yqp9KAl1bnF/usXJQp1srMuuPW4iw5GrdqIFHDbAacliiDrPoUx4bjJddLCf1IPPXSp+xWvGZhv
7Oz2Qeucbo5xLTbTCctJeE9hqTlvD2hbmUGok4tPJfpxzlg657GKGSqprSNUTarKGA/QswkFWbCq
ujQly50jfZ1Ay/SAgm+7y646yRtz5LLzfoRo37/VEE21Mcuuaf+oh59tOaXZgUctk4bsiCcH1QsW
4TIQh+uV4VGv9BcH01LmZx1ovYq5EDrw1DY/T3LO5mIorUlglEh+0PD+7+Z4Y3atI2xSY8WUcRlS
NALuJBrK2DiWHHk9IFYYPSx9S2ONBoqE3JptvmWKoRm+D9SRFiK/6bKwzC8iZWbXSy6gdJiuk1SU
z0BupOz81tcdEeiguj/qelnl+rTIRpKOni+aEZn1dmvblKRl1v/UBzkiH1f4pCqJrFH4JU0c+SCp
z7fMENlSMWrw4+uMPMBVi8LN7lMjRLUXvTjWS0Xli701mhMgSBOMeDyBF3vB0mwzhkSvm4MjdlPq
pNY8uCgSrc6WZGVYzXxR7Bz2An+QS6guR+piN7R55oNCgiQyVkf2Q3VAt8TwB+eqb7B2DUX1KDLM
AEl/MIhw+xVVhhjVB3K2Q0jYG++oA2edUZrybJflND7XSW7RV9JBrfpzc85mrzJwkssoB+Nf3v0l
LAzK1ZLtCa1+rlJLCVuV5kRAF+e4E7p5Sw86td6CLN4hAMarU4cfmwEGOCi3VGkKy3A+WxVBHIps
1I3euWYc9l3473wZI0t+ep6pRej5hMb3Q01rP31C/akaeuL3Q4HPqp03S1IbcawZwBjRvJiwueCG
Fa5wpbXU83OuSUqwxPtfkYPxJBpuIZ3bsBP37XGZ6b9u5g7y925NWTd8GakydeT9snUyHpyZCcM6
I7ECTtTmJV1uqJhP2SnryPiFtGj9yLN+ctLtd5CGLZhBq6tgpPraNKMcBWoY5kBMiPsN5A4oPEY/
B6KMgXcIq7KLjs9Ea0g0q+5w3vmXdC5ZRfWVringM+y447JCFkhphlOVc0VCTxqaOjuu7RUaLm6Q
VnTdWICc4E8+jmjpUJVt7Ow7ZOBCNz9BRohNtJ7aAa8Yb83+dUpRV4GCGDhYvU0ICFQJEb1jecyn
qphCw54+YWQLagjbYkZFJXryRsa8z+Z3ukyy5H+duMwysdVSIcRA/r+IFenoMgeOBzRlUfGDFAmm
l4HV5i5g3ljMNExAeoFlil3LTF1N7eY1bB894JGrE/Q+eyMj66Ztdo+v3g/SMddHdwEhwdYdsb8x
2buKgWtdvKoU1nah2/Edcn445D464IoEayBRP3NLz33DT7GXkWyc9alrShpd80hk0HGGa/ZWvq+R
gBqnTcamBC3kmXzjnjep8CKK9pDINn3IbWQR+0zbuSNW/VleSMIkhFmgNxXnX/nfRigvKO3cRxnb
+ecadv7T+BFK/Nb1tuydg/xmlbjUSS1yUiw/p78PsrZVf68VhZsFbrMmmkpINZLQzOSE7BSSvaFj
JFijvrtlctftL+edAS4TN8uC1OLx/l2vHCScVmOP5sd9pHNzy4drmhQVBpHm1vnQSWFXNTYWtGeH
jL6F/iHl2IXxvO2KV7OpikNCHN4Zu+CMyfpJ7oUQQAaY3GOnwHCm/a9/CUH/c+DdPS+Vvp1Pjwbl
Ms4qqDymt+3KmTk0G45Mr420jRqIwGwFZ3cPRNuzIBGab4vBzaDW/5DNlec/HaVG2guVTcSlL4dw
jksQGd8ucKUm5VJyDslYWjF9r4ewNSIKMp7eccJSFdLLGEVT7CU4o8R7L3UHtjLiF0qdf0XcUOCF
YVlFDFCiETJWPtaVTFtO6AHauKnML/hg9zmUi3lfW6M8fVnpuQGYMCIAtiLGuYZcaVgC1V4gbXYA
VHf2SLs6Of64NqUX8Q/Ld4IIrQQ9zXso/+Yq2m2wC4ma6ZhfgvwRr30jYz6rZWbpwISsU9pXpfrw
ZOX3G9O4K4wVT5g88lroVrhwamkbj1FfyLo2Z8lF4L5hBAl/Ix2/Ps0QakHYBw27QyZ7qRTz4hHE
q7tJMdDJSJyyMv1iGOJH71gGWHABk9I67WOUT9jxFJ0JET2ISLDCPYagmi1W7HYkX062nG9URpl3
WuLUEI2nGWXfUQjvDoxcX+hmCCGkOmS8Wqe/cgGlGDGtSK3kOUhI5KEwUlawAYog8vRShV63MsXC
VfIP6AngB4sndDwaoLTrh4e2u5Bxh+uxfqc7LvjcV43HXlNdbACr0qO7Lsdxty6PtZu3U/A7947a
IirM6uQ0NqX90Yotw9hiEVuqj1MInY9fe7uZUdCWko9SEkrK+pb5KS9Hruava1SzjLdsHuNZIvnU
JK2yRoKyk9xtUuDlTtkbq6uzW3CAslQtk5VYqGtxyMGbQJUMSseBF+NqiM0F5zevpqXuFFAB8cGb
OTaDNDsJkNvvyVCaqOpxxQ6PwZMS6VRcR0UIvBDQ6JsYnvMXk3dHlzOW9pQmGNel9hxQ8OX/7q0s
Tp+Ra3DY+/Tz/jRmLo6hEk7wdW8lHnrhOBV8Th9muW2qWHXFv3gUroeLadXkVA6bwCuEshWIqFuP
CAJfjG9U4XfUc2YTad50ntnEoJOUtptHXCT3OK9E+42Kftc3jdnd5Q+y0P14nwqGYUzI4rJm8ibD
dIYq509CnD9GyoWiIXruOSHSHuDy0dvu9zMqsx+Fim/DRYQvNayhmrzrKFOIOvN8+4GyROUOkddp
9tK4jbcNySeLb8isKVnVvOMHzE0UVPl0INgJVbkV7G2bfsTNIb7G5viklFUG1PIW28L7yDjpNwpq
3AXITL5BEW/oQa/5BVp55JGV7ExH2yQyhWdh/oLf/6kbpxOhpRFjLDvePQCDyXXZqnTjyTZ3o6j6
dWj73W7LXvljTpt9q0dwuK15VWdZwdAqwC7SYQTBeSggJtESgu13No/y43L+MhZGyk8CDenUFZgB
t432phDbN1qpx2teVvWQhCEJcuHQpJn44xZHZPXdyiajWGxqAoIuE2ziGvKtYnI3oegD4WbUaRtx
vBouoi9fPIjX42lnxZCEFO7lhwOvuC+UDpVYezgo/JmBL3YXqQNRlZjti9Q4Bh+Qd2BR4mR2jrIg
DqeakDStRV/umx4uJp2JUoSO0y261iI989NcGeXWkgN+DzMpNKD9QDXL6DAPxdOd8hfO6G+lQYiT
g8CXZqvozzbNQeVb0zVEXwMROTDnsx4GOQJD7WRcS2qvpSIoqBY8mv/sp5vh9aI+/KtciDcxsj7/
Rlen1VDNPbBoFG5X4TxsGDZEsFZfBPyv1IyEbrirxLwU0P3PcxE142btBFcT840bkiWasLuTnkB4
AS0FXg0Hn9lPNE8WMhHL9JCC0biwb2evO6onCdQwmGcVLC7MxJ1NglyV3UcLHpPT+uPegJLx+URK
s13lDb2qdHHOsqgIywPLICx9tVRdSo2ffEkgJ2XMHtZx7QKhxakVIJdDUiPKaLo4C4xBiVsN5z38
r2tQeLaRXpdEatzQN1Fl3kENyqdPiuIsfdvys86FB2KpwQ/VH5/vkn0ki1s1l/hGUDeNthSSvjPo
FO5i9ZOnNowSkUZzrNYW1L+U6x6fk1xswZUlrSSVG4Oy6FilMOMS6FfrHT6u3rw1aWSUIvESPe7p
zQsX2Crxx5WdI2+B9ibSxjIG450dyV+GeHEjpsi5yKdHYOGda6oMli+Y7UNKN7ebNKCoGwQ3M3ic
Bi40yJqauIrZ5aG77br9yx8NAbLD5EL12tsWZ9ZOiSbwHva+B5Y3TcU57hb6xeyndHT3mpNen6dA
ix07TdFp38vwgoEsXdkfDjB/cMJQpY/GnLZJwOSMJVJSXtqhgOvUDm/NpOwmZw3q+UYnaqAGcWf2
b30XxockwGu2ejtYfWd1GyVEuLzr9OlPmOBGLUhbSTI5fwdn/FNZsd1XDu04/CZROt9jAjUu+RpV
MZpm1/V6yTY72GjwuFiNxBNmLW0HWv0jYV5iMo6xJAu/AMPWbZ11BbBAHHJlqnQyOTujMcICvZXr
P8Ih/vkprH9p8zEj279U7vcUUnaK6BZeSOuY5/sNgxe1BDgZwn1h1mJVQuJwZr0AUN4rIZX7T//X
/XeHfEnJCoft4Tc6tZj4npJWxx0n85G0xA/zhmW3vHobsJZmRSjWjQHeq80uxSb29EVKrTD8rMcO
OWtkia/GG/GhuO68tVNTEH+ZxFDJXK8cO19CLuQItlN+tHkmz65pk5LIxB5G97H2RruhZZhDWLx8
BQZnRgbQMbsNZXbICGtbXln3ZELbGn3E/1p15nHuXt0+s2BStuaNIdEiMSkY5lDv6wx5OOnGPkar
a3tn61pw5uxn3nS0OUcKzCXc9EDMY61KEnEGo29QybFY+TJUcKiN6bFncrKutZtCzmU7JYS3x7Ko
Yo6eZk10qrCOI46oGm2SMjF+iKl1/PjmVaLgz6cayedj3AOl3vQ3/FJDZJivsNt6ye1IUrTL9T3w
fgYEtA53eqyeATi71ew9Uf06O6qekvDgKZDjHKQpw6YyDFTWQnHQ/kvFxtlg2vTMdHWh2rVSarea
cf265iEnN7IkVepocP+eXRl7eSpBPsaZYTHFp5WiycIBASUrnoG8ver/z2GJ2pFQtQOSvyULyR5R
ZJlfBjhSi/TH24YGmsRZ/cx0eFNV2gu7ANJtDXp64Hdo+cEc7r0y7VWnQSzTibFUqJZMCqdQKGzL
+1gub9ata+MPyyQffR1HQFlZi1PVmL/4LQYaWHiGz4d3eCZIlq0n9AG7O7233UsHQCTeX9VTlc1K
oKHootA+VqdJQaO0avKU9//9JQWiqWYRFJ6aeBiHQmHCTEmYpEFiQgc4PIA1hEl3rMD6V3Cr7p6c
WIsg6xvPVpE2Y5qeqvApX+hfstmoYDINMITjk+BCUpawymVlWobZNoLhbNvI+qVxkSquoIgwAmU7
yCyU13METJn0VCdyO5Zhu+1lD5FSWzmW5yjId2/3vBZlcx9tx0Q7aTlwScNOnpvUB3KnjkAchu9I
2BUVLZSrhmtDh/A3dUPSdTf3TypN6AIiBZQg5cW32NpY0z9TCgdX14ohVWgbj5ejER5hqMUWzXY8
L4GdlkEtuYNcQW1XpQPEy6/BLQdCdNAie+U9FPIBxAaGGfjcy2jqsg1JXHMQUI7W4b25LwCUalNA
vT9wWr4SPQYfnCCQJzfenS2FTXodV9ZtJ+V1YPC25Qd4Xz3b1A8D5Yue8lzLoPW9K1UJzIKlIYg+
DxRzoZ0Bs84vqR2VbggEGAlFHJs54nI0naiDI6YdJ6O/lECE5mvrqJBvDXmfZBGs1AmH1rnq+Bwb
MjbUYD04LYNNQwJpAAW7HCg3doHI14yJzjPdo3mN+q4FsRefGbNUkqNsvZGSYzqQpfTnjn4P5qbk
b0lNeBJTPsC8IaTTcpFE7kFXpTx8vrReCyqfSMm9RQ6AKTEibnTaSmxQ6DzQcJBn60XAV9ALbhkp
okOSQDhn0FNErc8z7nHL3LwJ4ivFYLMfClafyHhRGG+Ma57DlLa2snipDPMxww0iy6eIfU8EgU2e
9hM2iTpzMesqlf7e3uXdCfbeWxCfWPysk64DfyVpc5tR0OcOKL8ozQtUMwY7YiORDgNI9IPfN+kD
8XuqoHvIQHOCiaEm3v+XcAt3dCEbInQNke4rse/ITdC1IcA3DmjQhYzTemS8xi/UulAJ7gndoMxu
4byPd5i96G17eai8B6Q5z1sSFJv0Sqc3B1LTEv4jqH7hml8AQtmvAU6SxLUw0UR/4Jvcq44qfMcC
wqdbX1vsiK7cD1ChWSVZH8LrUWjlkSETHEFpQ/2Cy3jOVLe7dEo4d2OPb8gudz+qtxwCu3CJ8rW4
eTP5hXgGOkgRskbA0kRuznzG2/IZNzuo+11CodBjS4L02Z86eQgxe7m0TWqMzZPqQ1OGPvdo9Wu3
pb/zPT9rHUpbnYUpgjOeD7ArWgQLRQfoAnhLae8/IedWstnTiLK2W8/mgd7jumSe0O68+WQDjLYL
XR9LNZ/orfyb2HePJ9GTft7+33rkFQIsPaH+13PUafxtGgzFNsWV16Ub83SOkSu0ncq4m9Rx6hsZ
OM8k5xspaD794URrD4v0LoILgiVfpdnRDCMSdx2YWHa76kMGQI8SKI8OaO7I26GvvFVsYy4spcXH
DZp7IVPG4CEADrXZUIBKpkywzNYv7IaXapVHiKMNjBZlI4fjWvWKo5hH3a18llCIbnksa5RXx6gI
uZnk1jz9OCeVJHnJsqHSvgcJsxA9N9xLsgxJ+rdfgAtOJglwRawDdPi5bdAKl4Iu+E3R1yIiR7V9
XFreIE6oaCIjvD64pUDwosSMHtEOV9i3cVrAnbzWqAEK2wy10pQ4J5fwrms9ytFGOjxzlzv+L/J1
THdz4sd+171dDOXzOEGBaXSGQShA1YczuSPQCobJNJiUFa+UD8c80CMkLXevUrrmKOXc9vkNamR4
vSfqzFZjadxeunPecZo7TqlkS9eIiGJyQcnr3yrBaqJb6mrROiARM7NCs1Tr0IByNVuZ3XNPRpAd
eKpqfCql2SaF24UR+Gva+saMdaNzQ36RoCjs0niFSCRL7B/VVyqO9Uh0QowIxAJHlVVboNyJoU22
tHV+LaHBCbVR2iD0qiJolhlYSEvrCCMA5TNear2u6M9rv4N1lD8Y3HMM5AgTC94FYaRF/3WWGCQa
ZWCd0SSoqefrZWgNlwGYP6VHjK97MTUJ+JVYRl/aKOzCLl9EU1GSyO0wt3vwvpdvlAHu41Gp1qAR
l2ImxQRhESfxiOQj1fNDh32APVGOBL7HS/2+VtIvxNzYadCXdP8TcsFkN/h0qTA4dE0D57gOkCfq
wOEEK/hsEbMUMkxMQBl+VXR1Yl8FVmw+n5VbYVL19WPGdJPguXxnewLrhAb1GKOMssF1Jz4vJH2K
t0cRK6gLjZcHQafftU7IIw4UgwRNl4AXMt41XokfpIt79qnbv9SpXu32HRLyL0cGOp/Rrur4KbFd
zx0Fvsj5iCfasptS9ZHU6u/fyFfpKAv1FKZ54XuY9DHtTMrtdrMUARYouumZ+J4KRFQ7O06Sm0ft
ffcK5HBsIGRO9a9X2sZ1HUDbXxbIMVRvp1A3Fdw6o7Jib9JKpqwRHgatBwGqJtZIiqKdEZa5132l
TCeeg5FzxirIgEx0y8DfmGYkJkeh7g7x9brdLHd/x0AAs3EgFfiR95tNfsUdX5iBxX30/+6jgRsf
/cN8CaRWuQgTWM6Zyxjfymi7tXrE7xGwsYXIM/ifCsVxUIAxsMlNMWT11AZZmW2FQlTEPfywFt3v
xA8hSUCnR7QG3AtQ9EEYX6QkyroRFjLgvjtJ8O7aCCTyaAMMPhie+tNBp+UoLYGdsP6clU/DNOXw
OQvxWjdVdaHtRrL5ObEA/g++b1YvQEfjbA4DlepA+XxIU7oC3Igblar6lkNOgl4rUKhqI4RP7RJh
aXq493XnJO9/sCHxGdwy0Za/dCfkdJY4m77BIxlH8KkinR9swTN/8YH82muAu2EbYODFL7se+kjS
KiK3LlTsz0ff28WxT8lsQAq5NMxVjHj05NypEer7NEyBBb47SEgQFgtsH4ZeK3AnqZ+u99x2bPIu
UW5JSaYP//i9lWeHqD2HeK42QY+vAVEzA60oL9DboKOh9YQoGXUED8Zh7Y2x7cJ47H9lIW4vbsY4
KSbDto1s+ujCPNGpWNsCZeq2neK2xRfGt4lxhSh2LbwMhm7yv2AWK/igsF132R4WEG75yfpUh7wv
ozKn8dLzDnBQCqHUYau3f1XrCHFEEjZ08ETnf0/DJyuYL3OVjiR17nL5gjTY4laBxRlgFhwl+N+N
Mykh7DlilPxUJxdNkfGf8nakM/9D7R6UmEE//sbfvJdKN7URvgn8DF5jwoowxaa9xyT1DaOLOHa7
0aGgyzaEsPopZkV+b4ElOlkcCWHxaN7cETpO5jBdcWG7E88KHZozVvP6SuSSQ73oFhdv64Se/mcX
ZGN8ROHejSnBY3TaMcdC8YPwpQW6Q1gcywtRBwjDDAy3HJPoSc2IsCXsWHvzIEfaQq4lm0ftDoFu
0v78vNGSXZ6ScKOMocB1hA2xym/rhRh39al8DS7ukjMnSUiNw7SMn0OOXs/2YC2kwVNYEAqGEwbP
JLPB0UM3MS1M/ERERC3211VsDN6GTTQuAl3PJnnQ09sisxbVFVB4EgZi7nd64LM/Ik6RAsz/RbjN
hNKfXzO+5T6YjIJZeKhXbTZebHSknBNV12dzBPbaq8mQ1ogNYGcvcjzWBEszC/ytJEDdutyL4GZK
ikZE+5IlYe2wcnhtc28doNIAZ8yfmrjanV7TSXPmKPUmNppoDyV4/YNNq1ZNyftA0LXEMY1S4Rbx
b4PxleM4VYTr20jQfD/3p56WyfoRqlca6xFDCwJUX4lWt05xBPERzoOLNvLMMAQPi6tdgbibIQVJ
xKTj8r6cTaYNsmJT6YThFmraetRO/wM8lKu/xM348b3nvwXb/bdXGEhhyK+4ojy96gxDGGSaCFyy
5fWXzRwUEFqiQwvKRZgo/Jeh5FPjtnheQIH7+d/S0tIoJOwGIMN5u0y4WX8l/58SfapPd96S1V0g
6Dj6wRcKLYRoLWjhy1xXL29yG647FemHL75kldx49kz2uwrLepwXdAbAQ0Jf8+t0MbxrzbPma/53
8zQQCF0X3QpuYRKdhMIjh0ygrL6c35jvgc9wJPsJAfa0er9xpqMua6obf2LPkiWWxUvojYlLZdyc
n90lk2mBQjFOWhCQBMQY3fZT2d7uPMCrk+j0XGGVD9qOke5RhD2Vr37XRSbxrgSeRx7ASL206v+8
E4Q51NTGrLc3k6xrVBGaB4I9agTFPXDJHelakw6U7dabQbZTYxW2VA63puYPweQdhE2Fk9Qwz+7s
FMH7WtC0jmmbHqoeV9thjGpaHnpulujmBBDbn3HzTNctTakOIENOUhNX7yBGNkuwK26VKtSPFgge
74foW10ANrsyStURyxxpRPll5GVb0GG6Y4N1AVJFCDiePdqdQbBtaxWk5P1MQ3dPFc58innwhN+q
gT1HdKflXGxQXySwKAntHDcNjyFwK3L3xwNfRaNQyMyuC62WfN9/T0/ieACKbgKYgKi5hwfzcRCq
SXLWqd3VjbypK3zaobk9qf45YzesOH/G9+Yi4Cb3+cWHFLvzSiaRRSMNvbmt/443inhnjcbGgGqE
ivjV22mOqfut7G1xH66CaPt6vo7zT3RLe5AntKmO9cfPwCNfApSeBPm8mBmSrqEoeWN37j+Cn0mg
vuq8TC6N5hro71hx9Jzaa/YW/omvFm5Q8hxJ8UgPol1egjfXqcHoOu86plcf6uEAhPb22a2BbU0V
TTaf8hbeOkxMayA/2evWH2fq4gPK7PDQOpDrxSeJ/tLgFlOkN/3nnftjiFTyv8dfwP8ejB7+sJ5e
pLK6rbtzzKYwqzaMhiZ6FEmWgnHginzQ47Fgtfz/aIdKrw0YSMId/PrQlPkdQhnIlpUnK4OE0NVo
tHarcFawB4eyfqTdQABEQi9ucpDPpiiQ9pfp9sdMLdrTlX2mFltx5jbjSOcTozwtiHh7bLD2ysZn
1HyKCYaUE/p/FqKr1Z3tXU42gqECRm5uNsWxqX+bC540b7J0lKk6B7O3X1hJaMRYnkf5BHYTh5R9
nC+X7z3msXT2dVvEGQMV3KLTkN4yx9P4+SD7grmQACZu7fi3D2ujWMwRNenvW75D6WGSKn0h8vKY
I0t9tiUzNs9eFRHzD4qjp/0cDO1D5lJ1y3cuxW+vb7BlXi9xnStmzTNPN+VyFUTz4bvsGoW6rbxb
ijaLIWjE6LLzahQss4vwKh6vKIduwE5qOjughWgz4MzBNuP34sgysKQUvBJiGMWzg8TGIt0Kb2Nj
yqxpVUfy+dpKMQ6fkcXXRHmCYHb7p6UaP2lcw/aCsqmyhJBFMPh2aj1eI52Ud2IbAdYN1KYWpvgr
9dhedAGxeDeD877EOw83CToCrpGvbWWTxaAR0wcW13SSQSjMPX9Q3tALjH2Dz1/rK64w+UsMG9PY
WUyeJsbzGDoI8JOx+cYewvLbXWt4ze3zs5uiObWWBKhxPpL5srzHpa4q+1VV2k8SMbHZ0j7g4s/D
HDG9blqW0gHDtJEtoBIK+e3EX4N7Btnsnj85WkCitmegzLn1zT9uU9f/ESlGPAT/XYt5s04Z5uoo
6wWxfH5SbYEswDOQda8QKd5+RGeOGXxYyv5UwlU/0Mh1oeMrAOpQvUl5PpbJwB/wttWN/tSIP6+z
c1yAwncgiscvOHJ+MmLMp6nt1VTji5QtmcvMZGkpuLcXxL9fXq7F329CS5jyt1k1eb/ydTm33ZXW
ebv8IdEJ/YzlpmT1CZQ98BDVDfBMStRdJdkFt1e1e3HNki8areU0lXM/TL2DfsFoRhK2z+Fi6TgP
cytv/EWtv69DsP9fvmkgi4fu7VHTdfHJKrmyOW1sWgpGEnomXoCEU5CZPPd9rVqTZHNSuiMduHts
LRRVo59/ubo3USajQ25mYSwaulBqoZSaVB18nZmqoy3yjrf/dEsgIkp41mTqDHmKaW5Gd4lUxFPf
2/7m5rBpu8QOFoDSOkGzZgiluhYJn6eIymHDsXVut3mi1d1EdclIrEU7sKN1w/08lcdYhhIQAOLY
+EseahoQ4YQtgFj9wJBBLoogK/ouPoIl+h6vvJu3W64yP/UpUY4GKf+3/yNfRN68Q/H9cohn4l5Y
XilWQ5dLhaUUuTl7T36KIoQPKN7uqyQk5qo8GCBxxQ8ZQjVz54yG30bHOUtt9iSta3j5vWX4uMT/
IixxoxNTjPsFrOry1k5jY0DXajv0Kg7hXBWoofwsjYgTCKdJqWIIueqrSOYhiCCDQRYphh830dTG
r61YhpLm1dicVG1o5MQ+krAXSLBlAJbHMpLlyAuEuC/QRYWnMXJFHZ1qcy9giD+FsNymKBiESjqt
Ab8zLz6kz/LrlJdka29ythShjaOWSYRG29ZKKDDzcXZ6Ge1Z8HZKvxY8QyaD816lygbeva3qdsWn
7uAQQadMtAD3ai2qzicjWL4zZlsgmUFvGcR4Q/pAB3v3u0kxb/AnuCVEp03kOQZHcQFc4gVszvMp
1xmPYNt4Ff2cQx/YEVcovZylEjq6KmfUmXrOgWYIkMQW9RTUAacgguyJfCWDIVZxRrN5QpDawz4C
itUGSzasu4H7KI1lCctIMMZAnvDLDPvgC5BDLMDLrkXu8QLyZvDa8Fc5/7nkbLX0izGmrxnRitlB
B/cKrvaLswLaLZkUxe/MqXut/gjXje7NfS985KzkCzI2SMTT+nlHzHOBH4VJhUrY1rqdmEtp44bz
0yyo0I6ganOelPlgvum6sVIvT37qerG0G1+x/xzqOQxBN0bTkaghiynmfXEFBJlz3p37B9kyvw3v
1fkCmJv3cBAaWP4eu+aq6jQqcTUi/v7yqFaVg83uQZNDrtUf0Z1AxrvIUCEqtf75JL6ndtLQZkwE
QwPmQeFonWXocDZuc8qgEvGsp/zhAY0tHQ2ahJMGrG4zUwYzURjoa+XwpeGHCbnv8FhYJA/A0frp
6BcOVO+QIvCq5V7esT+AAX+0IJd+6a47TsrfS7d0L5Mqkk+f1aMJOhuUKMQn32RnLLwAoZ5vXpdN
XnK6cWbHeDNYCDEEgBeSXyRyWwocTivw8MVw+9GSETqhoOWFtgKQYHfYasohQPxos4FHpq1FMS3T
1+9r0N4EVlqJ7XSu/hupx2MSd6nVsjcaln5bqvmQYnkJAA39hs2lQzw5RenyD6jYhv/+QSFsCZkx
Xy7Jf/a/7jto1liDBSieg9+WvnXgR/vwEId09gtTD2o+5+vId08yMMlzmdFasmrWIXlMjFOL7P3G
OBOAeNRIwpFC8cBKROy/GhVtDiKrGt4QKAblkd/nmFwi1O3SaZSXqRTbM3skOEg2CF0Bizi8aO65
Km30drSnUGLVVP4lsrCDhHsuEwlRY+1zjntdWHOWjZyIb3hjAMgUKVDOMXTg92FcA2svhawq1PGe
LPqAHOhgiCY34RR4WNncl1WL0MrcUkyARmj8VzUTIz3UYnPeE4qkOdTfmrrpReGXEnVeAUw+gxo4
SeZVLl0JwdJARrGkGAfzxG3vNHKsyrPvdAWbv9cDOwIVlm9+/p4nxk2iHef1hpDMIMut9qnT6UVY
ch3bEY4FMyzqu9liLqZX0hCY1eDGTXV5Uv/RXzsKNTuBGQCL7oxvUCwX9msx5YUYTi3hsjlPXBVq
R37fO66TJoQaOARb+14nmerwe7jYSnbucQYiCEEVrvcW/XEmlTzBuqXeSKtl4pWNDdp9PkXc1dru
i65UfFfeOBb9Rrn0kgsHAOhkQRUMzK4nd3Y9yU3qqY7523qAfu4O20gxEAXHihqoZC3w2IZz1xSB
LTfayOeVsf0SfQ6M7H2ryLxNowZtIy+E1aw8S+58Lm+U+cumaas03RhTRnaIdt2Wz3RNU+usd5Lv
X7hVHTteGCA587KR41Fy3SVnR7SJa3WvbAuUR03kN3+BidRkmNyqMCxA2cbnQJ6BycCTeNakuI7m
5kpsyCSFxqL5lI1nKdepd98aeOLxp8aLmYToxbGLPQsG6j+u7Hq57jcYbqHUllZagVPL6yq5XMRa
t1K9os1FkbjQKpmFRvySqX6yAIuPVeVPO4QFHE+QQtMN/pQrk8CAY3sXAzhoBjuwL9Hu0e7dqxzp
xyiW7UILYkW9f5AW6Pf9HAh8rpeHfaGFEhnksod4IQ+dqhQoGgt6F3WpwmAr1GXghWcGSOtyKyDz
QJVXP/ONbOdNo5nEFzJ+F4ZYydHZZqEXMn8wjjUNID+kL5dtx03lp7FAXHenTPAwoAToD/Oryh0Q
e0cJUXrE5dkrxhu2Bq5SdVktGV67pRcgGruOuWgpZxqqa4w8SylVluGoiENPxk0/l+wWBw3L3hcH
o26scipEI+WlWPyRD2ciOAdZPWNTyHJJLGjhMrckhIV8r4Qysu/RO02ZFp3FlEOkCCJ3WnNXNTM6
yMDv4Vmfg6kmlQRfOwfKPkHn1DCYsI+NqQLeZSwyT+WcO/AMDlEaJc+qdM9WZqE9PrkbpE7LPmQ7
lJIOd1NGUj2+eb3zqsNbz2DwFveoGtgNV/MUa/hFAonmA0fVuBqpiLYVv92YShxfnun+9ZUVfe56
VIqTBrW0dJ4PYdRQ9RsngtSU4pqxA4aA0GDAEhML51tQNa1H+IeEuBFB2gcoUXpKyMbwvH+Z/cBd
n72khYGnDpSn2sxIJmkhDP1azFDq/Au1grf1fvNevRsAVxY5inzcvl/BXiPEXTsI2dWvIR6s3VEt
SUre0YUuRtKZ9QD/0vy5u6+gir2Vs/dzk1vWt37v+uDveKSAeAZ0xACgChT7SGbDPu8uFTG/jy27
70flhs70C5UYqaenfEkQfx4EOETqwwv7bP7c3/DOCUQdWn9ZR1t2YUsftMT+4idE/yuWznX1Yj88
CpA0Ee0EOZ0zMa2NHJ6AwJVp3w8cbnmfDDQjNvklNb/chYeyGSeYYUdj4i+f4CIy7kEveuIqnZFx
/w/1IXjhyvGe12f+FmyVjJqSArfg74aH+fnFO9lVm8eO4y562o9UlAKXRDLykN4KRz4KmD8JvF4J
yS2wl6Lqk6R1kvX9Z6k0RYpm1y+s0ICdHXczUnxizNcqpLERfwGTCoLrLf3aKd7poOBr/n7DOJI4
HD5bPm+dt4es29scAVDy44CUa3zO15M8qhpUbZa+m3ynU80a1R3qs/M3qrMf1b2UBsjCyThgij+K
R1mHub/54bwpbnlYBWuIKeSiC8CjxexXvSd1weta2IRNkcp4OH8Fxk+CIo+ThlhBZutyFra9yGyB
ccOX6P8jZPdFUKf1/Jp9GfDhkCZm0O0pxlGaT3Piy+PGLT0Jgzcf2u4r+LHHjvQKjPO3LbFyUKwY
xz7UFX/lyxDhvfVmlweh6edrWgZkEIiX5sQ38xYiiMqJVhJfdjsjY2cT6nbdonJEhbUgnmt55xLf
Lni+p8iPajh51KifAeOd0Uve14eNSJ/qIDfyG/t7Lx2WrvgkXGLzKx6TuQi4N4m399WOBzA+xpcf
eXUQLrmPiOCgei+7exBKxqQHDz+Zf46L5cf55J78dmm5dcORkD3QuaGF4Q8zI3IauWcBPicxwaSp
4EcdTQz31IVW5Lkw97fM8ssxv1V9alg4RcGcku9JGzwg3vaMN4RlbWGfT/tdPf4KH6OUitE0Tt+V
N4N6A9No84p0Afv1axXZiw11WBDqjhDNlHqre+RbbluO6MWaGdTmmzxCpbIr7uT90hmX/vSHgB29
LWNY0qCa/mcwFawXeTw3mLgkvYS5vc+ZSQ6/7b0w215je2E4yL4COaNVPISsV6Sa9LQ3WpuX2CbD
w8nGN2NYFR1jtM8jwDRAVPacr9zX9DkAeWeFvynAq30l0p4wSsFGQr2iFkltE1OpsQ9QHfyM9vFM
p2u8dEfanAkkwcJBolnk9a35+8Ux77lB3kTttd1fbtljjGnpeEoYeRUge4iHB01deRlJQEq0+2mV
BRYbtZmR2RFqeJyOomud/EgPl2tPKLicLe/vAdqrvlUpDcFu59uXQWQfIYbQ1O3qoNvICbhdQsC5
LPfosE4b+oY1OWSSDFBd7f2cclh843Fozg97zyhWrcr8z6+CB34lPCOOR+dOYnOunUaisMHZmh/2
iH9q+oYGGAIyxLc4kPOLrhprIQraBkMO5DCdvs/SwSFM0OYq8aQMI2XduJ0h/5iokXd3zXcu7ZEV
E44EH2xsNay13KLP84XL1uDqjRqHUle/l4yIq23+KsQxjyRES7ROTMSFDpiHHVE/r8VQBZf1ULv3
65R0osGSAO+42NrLIOmB0PV1fPrGTtsVUKfCrRIC7KVvO52Iabd8TrYzG9B7OIzhwN2f/VD/MPKT
lJtFIrTDWX+1d+8eSvJUIUH5r4781f49TrxEiPoFl+M4//oUm035ZwmpiwBgZxACEzyPQjUuGbcL
U7vgT5GjY2vNEbUl8j/+2xRt2EaSSncVJf+pdLeWE7ntndlWs6wn85rl4EgpCZZha6abUZaNc9Ja
EPit00ST1+4VIHylhiYrKYACS/5z4+FnE9dlRxCFeuOFqwtGtypaWqgS209W4HPBGjlvUe21kGJf
FbZADSQjJQ36H9s8YXSxi1dkXNILV6GIV5V9UysXv+kAKdpgNp9Qx53ARssCrM7olSQWwtndU5lG
Do5PMw6Yo64l80AtyN8NPlyOXsr+d4p27rIuks+TELwW8LJ2LRNCo6mZRk/ZllfPr8hjnZEaDCJg
6tnqHE0mO/3EY2dcEa0Wf/LuwsQGHmexLoL9xPmPLRAE0DYRvKBZ5B7qk9c/YNJYQ5q7oAKUwxbn
vgFJeQd2UnZZcaFOtqFCt3i9z4O8IPGxTCxZw0sUmxoIH+FaS+JRwmXRf9d5LqKZEzO21d1oKRl/
8B1PQvGQdlf2NRX1kFAaEyNE7sJ+dxxFFKYRigSWT1S7cwd4wBzrSODs3Utqy2TJ6UJmPxEPX/V6
i64x63U6Fkwz/7A688+DDn2QQG1HK+3EoqluWAI6Ko9ZXq6etO9AXbntMDvvPWxxkLPjLoje50ek
RnbbMySGaNXWUWbYog2kfa27B8SpbfOaaTjmg/ahFCUkI9tZhvcrkJ/cOjqK7T9qsqdmTlQzpfhP
ptczT5TF9vp1p6GsdKTXLyHc2YUSrOuAp4DnCDksLHwTDAkhUySR1oOe2uqDDOja9+ILEwUv+bIq
Ws+uHReUYIUdixOdrA0wvGF1nMUsgRLNRpMMM/KQ+XcRC8RfwE8w6lX7y1T3n27EReTYF4W7DHya
uuT9lp1cbQw3XOONX7DX6SSQEmmaIQSfiQM2VpNfI0gAf+Cq7eVFaF1NklavTEz/kp4XSVZAkYXi
T6TxFVDUniXF3UvyInI2d42Ws3rQs9yvTFi8HgCbU7NVEPS7CypOHYlZGhnOGrrBy0YAlJNLucVV
UjDIN0vc6ohpelrNhzmMb91vSGOG0e2OzI9+169CLbN0QFPeF+TBHLyec56ENvP+WGdac8OpCaay
Ii6ghlmDS+vCOQpzSX+cEgVzUgmEyiHTkqS5XIhOejBQjcflZF62Eig+Lk2XuHp51wBUICwAbE2D
Ggc2AuW3MaghC07rsMOcwdMeJ5wpSOUtlrDqyYEhqWwgYhRluCkB0D0pDQgHBPb6esSCLaZgd+ij
8HveqP71He3LD4vTv1DQBMQUOpE1JvABXzwZgvOYxTWNVGBW9t3FyBVdC5FS6L1XIWrmvzRKy8bS
pSNxOWQgUoLWwnuRdyvKkw1FhVz2Ns9hN1r97446IPVqWUDrejSJaod6KxH+JRXaIlIBgCVRq04r
yJUTOaRqKp9SxCoCNO8AnIQohnhYo9GZ9cmTLrC6/7cRPjkc1MGdNgc7qofTxeSjTb8XAkITSlIS
U+A7S4lKrpPhbj6ytIg2KU6aQF/Z2I1Ko1O+/lScCS5bmhw7US/HWppO4YNgQaI//BNTyXe7rqNx
++cmRrHQwxaL53FlYxFBIcNjSsxWtiwIyzf53KYF4fJbErjol163qdjB7UanMwvVTKKIAVg2Vcu3
PJs03fh3rEW0Cu8SWW7w1H5KGqtRnw0Cz4TYrKWe3Hf9beMuFyPLBBHFh74IwrGIZ0J26rozhYTK
w7Rv4kjQ8PU2Vq9KptMGULURtaWKsvHok7RGIrW5v28uDHlc7+oSuftaywqBc3uJnZhIA+Gly2kv
WQ0/jBrUzUGzdd1zmZ91ordxANlUONY3QRFh2vXyjmxyBQQ10hXvLVf+1tE2GosiykE8Ij7IvkBO
F2ZMkeAnZjzPd21pHR0l4pp9xDugIWYAP7rjwBurmfal1jVG/KBg4aLqNeRTueiGoi5etstZz6ez
suM84AnO3AsB0c36YOHfIqhhhHRyVjkgduMHQyLPqOFdzh5QImqefEP5y0JWf09Im0GrlcBI4Awx
hXyA7JWb/2hj0ut1vHhzAXfwzcoTf6MOgyfe+Quw+HAq9iWWdOt+y+vtLqz/uH7FTsNCADQBFmq3
o0/tDWDAvQp+wNYlx2EGoArjIYu+CcsNmZBdF15Y2N0MwrUzP/8b9DxhnYKythPfm2IhXyXoh/O0
1FmfLCvkJgDh489YXgMyyymvTdGAYpczD1nJZ+jPeuJNadNwNPwx8mM/kCMrqJlgasvhZyfThHMP
8lkRnHWZeas/toqlX8mUarR/iFul3UBEpXv4DhIPxI3XG/ozlh0NSxCeF+BYiXuNelyb5GnFMf6s
+UhjvS0VrXVVXZhAOC3sBI/yLhsJy0GUVA7HsACvozw64BLGfO/+MQFnkVDj9dxFtCoUzIu8Sz6Q
tg4piAkwDqd6Bpz9deLaHN2WZtbKNwIDO+NlKjSoeVUQXhpHY5gUevgzOrBaW0q/5kf7cfLK0F+L
Ry+59lcnUtys5aHszamDRRHVBzhGoGI1YKJEW28E1d008jGHx5DU/K2pb9wAVz1VlxfIp8MmOF29
GxKRU7IMhAsPvDlhajr8GJqDhhEJNd7gUfxhnO4vb6RTO1p75RAjBtgFIlKrQe26d6QZAVntmUKm
67OZa3uv29tkIbETNaEkw23uLTOm8hFDbpSEXNQkXQJG7ZbCj1Ei/qPHTj/WezBLTwCA5CgcGiKR
BJ9z1EnWTtnzzql91hZFMfzGKOIt6mD+1MDHGOZ9kQ8A3dV2Lw6YBwstAI5dZCDf/nQgQpR3p+WY
YBEeFLA2wa3eeBnqYkXwqSUB5/v1fRt7XA0wfXJ8LGXQ3JvkVoCRShlrL5zpaDdeqxTfMT+KCs/7
H7esZEXZX7CfC1O+p8wztMTE5sZJz6nWvvLWhIbWM9ogQr+ypkCH1+DHNripx3SHxoVZDUZ29Q4b
PwxWRgF5rxai//1ZTfwfF8DFSDOvShKEa5E/XLXHcrEHXjtX+ey+ExDTgQXsIrsmTRg/Xu8j3Qkd
W2QW0fibweYSYyy3OdLrsx1MyVvSBrlkLFjV+a4e7LgoQJPr8CzluyyJneiz/B5WKKB7WMLchVGn
x9NJEunMAP7iHmnpzYqW1ftfLQB3b71pyOOGdkVDVu4vp9ikcdN4eL1AxIXxneZ7OJ+FJLWzJFl+
eT+GSJKdY7owvgOjlESrp/02v/Vyh7mzthYk/UzcpwetgKwk07fo/eIjnI4R5HYovkm43SQ5prQh
uBcvO3Qpbv2THXE3qAxn/sU9x6i/4aurCipfA9HHLnhgfcb7z0vywoPe7cC4G9b9GvCMOkXjdlN1
DfESIT2Gld7HiZvvNUd0ZaDDylqkpi9NVRyv/ugtSm4aPhPuWyXV30cwv7OnyCLezCBzlfIY0vJg
oyzH6crp7OPMg4dwur+YFEzmMsk7KUVKOKJ8+WUTTQwubs9Drv5v/SS3s6/GPRBPV1uwV4mig+QX
pop+tW9X2pQK+UyK3swnGwdwX4adNrgUNS8eGirQLPyRTHTwo1vY83DvoLzl5d4Uoc9KXYXjYywh
iXI/YNrvkBMxuxCzMAdh5/A5dNQCax02p8RJOaLzbsFWcy1FCOrPYLs8pdxk1KnUGmLsjlP6Lxb0
HupNDUSwfQ+LdDve0RzTOUI67TIpSe2gJGrHG01Ifm/EN4UyIO27c/mK9Iv+7QjEdXY5gehPYtvr
cLufNkedWEEoiQkAwwMCB1IWvLZLlqRxGyXahHcNx3DaI1r0AXYR8hFpLKw9DWPGrx1TlzOdzco3
r6hYaqS2WkdGTXfcm8JHZo3u5Cife0s95WWhCVbCl77iCCHGl9Ww0hqvu3XOpbUZHmohUO7Za+8D
ab2J88XMMhO95FibBWcYuj76g0LrCTu5UHS+7ieQceBUPkKydRqK9scOo+qE6vA9ywzfHBBNfq7k
7lj68r7rNav8SXXr+rolzmEesS4mDer4KPLb/pb0l3hYSTedGugYMSMnPkOcp5l0GBivyokZndT7
cUufegN1xjrK+b8LX2Cw6+4VtMPrnGaQDgtoYdhVQe3qMOjqtpdM24pxL2MGfoHSuoBSETGR7Ww4
t/V+8JIwyObvkXheksKubyCj6vINbNoA529l6K0q2GIdxXiKPT02DlJOyF3jATuAys4e2/L1RnpK
YHw7e0PzH++kbru6+XcOsOT8kDfkpyiuQBiQTEW/XsXYZH7SSbw5/L2hf9wcc964XjMotYsNEvRA
mphGaknYG96S2zB2t1glz/UIZhYqmPiXv/EX3+3srtzpLKJw56bm1NeVjYA4zy9lY/I6soXoCcUj
dl/EwaNoWteZEOLL+gRab9E0qpTTLK7e9aVLfMBR/Z+/XNSJ03pwdt+t08cA+ECBqIm8yQo/U2Yi
Nmj7JYjUi2SY3GHNIeJj0SjvgpME2BSrZLg4jI5qQRucT3oqGQWivrFQDLzPzDyattV02+PojUlB
7M53GFtxkC5GTYjbYM//ju9K/TmghgEkIny98rKT6qiqnZqyWzmdIxMWDSx/97eoCrGLjzl6ioLY
Qv14lw7NlP0QCvFR7ZpZEC/iNbVpLfBZZJBwHxviQDbIqAE1N8m/t7e9D9800WxK2GGQRKUnvAmc
qbKahssMCO1yKLkAOXzwTcCk8FflqZ90NOtnQ3pc7SfrUxwqw+ftfV7wi80vXGCQvZ3HvnVB23oR
4N5ayV2ejqZFoT2mC8iVGU6KpU4u0aL6hwNR4yjkHYOFhwEw/B/HSEmKlFTd/x5irYgKLtZ9M62C
Sfkf+2D1eVXpbK357jQAo/0yVlC0rXIV4M6PAMRWEXlU2CuorrzaNL27Q6UKjqVuAZOncZjZOoWh
BKeYaiH4TslFnfrHNcGxjbeXiZEvN1H5xtbaNYUHPzfmzD6Z1AhJYY4sjREjhpKmlD4v6a+jvxfU
/EQJ4iSTNYN8qSDehbrBM3fpr+GKQ4aGq/Gg56ntqKV5FT6yGLI3KkuJahXCwB2NThE6lwzaUJNk
Q4ixTrun1v6oAJEA6fAxW2xMntzGyP0dxSd+XyKCKc78hDqlcnzA1UbpbxWNnJLWU/9fefq/MPzq
2qln/0jpiCUDOJmKvbexgMbn2rl+e78As4n3F0YerOwrfd9T6mGhTgq9Kv2C34F7xQGlKeT5saO7
2iIk5EW3Q2uHNTEgXHYLSUvl01mXcj8VYhASPA3JXuIQ02M/THmjHyqmSJC9/8Y03Db0cHmpp31j
Um0RZ1LsvnMXGL1svf1McTIz2ii6oVpztNyKwVE9TP3eXnjk39TfCWV4kkEJz8V80lusJXFpK8jg
wg9hjG1PmCS2Mnn/s1+9/eBA841M6JcEvw5ToTki5i09Zlzsy9+40z4L88xYYEHAp5YVvqCufsnu
C36QkqexDFtoXwW7aoCdPIG9tq1gWavmHcO4FxbJMNcuj06Ih7d+puu7D4dMo5F1addsg8sqJHfJ
VMxv1BYiew8QACESKF45UjiDTJnCtERhoueMTCcKuFc8cR+VumpFjNhQbfzHCG72N801dVqoMjr5
U8Wr7X6r/LXy0xD8v4uD2G6m/XpM/S+HzuP6CmCdv5/IwL5X1qfgpKRqT0KHeqsjWDozV6tJk8MC
cd4MmrTq9PNsgWhsYbmsT1ZjE2dVKPHCz3t9tJfv+t080ZaZIgwKAoXeGWHA44eHx1W+fl3D1xS5
vCz819tDyv8CvVmyj+sUJAbFGLvh9a4k+S58yTFTohL+y28gpQb/nPZ3a3arNx887/icKQcEaHy+
erHsOPVEgLe1hAkW0vghJyu4Qfx8wW/J14bYXSYoWSxyYg/JxsPt56ImxjGgL3Y/oxee+WuKhMGD
6yxfAzrOtzklsFqgCL/zCQRXfhv0wVK4h4p898ODPytqkgAXRgsOKqprRbMqebV8l8UhGzYXeNUK
LPWRCPiaZi6e0KWAZRXXVVGLb1hPcol7ZNAITiXegn6U8kIQVQ/7KBiBE/mrX3hkWjeh31kaWDEB
7tiB4s9zLevY/51lW+ahbTmeMBTrL1NOOfPuGPW8NAEfuni3HbeVq+mC08nVJ/JT1rLtGcGpMC1/
dkWwDmjYfLTlo6l7QeKAdf3r7gU1Y5NIs2bGj8di7OhseGKmwVVCRn6U0Icz+yHIAQLzLAewRqYk
QHfxH9yvoT2a68dPz4pgHR06hXiQd7XnQwGQ0zczEw21AI3mtED92xtwCem4RgbJl5z1noeVzots
B8NCqkI06mV2Kzt4Np5GO1XWce+JpDfYJLDqLrEgq591PlOh7XpccMsv0PZIrwaBYzU6q/qNISfB
1Ru+EfF0OLv0GMTZGQobVaqX+/0faPSltbeVoDCDo493FNNwkphYyFgJb49sLW6VHum4FJJp0Sjg
kt/+/FR/K3jA4aPMxlLPQU7Qifcr0VU79m+DefhHtGv1QXuuMl+qyHuVJr9bTP9cW7ClD7tEis3n
TVr7H3b2q+W1lHzletzCdho21bGpidrBk2iE4+tbkWGE5gZiBUgdAtqldr4iXDD/QvS2uiC9sdmc
04G/O/VFhXO96cY9uv8qEWpSG6pmFW44n0YXLYhOXVBp6l2mE+6N1UhWkjT0kEiB2+VyPGL1SEaj
Eqp76W6EksFbd5VwWpk/aqEW2nX89vsFYlAb+ZRUzayCZmqcbOUY9va61UyS6VmL3doEq4U+n6kT
OT1COzV+qMFz30jmQpcneE0wWDSQFGuX0LBKTBcRoTNkBopRTlA2IYz5r0bjzNF61UYKsAPcSI0h
FLVx00SDRqQxy8mEAKePM483BBhok92LAPVk13aY9TL0/d6sP20UI6sElYRL87RQLWSkLkE6kx8/
k4sx5tuzlPzUJNWAXXzWgGmKKzuxILVZQLdiROzPHZOIMQ48ApJ1ALK52QkFFwZKbolk+M1FYGZO
moH6fmC2IkX6WT3HsHSJRbdK30DH/nHbuS2Jg+kjlFR38LMixmUWllYpiL4Q2WoppsBGXKHmlNBv
P8RKdmwhObVCamit3nUtRjt1QvXmkG81OxtryTKfcDMyyUyZRZV12g94O8UPbV+JO5XM+Wxx6A3S
7a+VCIBz014Bd+Jlt/lLruU3a56zRLQ5MwjcLo+KcVDC9oq377BpiqTOjermf07Boioi1XcDumkX
NsQE9pNz5L95l6c1i9SVLTuubEdoHDoQ7yyQLedckpRqlAC3XYRdJKLyRvS51joXGnyxIFngLhtj
DAq6+0u5frm7xX6ilXDsSokrzCxr9g1CMiG1OYqZkMp037/LB4PQzVUT/V5w3rUEz2xaDOZgulji
RLvdgWkDHgsHxTcfoJrHJCaD3Ninfo1he8ej2UOmeiICR3Vxykrym+ZCibkrT4EPJDiFxpJ2/F2O
7lO3CZtHD2sfc7yLLZt6L+5yJf/pFadXCJvsf4QdHTi7mm1WPxIP5QpOxsdOtNEF0Z1PPE+LY6fH
wqRNt7ttGR5y5SS8EBNBY3lHXNwgzl6/Xv5n4My6mjPTVP/fulOM/jiwB0fcFSnBS3DjrGirUZB9
nAVk+IOYekFaRcu25Zzt6aurq76dvC2YFxNGsuS03w0ICXoOz6k47xJJ1I6GVjhDUYCp5SoCZ3EA
kNyo86iT2RuDVdydXbNf1VUXPJ2PaqhJElYfCL55rd5HFNu/x9aPtC9DesKZ69mkz2nFCN0liNXg
CljkXReILUYiVVaPoDOllkz3uIi/RuW1lumVAmz/475zN0SV/TT8s3NzGsOo8BGnJk2IbA4jIUU0
vrVHiCuxovXEWAQCJgThmiQfCpYG0LjdRSZaY4Mn4tmk/B/PZNTF16iHmP/R9Fa+M3KsRq3ZGC/Y
6yq+9WdwZ61b8zsmS6H1djrbidUMShBmiDIkB+PLaef+pVIGa/hc1ho297AX0LX4Ub77w/EJPzkp
j+vtRfj12bFRh76w9hMi4uNCgR7++ZWyS5eXZjWNm3sZU1jod/iZOUZGYlDdYaGaMwDmhiSm2mR4
z7lA7cDEJ490Wyi0a8FwZ5q0Zp87NLn26MksMDAXcaTm1V/bQZnuvvd6+V9MevVl4fPDeTykbon4
jeKZ9FBDgpKO861Hm/vv5KvIMqbk8qPaS6kHJFWMl6aPoHSnB38yN0XFdZ3i8n9NfdfKGUf0Qbzx
1iCM6nmO+GzwN3reVEquxhUU7W1vuu5P9sPaZxDMHN0gZQNsTFnqDW1xQ09XmJ+0tyPxhxMM1hgt
bSYO2Brs/+2AfX9tNm9ouiE6dC9RP+WFUTBoFg7Wv0wCpK8HqZdMXjvh+CHJqijfOSCX7NnzPJsh
xaWElqaU6ruc2kbdA9L/SiiF5VGmT+XNIkJbNR+eZzididaUpBLsknRhonCfayOqtcOMV5rJyql4
CU9n4y3aCG4Rfw+0qdTxzFdddHChGIwz2NM9sf/k8GGFemdpUmclzWawqgV6tK1khE/tKaFd6IBP
i4ZmLf5kYgmxnIjB2cV2nrPv/4OoVj8GBP+418JcEwhZ7qpnVSVRLlfeZXgSkDL8DwYlgJ+5ggjA
s+YYiP/HxuxEBy8b7O89W2ycEmxsElFbE5lY9BVIdqjtrc+m9EGcMW5RfKPaf6E0qQCSv+B0QJWt
CPMU+qo8HtbB1gWBpISvicKfv6nO/jGW5Vi+wvxmtmkW7cfe5WVe5qALCDYpwtAaPFy4Plr9Y/xB
w/0WyCaJuW38gCxTDkCzCkNpmjgw9XL2M/G93yMGNqza6uh4n6UzUCvALfVY4GkpRlZaLXRzceex
DIXJ9hqR2UR90uUAk8BD8rH7d92wcDp3T+O22wUb/6SOjzJjUsnToppbldqOO75ce4qZmbinZoc0
WHIK/m18jP+3C+JfwLg+gsV3tBc4BVmNVJqaWsUkSeP/HZiKWVpKXPT1in/BpkjPafiQ2YgLIkJe
09VVQ3flKNPycgzeF9iOlf6WFqj2BhYlQdU96shnIbc/sLLO/yAQ8eqszRbLTgtwYYLY6Z2Rpikl
7evnUrVEM7qEQ7y8flwyL6k4AN7mxOEXzTAeZslxuXVIowLeOOrcwvZX5992IinUPl54qbRKFh53
VZ/E5ltDDwnujOHQS9VvgCGG0b5K0crYQ5pd8fuq5u1zkxW5El7TFEOQ2MA8bsetf1+NhdEcE/8t
/h3R/04C8CX5uIJVkvs3WMeEAM8fBP/B5KLYbcib9uWPC0cxVuDajaSeBmQHWWuPNFV+H/lMs9dL
IygsDoTtHD7TOC9qw6r/Yu3PGtWd5vpRVMeCGEJi6NP8vlf1Knu7Z9dlSmLVuFMMvhL73DwdcViF
IJ+wBduc8MNh0+CAt+dtp2LLDtZ0bTO8jrdsXithdJJZKrzzxE3z6GRjOEtHOJmn52ufe1U8pA0i
vTPuXlxR26vL5HFYb3PFbwURDbYuLYD0CFojUeXBlWJA2PiD0CAMMB6tbGJzaL0rk2dEOxaYpJDV
YD7u3WTcYcPS38rTRSq1poxj14JbJZmnetpQ8XZzyT3xFX2CtU1UZoss5/rlKzUXEObZJE9F+nnU
10QV40fuI4bBuH9lsiTFhcSiINSKfOpQlZg2UrzukmyukmMPdVcE3GqS5G66HspQ+uxgBdTKeUiB
EFkQDNfVFAKntwIAZNd0mynjNbFI09Rx2ZRFAWij0MqdPvFyjCzq91TAw1RrEKY7rs9VtM4npG9L
sn116v0zQJD7qizznRz82OGSoDxAuxJC+Y0mpiBdIybY3A4VOlVTRGEHVzTpOXxgoAoVUG90lvog
zKckJzx5LtMh8DDCxAJeHpTPBQynuvhdVca1sEaQyOvLwul5NfjHj4GoOPP5V9s7UcCAlX4cXEHk
c7j6lYjiPUVcERuTYOHOCoR5GDvX+QlLJX/izAKB/cFrzkn3RLH7ZFuV+xntVLoqD3D0Ry6KVtAc
4roVQzg9bu4mSAljPZLItaop59ccscuUI5qKxHh7a+PV3AgEiJ/LAMxRQb1vmfM8TQrNNGJbi/7X
+8+AVqZUGF14sgAy/vb0k185LUPGuqGiaSpzUvX/gToWZ36mHo0o3laP2gA7xxE5jQJNtso7xpo7
UAbxG1yMyOq/9LTNk8sjkv4j0k6NRA70S97/HJ7PA9/yHgRPachzb17EoFyJb6PLOSWbZ38sASu6
6jqrzJWWVc3qX2ENFy0hU30U4gaNr56B7GJR1EA168EzNSeSSIcR4BRz8wep3vvzjZeg794zNX+D
fuLmYD5G0aMctLQ8aYP/7/mHtl+AtrOt7aV+fUH8FpCT63omeDudhyFnC8YUQX/c1V8uqke2Hjbl
Jqbb9ZBVhj09iiQhxc0TiFsw8tsypHRMN9K2adSE3cvUh6842zXb2EdDqcqB5fCHjSNwwUJFjKGy
Squn+USsi7ODKAEheyw4kw9B+QFCry4dOvmWbG5V5PBXCdlT1XMjdTKPdWgeNevqaWeXQ3fv1D/+
NavVo2/W2I7imu5UdnTbu5PoOiQPRdm/qyOCRcGr18JKU3qSz3oXCO3WwfhWBUNE1HZGT5oNexMF
aVrpEyS0yNQGGnbnqLpsJ27a1Bohp89G/oQgcNPeYzIO41hc7Q7JAfBLudRWzhOTiIdsdbkf3z3z
b4yeLAxCX+HWbhsGkAAp4ii8rxfXRqmOf9yFA/zoj9Ru9hJjZeg7eR74ppAns29c6eGjuCUpuaK3
BP0yx45V599q1ly9L0Ixs/vC4OcIA94ilKX7wdNVwusLrbKNkH4B1xZtbj8Zy+zMVKTYFlCqYllv
oeU6r92osX/x62zPHQ2B1I9QDwKpFLTKOsh3FmbDjPxPnAwiiJQq1Kt8Q/G4T1LmCUkKlzBAevOz
lx5TjQWyjY6j8HN8hooB3D9fXh33Ttz6vxgVozQKIh3mhri20p0h3Hqb9SePz+a0BGeq02UTh/7k
joKhonvIjJ5/bDPdkEi80VxWFQiwNYeaUihsVBWR/muzgzPcdbYHPpLQdLwhB+rk+TqNrJQcRJEs
sM5/Mwgikwhc0Y/gnHx4Qr3wc0TlSFzIijpR3/4LzWshQD6DsVG1VAxt//0v8NHQ9VHDLQmAXTKp
+pcJfFSSWVjTQPsUOaFwhq3YhzRW1k/ydboPPDQKq+JUPv5cUSdNnzECZFkNj6uy5B0T93STd+hw
VdQvS03LI+cls5ummmYDqtblnC7VffjBYc+b+I+U3Nz8ywXaUBXbXu2CSo6wHCzn2RBUd9QPjn/K
NMRZgZxfQlwcLrQexOFidK4EVFd7lMMXiRy7MbJcs81PxjV9ENWvNWM+7Bsbn6BTExL+xNnxYbQ9
wrxkoUKDPzCW2e8Br9M72nZ3BZsq8FlbAfIBpEUKOPgM2K5HvYp9cmwEZn9JWOP80WkzjlHBtwMD
a7h7txal7BdJZ3vy/qkV/BW0r8tPHmIMVOU1geqVxwFTHKP841x9Dlh6fLfOlqO0IOZEgv0Hqpvg
+6skPLoamdJVDCdDwBC6InnPc+Kj9q28sfBp81py1KPIMIqX+Oo1XXaWS+ZXxtE8S4wMSpczkRal
yAxHMc/cYxJiMyN0A+7N+iVxkNZxUiB+9p2UmkZwHvPNOuz6bSnGuWv5ACfOQqiEZADOgubU3l6J
5KXS+q5sJpwo5hfbNc2lpPLe39kJJ4S9jWdtQDBn+GeYIwvHymUMKofptxFQJO4fFSklopHhXzeg
tb4eZ7Ikg57ZYCtq+M/nwS8dVktqlXENH54YLyyQJVOuN0mPMSjz2sOCra/Lp5oaXQ2FHtMKiCjr
yvVRYYLEvBunhmoq498Ng1qdAMEQtnX35kSHibXrY/csSZGM4J+Wt5SQ8hIdbRDzAg2aRsya+DhK
NS4RvzTtQsGPewO4E0wzx2KXqbo7UeXyLSdLGoeU/MGJgD5GuWWTs/iOM1AYfBKXhFchClaKG0fX
DQZ4nceTtzuQCgBGEC8xlhomK1s1E8sgvj0NO5GJWvG1i2JahbS8YInVpONqyajQOE3O84saoww5
QBm9MchcB6F/0BZRTGrFmGrkQ7UtGh47YieoJzZZfl/bwIyAY6lORVBxrHbZO4bV3Yk1h2gkAJy5
HJxCPCW+FHJAbJbMzHfb1MzDnBCO9ak2MTJ25VxXVMwG8MWlFmMQxof1mFcygYztGgd4mobTsWYi
KQ9BOVZUlHsACbspquSPHf7U25JgGus+d/wuwGgtZ/WqSqUgMrDsv94dnTvSWcssgivEqxMWSjvO
6kGVRe98INiNNS4ui0V+r8nCj2DVK8Gw34EnsB7YC2lAT9wYs3sVe+s4blHLX35D5cMMD0F4wpeH
/if42uF+duOjbhuP93s2LpgH7TMzQQy4EEwEVbQqPGwOZkcZAq0jA9yXK6+NgE37gqcGQzHgfsqJ
PIKGClPzox6ZKVXKdXZWNS8F5bziQakXLzfkZRXjDqNS5Ph1mMQQIFsEakU67lj9+4Z7yeW4UY4h
Sde4P3UyMYnDKNnYInvfJqWxN4ZixlHCOWbDNbwdQKPizFcjYWp24arcn/DoRSDMA46C/qt5Zdua
CsaH4DPgNn+fa9FtwJLkO5CyemQ/E2hbfdvx0OtBmJoA0PRXPTrgQ1kgNE+l2hLkH8fW1bDUmXE5
dqr9QsZBYWoBaYlM7sOMSLJJawv4P8MvkNF1myyeczfwNxai44/KrWVXsCqQ8zq6Y6a32V18DYX1
fa0B/FBrl71BKpvaM8hBCb/N7Lbc5UMoYKu7nCV7N6TxySkIm3t3FPvDQ8cTmvTMfBfjgsIJTYlq
nPkBGSBboOqiq5wDX2QI3mDISwRf173CefX8JMY7SC2MajEMDmpKMOfoJpdvBs8Zb2klC4W59xNd
EgYBBpvYGp7SLkvFbuRR14XYTMZkOsLpe60okDr08Uzvz3pdeOxH2c6FNj3dtKfELfU54Ge0E+r+
6tP6vsvkXndYw2PltrMAYtYdotwqWGyc3ujwEvwIaH5CwqMq/8AgJhFI3BqT2fqmd/LcDi5FppnR
6fd4BXiF40SUQ9obgE2QSF0hLF9ssKrukqFUkznnPlKI0HS/ush7j1ge2K28x+w7KrOQkUIjb2n2
PVMClZQ/Y4+V0O7qFFPEkL0SEFAzSaXn5r2lIZ9ZjZObMSTRpjaQ78moRebDOsCsGzq3utuvjDvW
p4/AiyLdpDsdE/mSzB0oqI9m0wmo7eSW3Jl6yVzbKWhugsyM5Mjzjdn1VJa1CV2xqWqVXZH+pS1Q
zGD0wDiY11Y/zUF2hDhEi5vSTEwuwa3xUXad6BC3SjzmAWeiA1JQZt3KcwtKfMEnoMxEHSt7lVBW
H+JSQmaFCpiCYcRH7SjWbdaomxgjzpjQv/2kY8tdw8te5Xj7uocCUaT4/lP94zLn+EM4THs4ALUH
LW/0/OBuTYf6fxTqcAk6n+dBEcAsV/FE7MXdNIW53djzZUUcCf4vxJkJt90YGAG856s5W7DYMyo0
sHFa54EyM8Vso3ub4ekxrMHULGoEx9bhmdqaeCc1vr5p8ycdiN/4VMjvIzK3Sk0G4UPDIw9PnX2z
C1FkLLMmMR5m4HcQAUaV3cYWboNni2hc+2QZP967VTQsk10tmd+GigMJe8usPpscy8OsbhCcoegt
qwV/cOcKJYMp7UYTMoaios22zetUc+YYK2dTv1tQwSYEDA3fTbjgu+j++OLKKGNFCj8b3p7b3k7x
bcFUaITZpdMLQelQsAeOKWSBlvxU6pkyo7HJFUbSmq8uo1ut1IkFQDsadNKJkcSEFU99A6xKS458
E94VYn10azCdTLEAm+AgIO+QckgNzuwtu7G2gnkrjm7zawNLABmtGPAZHOh+zLpOVf5O1X6WS6dv
zF8uHKaGdw5AzqlKu+StLy2PlUbI3BQqLj5ROcAN+7dL9xE75Jil/idbwaH6xWJcCVLgITMNsruH
T4QV19lAqLh0Xg+iZEKl01GS1YJPf65FeQTqLN3v6M9mmtxw2UuGSEI/aUXzBbrJRtxqTYHa/xMq
gZTWrN0msAMrIx+qnqYDrJ23HUigtMqZnk/JVm+TtT3uwCNNhpVCCGsco5MCOhFZtkLWJZw3kipY
U98XkYc5cnXs5ZCtdyEucXdLUbyrqqWBtsn2TN+dkw3wULuwwZcgr/YgYnIL7GCE45Fv6f6cFV/5
SbT5pbVZsw3byu3wfwFmmPxpxm7dJWodvpQPAP3O1S3W/k5MLC563GaegXzp4aTce1fZ3lecrHrq
0+pYKHpi7Fe5lg/x9bAPJ5NhdiKzgHMQ37l5z7oJK559iKrGgETslZQ5f6lkaYld/s73iqr2SICa
KToDKP3kzxHeY5iHC9s02n3NvLn6a/daUFKGe4nypsdHgpLNB6l1APLMhXFTNS/Od8P4UCTdawqy
mA55F1uTNFid09/mGsb+unxiN7YMmjYpqz1LrpCMBkrTqNg+15aK+Wvz7h/Muizav++s0h5EdpCe
Y0uCU/z4RPw9MoE3fCdQFJH4/nB/vNt41+ymU45lbGHMBFHlJyVtsGEFEec4IvnyWvS78YJPfIdh
Oryz7apHuRK6y0IKWvBReUAF0ya4vov4P/8awELUH6X+4k0/5LauYPpL7j/MrirSlN8HGFvSrZwm
ZxHvSYXErWmR4Aj4k7sCcoKU+s7yHTjxjKi2mvtYFCA3HQx0HFE3Wrv3xHMzkLsdDjJv/2KhW4i2
KTJxX4DL7rSGEZFH9ZC/eKsusDarHWQ6pjHU8AyvqSW4+yhTxRudbY2oCFH1/reb/3exPX3W4wiZ
oN5aoBWlC98bZ29gYLD09TGTcm1kS4Mj20B4Tg/righQuZwHkSYVEDjJeh0HnF37YfkitOTCGCSo
XWZ+J2Wfeh1rLkuBGs7N1oAt49Wku/+YF1rkoh/T28r/Z8LmQyhPKUTIAQWI4TdWJgvsCNZ1ywst
AyrSpD/J/ZUmZLleMo8mZZ+w0PvQxODygrXSI06PH64OTbx38TGnFa+cgoV1sMnjpzx5FcBPbHtE
eqTebK6YrZWqVtlQqOhiuIceH2dGmRDefVrsk/39ARYENoo6AUdriuV2J+Bx4DqJ9pxCzN0WnV/q
aLmIGrw7i66gfZmZ9titx2ixDaWqcnhmXo/H+7cXaMr1VOx9JkijtowJpEVMIDxQQM8t247a1vSL
0gTthW3OyG80Fa5fhozZFR3miMdWCirO/qV22dx63bzQTj9wMdvEDTExxWAFrkuc2o2ac/vf07Bn
VY4uvHFBgBNhsR7wHRrLojPRSnQuMI3Vf7pM3gSl7QPSEK+au1Aao6O2SJUN5rNX4xDwSzhIuGOK
dqBxbmT59m1FDniRWR3sVDaCI1hXx1Gv+mgKHSv5L+4+W22enGH2zBLnsCq2sys+EHQtPmjIXaW0
Q1mkfWyRZugPb12Fk2AjQotL1PO+4s/fA9DaPxP6Px7qED0QnjsX2whDze7YX0WeHbj6UFCRdXTY
BuPW9uyAtFWmwRBKi302gzcXOuuTvKvY4KuoF0tpL/CEbTn7/zevrUTV5UUfdSX7rhY5QQvTvs9p
RuIcpG+WfSaRYJiHHac/xv3x4wgCsPrvHtpK6W1FhdpwKeWxN8OO15sl69UBQmTH9hevy4T/i+V/
y8XyLEYs44SbPTusS+E1g6Cl9tMp+UHvY1xg223gqGGYvjt80xyoONjGFuVP8AzyFwnSz2CRyCRb
x9ShEz/I72P3qQbi+NwXVdbvsEUTiRXuWb0IcCsLmQyNK5zx6G1tx8hO61yP5cT3yqO85iV6ZQSb
Mq0ohTTNWK7xdEh47R+Dz8EHDTcu0fjFVcWn/ZQBaLElHCTeEMYkmPgv7in1IK4Rt+Clks5AofC1
PbFWHgkPmuS7fPrgHV/8fZ9e4L2f7xeD7e4703E3A4ZroiJkm4lldSWq3Qf4Xq76r08M0ZYzJ9BK
JLZYIx1aKBwpEftV85EPxVRMpztksi9yJbJ+9TWQB0kr6t0qrpP33d6sHsSHMEw/Xe6XKS/7qP/L
My73BvmOTGRwu7iplt6y4OiZ878kjsckbs9diYlbrvNsRGZsWS/0BDcz6xxV7o1BqrlkHWdVI6cj
QvlsWW+dfVf9sGlgMkLKhMKCPrxNjr1yZ23EEbSLQ7VwgL3kLVM1RFOccEm5apu9iUHV1KyKi/I3
EG9nM9iKGnJM2Jf25RLd+D25oonvubIsbKe2gE9ne06Q1u5qcxtRc15kx2DKTKP5MMT230YZ5TyO
OAT4DpoV317DjjgVlNjBXfs9Hbz4OVJsoWObr8D9gi3b/fyDfmvr6WSPyirYSBHYbNMyh2mq3izV
0glzqxxjNEwJpv0fXaezvYBFs6pM4mAtU9Sgpf9Ia88aLMQ/WpbV4NoYRe0ogxSDYOw21dBwZxkT
RudTNsV2C1DqqM1yUzM3oo091PZ1VdQL+oNZihil+jID+nAwOguaxaZdxsrwerqaKqQXz7KNAImG
dUFEvCHx0GmxAFSctoyXdIw3c5mmUwSn98A3a0jzsR1o0HOth0TBX+N4a8j3mDTX5SX5FDoNg09E
yeOfKfNDlSt0LbDjE+xxVzsw5uOizKyeowkffHeABtrxsjT8pXfkiz+VEuF3Ru493CwfBXlMx90B
jg/LnfflztQzvdkVNbqB2Lp2n5d93JD0b5VvchYQiViTwvKjAAZ2VRpz/+C0j9Dh1gElVl6rW1gI
t15kUl2+Y6g9aT0kLoxpboOnKiqMbfAeH9tp+ndckErrU7552fksgfaENLKy1PdINWso7jjZRpQk
+qiW2hEl6PUfUTxJ0coBXZY/cFs3AQu+1BEIKT4rP/dcxLPfFvk/zGKh8n/PrM9ZAWNTH2rJioTY
k54YZLJi7z084WkYp+mLM9S9YSiIbHW1jjrLCzsRaJ5qAX5LEsMI1VApfKRWFQcx/NHV/IUvmaeG
uaEgLRLYjjItalZC/4S5U8Y8LpAbREgkswWzuVEoJWsuyBeggg0BlOYx3ZdnPHMH0z4ZTcRTYu0y
QvVZchKed5i70A1XHjEjqApxtAo4buMpVcygMgwigQ25QNyLMLVqqwcNLSu+5T0QFTld6Qsvcl49
mZjQjptEvqqi0LfVHkWdkYXuoeRaJohSuNVQh8mtIEs05png2jtBJu4ntWrHU166jf/Jv0tc+85y
R25ltrkgaaPYo+UT1a0ksuf10d/McfOmSD/99MHITqGJdtGK1y3u7XeKlv7b4RDu9uNA9bUB8uTp
n2Jk8YTUdqvLgVfnHxt7FFr4AmoB5xFUaH7t5QKV/hYphBed2vRi1eXkKi3aMYz0SatYT8On8pAZ
v/ez7WVt7oe0atFuOG8OnsPPDV0sjbD2Cu9UoBlhvvHjIAcuJQDgz2sFA9sbfTfj87p/oQ0kfrZw
gKYxDmwA2F2X2yELQGs6RbrXMNUpZHQJKkc9/Y6rvaAVgRraZIsRKR+ySq8GNhO4LrT4gLkOnKl+
A0TIPl6v4uVrr+l7/ggxLQqfdHz4kf1wShzxAMFUxUmIYMowhkV20gfIkKEX96JwSbhMpXi6xz2E
kQJSjjaXt9MWdcWNwqucWGiNTqfGxRuExX8KxBiIG6sYvuruNmRKvPye18rF8IHUU+JClm1eq68Q
yOOYPiv5AMZs+Pk/tm6ccKfF7ZBy9lS4Q2/4YTsNVjECApZT8jgDsTitw0Kbc6QVMx4hmgfbC+Rf
fTt696wa7AON7VbGhhfoDX1eEO7IUWcbAh729HMjvYUWHt0fgkCLAo7DvePjVQ2kyM6SdHaKX2Lz
LySDXKMCb7YyPE89HgP+KLXM1mj1DtkEw1ffiSZMjLv0hxL9boDjQKw82GsXfiZd/5RaTqPkDAee
s5Map7nzko2p9ixxlEya/OPQ/y+y2WLpnzd3ALSqbzWmoY924f0+HB1duzaw5baQa8CRAtQ12+Nf
oe2REPIyB7bgDzdGFK4kIYBZqgtC7rP13129BDjcgFSKo90GYP1wQWu7VTrD4rufRHmL9Wj+zCcI
CPs1qELkIyCScaDdThmwsuEv076bJFdiCrWPGqQzlIqvfT6AEOJIsGyYmeYsAGAbcmOZBH2e3JfM
luDe2ucVJp/GBFLGtA+jI+mtffjwZ+JymeWaEHZ+ieIafX6TqVwzxt1mToeP9FaHCpbkUf/IXYAe
uQQvXuT6CYKDwzkGhlUafFsH2k8sHPvfAYmPqT89NEbs81C6QSgcE0eMByH3Ra+xxXKKjyz3Po5b
zW0oaZc1NltkRe4IgP6wi/j6XYaSa/In8KhrTlDpyqSgkllViFaohinePWfl6l0WtSaDE6Iswpe0
Xhf1QK5xCdx3/y1F7+i7BMxKzvWjCGclOAMrChNFtJu9g+RW8tw93Shg2EhigJh0y3S+Fk2V5sjS
yeenna9w3pmFV9cSILKz5L1mpbe5WbGRTaxjXR9CKXHXvseGCbs7CI3uMnIWU3xx2y1hkHRVI7QH
b/Cl4bpkQIfxgha4OxeOL2QJnYb0UoX7C1j3jKCxtfrlMKzlBmcuRzOBpX/j9nyb1ipM8DqYYSWg
6DidsPsW56Pv8ka4p5u0JfZR/bwhaNEX827DtZrrS7ivgrdl3/YdBqfx9JzjAhA9tN3sE3m+7xuE
0XlRaijqit06eJ2Bk07DirY36vVfGv4weGinhDQGhxeUwqzN+jw+duv/NBfX/QEjd4j2CPI8Hzi4
10X49hTiwPAP339XiLu7QYc0vO1lXdCZlhl9rP73PpE3AWMuCRM/MdzR1hWj5VdpPSpABhlErrNF
hFMT+lc65rwdyZdoYn9HfYWY8pS8unV39KuFEM4U8bCZECwxwJOzFQqlYHVcut51Kobczn8wJCXC
+REIHHI1dvx9qaFhrzltmL8eVq+AKfBSsT8AiDXlppfsyqs7vLQud5XJJjplT4w6lX2N7eITSzRh
1e51viRY0Hz7CvZ1dYpIbWdltHuD2lldJib9+EPpob56Hw17WggFKxxqfzAXes0clnHErlAqk+Rj
4UgVu8SpDa/Uf2bv/60H6pp6L3iesoXaAxD0VSitxOoqwtxBaxe1qrS7FOzV8fBT0Bsp7tBTwpf6
ija5pvt3k5xgMYD7xi4SJSc2lCaiVbedMPiMyeCvgPVfw9s5msj2xIb6qZlCq0uzQ4EuQiDCRziw
UyAthqby+7fprqVQciErBZ9Gmc3OoRac0zbIh6TBwqb/+RTIHf4JyiKsfzFu3oRGGoysIfFv3xf1
au3Mdf3nTP2NY8o52MEheqKqc5wbiC5qYOCg4jKHvfJvorYVTr/f9fA0znAYWTwocH63FVRbFni6
0ZN8ztAsAhDRtjXXXh7Wsy/7bH/2gCuEWys0z2TGa538Rs2d8x398V8cOOrJJ0cwWyUChfNrme0R
2RezWoC2D+usaNLXhZrTURyrZtmPupXpx7A6HbBAI3FG98qugyLSYmH2nfZoHHFM+zDg7QM2+NlQ
UiimZK67FMI8WSH5eib0Yu1YxEfl6bwrQckPYJxFKXDhzxp32dm31KQ3Fr4zA5STQ2qiikna+Llu
blVFdCLYCxXhOaJxPmzxb42D7Bm6p3b1Xfy+Z6/iukF+IwmucfSX4NV8MVyg2OoNU65R1EjJLo7x
47T9Xm4+HpYccoMDVxE8742EhMlzBf530RiV4A5NXpn7oQGY2buRtFKqBMrFyAqeq8jJxFoXGikC
fu151p1GjxMSnTRi6idTQWS0OsGiEuI+UMEOLFCPFDDabExvD/uxxANsNB/Hxrk9Jid8T69408lg
5JkMlSLh3p6yj8L4tTKg3y9hQrEJSaQzdb5aE+0rlP4S8dNdc1HzFl8wCwjmkJ+jwemdC7JYrVTy
n/1ByLu/Tkix1G4/wXXnwt26phI4vPLzK4cOaI62zG/mQ+184uYW4QCBWH77L3amGx2CEypYCNrt
iZPKfc0rE71E7zpLYhqhQwFgMQyjkCtUteCqUxKDWCXoWdzn71KSjHRHCLncq8pzFh4W6YFX99hM
WuJCtddCstd8Q5ziTg3a8CfAP2mjQOCQvd7LtIsU8OZxVWrNWR4VI+abhYTn6RXVhSxzppsEoyJq
jMNDhaliGU0FKdZe/I0eYRVIH9B810WCkobPtLhV29e5iCrLmurGvFDwIN1s8zTERm31MatYvuFk
KuitEXvG9CsUOyVZ/t9ZP2lslobk1y74n+J1Y3/XgkJzF5c3btT8jPP87Oz/Ru4+gEfDT2P3F49O
h+AND9CykauKmV5NNpu8mT+uzYtk/vk054NwcJu0UIsTgxy3mFLVTp1wzykWK/GjubYRo/Wb39QG
jGDkIuk17bDYGIOcIN1d4sUv7f31Bu1urse8Kp8VJkT6B6VPtzu181EF15pSvekn7TS04WZIQSKB
mplxLtwh4BRPnEhubglu7sb33AwKlznlhxrq7+uvuAZHbIq2oQe5lpP2dUK8HRzMf8KoanURAQdC
WG11kCPUqkALZ/6tNhdL2omqjsiWCb3wEXUJo1DrhrAih5DNC3pxM5jv9njhfvctWUSF5UlMg5uc
BXfs2puBMxvV+IDqLWnFgD6Nu8wmx2oj9uD5ffQlxbglSPEm7+uvvHpkniEVkbUuUW1zBNDAWQys
lnGS4cgzIpmJvCo6tfNs8ZzPmx/xVLYZeS2fZqzXq8GgyAQdMiRA58nFgkGkWoJIvmoCeYfTM7Lj
zdxQacoJrTp2P4ty/DFZ2M8mlMKHnyh0ffBUcMBIwQh6UQyXAFtvvNw7qFpVv/NlSTXWE6tsyYFo
kBv+8grLvRg9AAehIISEI8E90JxfGAk33BserlsKAeWR6WnLekQmoxMQe87ZZZoTbHaZ9AEt8kHX
Vwzeo9JetrGqwBVPSxIAcPJ/c0inx2aiG9EIAg/uEYbkw4YmEJj/7C1ueQCdLbxbKzGzJHCecE1n
Ak4KJnFWXao10/VgkIFWTx24kRjbFl2qpes7UMRAKsR6eEytVkdad4M8pbzsEUHCdd9q7iHVQOl1
9uOcd+lzh9wnnwRNUMkDMq6BtPpFS9AiYHqTTys5niTEkaFeKjCwxV+avqqx/LsZ0H+S8l1bhekn
5QE5jZTD4u8jssdBwW0jYHjDT7nrTV26MqnopikKG4itQeWUXHfV0VYmUypST2+fGzv5qtv5A+Id
23qt9oUfQBZFE3p7ICzo9A42ry4H97QcF1VrPv19ePJinBoXzgGbG4HQIW6+FYRHc1deIk5aIusW
BTZSO8VEjTrk9NRkOvkk3iJHWAHWsf1HqjbUQttNQ5GoObGGvtvbI4+yUFT6GRFQ9IC2zXE77vur
hcIfitsIKETdDoAWIZuoTc0hNVrmPzgPjiyzROuOCGgGeXgjhBDaRVpXpSkcF95FHN6J6KMkfAP+
gnFmxeGi4tCaw6BKXkB79h4A28Th6jWTH7vyW4PXAUsCPel5CPbwtR3nsu4Oo5idx/Kmerk7h/Dm
xGW49luafwSDiJoJn+OpmhifBD7P60yhjamV+UB6d3bkRTpgnvE9U5RaP+PqlzHUKNzzC11xqZCf
0Y9RS3VjjoqJ0bJI3x6Sx9sBVOigOJkFoSXkqpn0bamDWXVNflTzXOOXPBYO0YLLjsLIPTAujRH4
DrlCuWDBxGXaNxYEIxUlJBbZY3CwBnBwHlGOFO1x8C3WLTg2FY8WtyWvy99nIYyJK8uy6tQnG7V3
/a5bQQy/FG+/hwxApm8R5RclrQJp7AdRa2hEUYJN7HwYEdLjylnow0n+5mNI9fwgeqyjX+8riZAV
B1qPYfrjMlukpvqzW/uETaUBqi1c1tykruWUARmTJFbu/lanVAYmBUkuMYeLhB2wQv/sSf3Fa6gb
ezjVWpc+MTRrFHIMmrKm2JEhSEXuk1JAgjI152yaZYs1u1X+qziMxtLLyrybbaj53qk91ABs+lX/
MBAKe/0QE/090noU3voAGYKnCynnKy4xn65/1C+lfCinq9Ll9SlVPNoZK5hLHBMv6YieA38LrXsZ
dkJvPy/8dwHC0JpKWs5FiDhcHRGlp8j/rqt5ImggYnK4gH7ZSe4nWloEsY98rrR0gpW64cjLi45t
NBaIMifM+bJuUuyg3CLbRqJT2CgREA9/KzGM7YFvLLD2yKFkVTMgpKWcPUMvH1d91Ht9NlTRFVX6
Q+Gdl0A9JmdSN+UbMYyv4VljpZ8YYyrAldsrOmG8DIjiqSHLTU9ZThj5xR5DnnvC6WLY66wFXDgi
rYiERHp/JuxeQVFTo7mDJZOL+doo+Kpq2yzyWLqdzWeYzW50w0wFLlkwSvEVJ6KQemeTBmfT9xeK
Lt1WG0yKs3JbpUm4P3hcgi+YbDiVm4Qv63hjd42YCDrz6Ld2IwwmnAJNln6OLeOk05to1CQax9tF
2gsONjLh3mQ/pLiZWZN8Lw4xikmMB2WW7tf7OeL87tyNfnqzImp3k1MHsEXBgnZlV2DwcZpq1lWA
D7HqSBvARTdmIiMy4Qnyf4Go1PO9iu+pbcdS8xLnIPMmFZdpNPrfA/Z0C/0mHEi/BNAzr6Hn0fyv
Ad6aELvC3lT4st2AZ1lnszxjQgCesiPOuWG+NPDa2sOs6Ejigw0wNo3C8J0io/BVBRAFRm31Ht73
EQiBiTTA3U2bSST7Vvj/LAzg5+Fw2cXicHwHmtof/MsfF9i826DqgI/8oVaSdq8aV9Tkg97z+zBU
hLJJ2yywMhB4CDgI779h5c4UAIWW5Xz6VFsKXuklXMIh/0ukaj0YhFlwhpxYpk8ZEro/ODRgYX9w
sVKlMdYmjrqvEjmi5jMyWOovcQZgQBBpAjlipOIwK/Cz9TATyC57mGUMF20XTolVhSL8KATL/LTT
agafsJp4s9E4vB7EBZCNxHGMwPPBSdQTuHn8SeyNllDOkPIVaNX5Etrej6/kdOlZ6yCYSUt2/Hp2
Z4gu7PyW5eeHTUKaLhRsle76Fa6r5bakvb82SflE7h2/ioKTFxeOs906PwfrdcbiVfVlnUHQw4e+
jFkoHlGwRQlEc92/658eVQblwArTHvgRp87dF3aS78rQ9hRSO1g+5Y0pohgGInmQVb0A4jydWQjJ
OpkGePNzPTRUMZ8pLgL1coCzzYizQbbG8cfTLaxtzscpu0dvGh6VWPVQVjtpHX/ApBJ0atcMLptR
+8n1xbny1kIvk8mXoSlnSEq5US9Xek7r5CBZcgcd5mJswFg0QbmqXQK0sbvi6jCW4Kj8xt22BOQG
Bg3uNMPajAcN5CDXl+rsStqnVq5VRCtuKxuxZ/oc9GBKzK6p+oqeUu1qn0pzAMfSWCjOw332fJj0
JjqCvUjfEAPowGMegt1+lzCFJXlXyVFdpK7REmZQeJq3fuehbmSTuhLb6fJ+OmkbyyNP2Gws90Fh
UpX9ovsIV5KDH2P/b6LMjLInfiFdZnC/J0yfFCLdbJ1ISa80e/LhNGVaq5x/tmANDMT2eWWhGAJA
MXAsGnPO5S/qc8HZo3i2XdTA7gHl5gTxQJ3NdD8IgKfojWGH/aIrXhxS4GodW8kbMx61H+WxoxuF
foWmfcQnVerqG2TbJwZvq921cB5Pck0MTH+KAenDnHz6Faq1Otkz56FYcI3S9NF5RW+qAU92ot79
AU6xyrX+xuSasHbqRcJuNpx7cOlJ2eTd9WL05EOivorF0Hi0tLuCeSG+1AFrxA48GTffCL56DIqw
DAwH6aLO5hwekY6JWnPdYbDq08dE8KTHZ3XkTDx6g0pwXknAN+W+u54RpLyJ6SBlKPsOvTwbdP4p
fiUcMscds+LeIjBJYgqVj/b3nBrncyd4PlQHlfftXEXVlUmeBuvs8PsZ4w/ugsrX2FkQL1hxTsSo
WfL2AT6OiroR3GobaTZkNVJ8IgN+vjg6FuWiaEb4yxuvq5y/o/K4xN8lQ7RxFJRKnuzlcdJcZEGz
e34T08cZPTZKauwKEtf4zVzM8GLkl2LXeqZS/2tUS3GoUVo80lEiRvi7KyNsKTddTezj02mIJnPV
6WFgH5Pzroju1SjzHRHl+g6+HCgJktatQNozCJafo2qU279TySWfEfOD8iq8hjiHgWOhG/adjCcA
/iNzn+yYQzYDWPzqCGT4dIVDSnZ6bH1CwFfqH76s8sbfK/0Qmsf8Wn5iVTbjBjNKGKFJFbE1XViz
rAx/60NsZB638UTXQlGaPY9LnRjzaO6ZgIGXtgv17QGfL2YnR3Ik5IA0reRpdx1xLeaO7MWfQVni
HUv7AfAxSDHt47iOfrMKnh15lVKptpbY1p6fbJxbURmBVwtcPjPrvoojyC6Y/IKjTBtqycfqu+2w
F20I2GMwfpIV9p4WYei1O5hgHoNweibZUVyTYpYY27/rEJ0+Pxv4JoYtUze/M6peXAdUxZpXpmh1
tYMO0JyQV9K3VfFpN4WPBeVfYe2klUX21mU9SS/wJchsykmKFdt1ex95Z7c5Cl3T9xShVO9w4eLF
nrR8mHM2DuogQBywsKy6FHTQcwO9lW1+TCxRWcz6BSfcSnP0eHUXyG7iMXJUTuhgodCTmyvptOa1
M8TcAKgvayBvIKQjR9CDIYByMW6kmzlw47uCmuoHUEYmhFEfUZoT2LZvSMY9kObUKnCtJN5SK61j
yXF8PAIhzRPkGJmmXbmM2zcFybQ9jQa7mdxDKJBEF6mol1EJBCLb/sYwqineSaItR6QZ+FB6vZA6
/96NizDWQesgIsottRrHXsFoF5J4vdWK0sD/LdgSxlbgWiLMoKiPqKyQSKFzWZKgnsFZQGIIjHun
8wUHo2DPCDOzOeiizQZNLg7AqRLOAGq0DPRsk4DULmX75XTL6pger6XFHRWL95Pv2AlIkMznYGU6
u6NAycbMOpkt2hOVKU5oh1K8Nycvl6kHRAD8ztcB5mBGaKXvBy4CY+jcUbRQbLXP7PeolhDOA2hE
PO3KttvavVy0ma/laX3hNwr2h0xVgID+OlzbHNhTOF5uogEZ5jrTiccB1MVM9uLnc/qfvBrSuF7r
BmuHcJi62KvmUGNe9RwbUQHnyLixMcxiz1p4QgrG240aimlOdq9jKJbtnrqw8l8ynShw2Ns92+HS
cbQyjxbenEfU68asGdODem8wABFGg1KDR7Ffint2tlkjgE2VzMKJq9CxaA6kAhYxCY8FlKPpz28x
8audGPPWX0RuzB6ok0EgUsDqIGwXX63afrsG0/F6H0GKCWvwZLGb8G1lSajIo85qmqmuDycN4yk8
IIxWMt5SVIS1eXU/wtujWpAdPyMB/vIP4rWXM8Jk7h0weUwt+VgMj4caDJh7PrFdcdFvHbbMWBxM
dddA9JD9Q8hZ2x4zii48V1W63btmbEPoA1meJcbvSnp9YhX+Uqm42kDVkKXOkfjlSuhUwaniSxmu
f/oEAAss/gQzKvePKIuKom8D5c0K4jyiDlEXsgDB4t56rEwEh5FpRkOFruUWFFD7Va0qZnqvC4Rh
uEuk+TGEM69rA88CPLJ2CCSU42dGCJFadmEMvdfDJCgDH71VQI6zVuus9Loh7Gc7PBVkugeKm5Bs
1MVH1ES+TFcyPVAXPqm/m3k+Ic0Y//Yw5B5g+tfFGYjnUEe6g75qvO5SloyofIZFne2QjFuTy8tu
d3tgVQz5w3SGxHmabnMXBlpGkI/mcYQ/r2JZLZbXP9z3SWct1pES9oyjLKQAwlEg/faa308bDyNB
yl0ptg+5td2xGNwwpPmwSpSHMJ/axQqjYBSGLiY8r888aTS3seGV71A5X9g92L+pHYbBaCFp5j2i
+PQ2eCl4iRYlsnF8tn7DpOUPeoa6YNKwcvrTIA5tm6BMmS/g1Cmqe++GUO97cZl5WvUkO4LxYdW5
BEFJYkZAX524c54wt+oFIGqvBdu5vW5v65eqXsbkq+VStX8tUuEJQK2RLPUynlB22tf5bqbQGy8I
brcoiTTG+JFeKsL5LEthtga/zNpaIUq8AX6TPx3ZAqDvJOqTArMB8nO4YdXLQ5r1b2K4onuvD0nW
pU5wCgofzEO0SdzV0+92kyJXB0NlikfWHXiXJrN4P6lN7FsBs0sh3+uyLvtT5fd9Nxy+A3Y+ZCc9
9CFaZ9tVwvtnGHigEt/y/+3lK3FtVO0L6bi2tMpBNcrusN1su7SBBemzspmO3rbKxXs7wCw2SS6z
blb4zmMDGzeEPTiZ6lZ7eVJV04cSrZAI/srzrRsSE4hMP5ADoDvnpE0m05LjbgYyWgE/VqYbMYtD
E+MtHr0cdOtlOIiGnGcm5rP4i0d5eqdPo+GnXU22vIbI59Kt3GBiD87ZKl7tkWEJdDJkThko8aRx
S2YIXSlQC3d/eD2DSL507SPvVYXjnLEZFADk7yJLptyXOqPcdI6GcE4TyWMjbenUmbXSu06dT9lk
u6JfcB8/QjKOnt3ERjfMiS91gxOkrgw3HMi9InI8SiAsnfhlQmPZ0k4J6hem+WXpu2YrjJE/eK8i
it8ynT4aNaePYgM972x8OXStCDJv82Jx5MyENv8qEB0mca9iEDp/TUK7VvdEFYZ+hZI6MclFHUq1
UFhWWo4u5n/rqdX5eC2yqUdHgRdDxa3QVyJ6vih+BFDj/Nahrjhe/HPBakF2VEzOmF2ASK0Et/X1
p/cEsu2BVtqTsfJO3o3hss1XhikKdhf7ttnnxnFebhsqPFJwfOaMv7o9dtEIs19YhVOlZFsHyLzo
zPd3dnzAVh4dA4RsCnYNPCOkHpz9VTGEUDgLJ6Z3q4L8qRwyQSzdE0lqNzSA42+XTzC/xreq+ZVw
y57nF/Blw9L1mpj80AVoeZhObP9ffckASnrECGeL5zd218yV2+CfmP8/Ig8uTboKyeioH39HQnNU
WGbAt82VFS1PCOXQD9Ktv6yAMI9K65RnXDouM22bX4OvrjOyWIYicaxvJbJx1AP8kdCGK7kLrl/4
SeiC9WjyaMstZEQPFiCy/nGMOXXxLdC/bROpTSPPscSkaWepx2fu71oguoKiPj+Mx6X2SjbIerMp
CWGi5nnbKIk4+MQLMYrQbeJsjRx4jc592V/qjHhWf5OjMIPS/TfNhpYsHMalbwvm2wfGHrcz2zWq
kI8r3Kq5roWR+OFna5RIIRon0s1zkrPwvoVHG20/zhYsBbVfeXNDeFIJw84uiee4VBUtVpR0GkgQ
JyPBpX0cEJ26b5ASR70FEaFd6B94S6dlUGQjNjiEn4WsaJxSFUhb+ql+uiIWOEcFmRiTubYxYkIY
Whu1ipXoZZvxqZmYILqBoRzTsjZdz9kBIq2gp5U4O/MXkjGeZKW8U+LeMlKFmL0nHHXYc0hgVEzi
10mtHKk3yxFFSYkW4cTLxRasqXEUhJkdiR3f0RqXEQtDSfAtOBkTV0liuRNWThr96fk+Yb92HktL
RrZzmxdinK1wLNKLAHbvaP3LYa+M6P8kPCoaRScmlSQBIuQgXQv6oZrmC9RvA3fP9rMRFcgJvcuC
Mcrqt66dxXBFHpjoqPR5QSWCgwOOFon6vpDqpPAj//ohpmFyaPzVIuGie0BgEPk9n3MDSZjYJ9/D
VtHUb5ikzOFqJdtMsMYC7Pp6t0nHX8MerE4lTtIF0ks/rYfFE15bGmTcjYyBLfxmQ7m/sibBkcL1
f5GatV8jBM7t7OkdXBj/6IJwTb3+AEqdVsSkf6hA+qXkoVbP6kPpI7++z8VWfpbgGzZqQGM6TX7h
ZiA9Ez/vL625Ak/fDzHa6Y+U9vR5lK6sqPtIJi/sTz1GZd/QQUbz+ZT6DbN6oix9BIMR/5QvPEAq
ZHBqY0B2Nl3FCoHyXxcOFmU0QyHbTVdVOJPV9yWub+Ikse6szNn0Ovus3TUI3LxmybPTPgxEAAXy
HEhyo8lMrE1hV8WFJEq38fLydp9u23BMtpfBUNkJILRts4FkTezLRlzw4uF7wzDNumW9Jq9vtR3O
Cl5ZtxmERnytXZn63ZbFi2+UFtvcqoSoa4ekpupXnKEtUMUCZ9ygnzklkSP9BS0XKwEpo5X173d1
4qPtFBCgjzVP+Qo5YA9SFcjRn29/RTPJe74CD4lpJlJIaFkLHSal7hcZnGpqR2SkwEdjqqV88M43
K8S9v7Hh/KjAVPjNKpgtEJx1da3fZ+/s2BEguPBNsbiMQxy+fU80dgd9BLr+AOXJ7R3PKsDjt6oQ
L5t7n9jFNJXSW8ZUZJEnPAusGMgTh3mzB3YjtS5dN38wq+v4VethUrbRq+2xL/Q6/hJMDacXPBzV
M0IY+m5RoVFEzYiN4xXZXGL+dcLQVGJeMJqTivORxZYgQ04rwlLCp2ZVUcS3Xj8cwOgoQkBt7gkw
PmxAdtFcHSKHgeLosjOP+yPVbas4Vn2/lXhwgFz3PAou2GDMDMJFl9Ijq07ZkDAAuI6Su14tNKHH
YJsX8NA+PI+7iZ+AEGJJP3CxbXT5UuxUIznJHGEAhJclRH0Y924HUZWFVo0GTsnmLENdkQwyuUc4
1AERXqervOXQxivnZJV3jZ1ZySccEbdJ9KfTxxX8YYmp/959xFHV4GanpRDlSjvBRMQ/kbHJ7hW6
BaXIdfOM3BiCaAFYLuDA8X2qp962ntANBZevXIGxWRXmKFLY6KlWjA7FrEIvq0h3YSvsCbbgJqV5
REBo4uNH092rljsbdUoNGMlhrsBtHOMDAlMlfInLbyNENV9Fn17mVhmUJQsiqpewOyNSOryfAXrc
VqHA1Q1X+KZ6/w1LJvowxOEI1S1vhpZQQF0RUOIMuB1FM7dNsRpZ9vHWJhd0SiFwMU7dS6rxO0hy
awiMUCO35zZn6aovCNpAqZvel0o0RT7nsGPdKaaYAIJDeS0tH30CkzDniiKpwFYDdtzuQUp0A+m8
ittqigHM33a6sa5T6t0CHAUhUeZzQFpkotCQskXfGacKT2tgjOXAgTJcGzAnh2zttgnrBPa3VwwT
9Uj5baFLg+3+uQ+aYAmMziqXzAzDeUolo29/0tTecmD2uYyOAP2SlMi3L9sCWqX2+9/e3jxj857J
KHspJHcSseOHySfyWYv9L0pOXtNRG/wwMd2X//W3u75SZ6kMOhPgegFxY3yTAGOVqhUPwpbEil1f
mJDNdbc4qLWJ8ERH0S6EkiKmijmirnUi5T89s9lRgxGVeaOVLAt0QGLD6k/+P7nqnsNMZpHGXJSA
h4gJu1le+oMSWgsO0MbQxE0Z2v2r2Dgoyd04ZD/kFCJU1wCISFSNs9QBo/MNwUnwicREGRk0N6ff
+o8ty13fAEgKcrAitypYAbfKiLeOyU6WEPjQnbXGRa+Ron3xKhRykatominJjLS36RBXF3Q8vMzK
eoU3zJ2P/BmxI3kF0315pyf+cL750ti3X6Mh0ray9Lo/xkiVxQDhF129YCseemHd0gmOwKUxiJ3m
RZmnXDmvOMrP+Q4XXAYdwEw7wxACS4w7WR/l/jvHVkCHLuroy68MzkvE3ShI98a5w6lqOX7mUrov
Gmgo6ZLfYqjV1HuV1lRDjUAuLrAEO2djIxib3wm6ib0Vs8ZIqDdZ0UdQ5phsvyHbJKRmSsBzS167
f2S2LejunzJn46fWyNT6sufyaigvYwB8AGxnhOLBr4VBxMQecQS0Rg76fDxXH2HrIHUUkbHClP52
QRiFcBCc/fEbKo/DOskgp4Pluc3zwzEbPG40IFQr0uJfKY4DwdltknuLMNh/VHCS97jhJNEcD6Ux
QiNrqIJWRnE6FmVVfcZxxtZLNRvP3CaV3VtvxR1IikglNUnQ4GlH8tJc+8r/0plNJajiSNJGxe1V
T1o1lcbhNZqyJvwwWfxF0KpPKTE8WB2bOev1m7/3EgUnddYVbJxmk8KS5IozoFjOpIBHVW8J7q2G
7gzmcWZvIbb1H295SnFrBIwSA/7eHibuLJhNirxTZW6LPnnbdeqjDSxnwN8zYzeS1QO+Vg7qYrqj
q4KZ2jlQWKvBK80Z3p9YlVL+82x4dzUFwjvTLchTjI0sw9E3kB1YxMuxg+XfACoPhr+RBXkC/xAG
DQnBSSeoUP3Z0x/xllYqs6yY2f8TG+hd+MMIB9n1ONI0s8zUVY0fKvXgphaqsit/LaKXYmgv1RZ/
60ZpP1Ctpfp3715FLWisyFRPZceNf9do9169mcGj4l0n6G9e4c+bD0ZjyERiWqSwqMvhoBOkGSri
DUjIbfrJJKFkI2CY8cV6IL8N9nGLH8JOy4VFl/To/FtSeh6/8oHGaYbgdNaCs68Pc+Dp2YprveIc
pr+BHAW1jNsEk4AGd87JcZZDNShW6XSpQ4E=
`protect end_protected
