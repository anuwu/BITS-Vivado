`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mCTsLEbsPZ2vQwU8/7gCUSK/pChAk9a06Ca2pzXOPgWuyZNUN2/38IFSH3fobTOXCRoicKPjw/zS
U5JdUhkrLw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GFPI7s4C1t7CtVyK1SFEMXCUuPDr0XM3dS0SXtjjql05Q6JUKrxMZaM7re8CPIaDa54K1WYrSiji
LOfE418BW3NruEHp6g4ffIGVmqD/6oXHlSP/+pZ+GD8J3ZZ9gHEnk9BLpUeWxtZunteh6jCktwBR
rDRNRE7evKc0RdE4Dzg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sEab41ij0Mmj3TOzy5LUFbrA1DGo6sn7RpcTh4zIXnxchi7xaGXTH4JkUR4ERWmrZubZVNuDty3G
4TW7X1eXkIYL0g3rTl1BN/pYJcBojhcX71F3LLIf2z50xQX6C59oMYwkdcd0PKmDVIlUkuP55LXc
ILCABg2L8H6UmzHAHUiOb/o2/XfUUvzZHBTzPfY1N5j5wGyuLLxHjbTs22mz7su4SFA4cDz1ALYw
WqIXTEkTzRpnoV5wAq1v0Vljr91e3XWzZQtWtVlINSogSOqFkFryC5Sn6XgFKHe60XmBBtCyjXg/
RpESrybcLJXn3Sff/R8O4K5MV88ExUrcKlwcbw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kVMOfbqeAFbRG9AMrD5M+safOIxNtaCf7vbQo4khE4OGfju8gRGpKeH/RBfeF976g2hwQ3yb68+C
IHXa4Ggqv86YT+lK0cUiptCFUEliyQqLgeutmo8QT+myFuhOCigkd3gO/Ts/HA9efV1h3pF/80pX
hqDlXlXuHo+cqoUwCS3vdZF3BKdibV6EHy4qF/qVnECMkrspJXIVcIRc9rRy1y+MbXqEbUCxtwrJ
rm0ZY0xzh+LekunkI6e2PVdvd0g/qtccEy7f06N3TOMMZaWTSw0x9HhMloWl2ouB1S+bvFs9Yagk
Tc5aSMQNzOW5qRZ1mF48mVKRrN1rrE5D2xD5JA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U4bopG4wSqgAQnZxL2fp0S7FrDx75jbl15bXkH2mvALsB9XQUE3qdDMI92sWWRV/uzMbbqIMshjl
ZKIENZsOxjaoJ0hVcroFjOxph6nTzkmbbFkmudkJ8slcjH+xiD9RfeQFHMsXkBGLzC11PVdamyZ0
P7LdruCjryCHGCn70pBIZuh55AEoIPKbMJ9MaIkCgo37fZfwGMHUIfcvU4aDBBuf41xMf2m++S9u
RR2xaqwnsNdfcKXb+gT0yVDNqNasrMWc3PwHJvsNiY4RwM7ZSITnu8GWNRuKRlIjuYg7t9pIPzTe
eHl0DoLjHR6lVlHoVbpqWfaaUa6luuIc7u4PNQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sAs2oWs8lBD4xeSCwEijiqMelKmseqrG/zdMgpoP/wZ8fFRCLUax7WNKGlE6cPnL+y3jaA/+0fhV
ndzyEbMbXXM0aG4qQzxDsJw+4KnEUAFIV17eRWZk6dOo5MnkmDxgjZixEnxP2MzFUchitx7IleaH
iKm7b7mAy39oUY8fSx4=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eWM7fRAz99edtylcrw22vOsawXtWPeHz6UHdrRNJFlHrb+PoOiaxgGrcbYNHn9NMpDY2KUERUmu5
7u8qEumSCoU2dkcWNPpMNn9MGhIh1nzl4RJ01/o0OfiS5LtyOXkCQkzbuE2yNIPRfiygQYgD8Q+d
oGEZN/9d0Ds57Pkj3hNfGS1iNbu/7qlhcXQhcUh203/GNMxjzFCRCWCrG3EQCNAUSPsy+sebZDxg
X72jBoFo8D3NZ3K0TK/OR6j0cYLSAEvX3AUz7+0LifAWGDopG+i3152NkVbQICrPt5Wb1h01Eyfu
TVCmOrE3siGLwl6+yYH9uKwyU4tc9mQHm817lA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oDZ/HLJGYC65wGItiCMl8rUIIcjy2vdrgFYPPFItMXWLV/RCwZ+IAOrpA0FarBzttgv8oSNmKzjB
mNYdICjl0hImxNi9hHbN83CfIYqybRISD/cmAcL4S+aHECMc8R+FMJz0l2qphfvF8mdgxnGjc8zc
y+aB/1Db4HQH4XHiUY9nsNK7nnkaV/RdE6XIclPHqukKyLX8Tq2w/kKoBWOoWSSkG4uOC4SeEJOs
u8U6ALcCaYIStFeSuXNGAZmJ47B22XlipvApuzKJqQNsbeg5KOvWKnof/xMzPFgiqYJalJox6y/i
wpZarOwj/eINR6KiLV0yzqadWxDE9ReUY5agEg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133280)
`protect data_block
XLcDkdIVDeccJnN84nzMw7DVnWYROIn65OVr2Q/U0HFzj9EmZEmXbKeWgGv910agobtA1Wcl4BM3
urvD41OEJxR9f4EI8iJa+wS8xJcFkL2gJ0gD7tjyOrXbY1whlYt2ZvCxC6Uov9h32tRsWLoof4sd
a2h4J1u+rQq6Z4qVw27TfCy9uQaHJ5KG3T/vHIQrajtOb/rHjtQWpA86th3g2IeS8+z/wAW+WAsL
wgAG0in8ydsN6Si5bdYda7J7Rv0pn7/BnTF8FAFMZNJ8ACEHx0hsSYSiyxM2I77TldqBiGZ0MEQI
NvGP6r1eE2WWSnwO9lPN9I6l/N+E1sIS3BDEEt6YpF+G9pRjUc92su9kg2lnIf3nj+QOdije/zep
+4FdA5WKpvIg7MErgeVysB714Uf6f4Oh4mHSdg0BieStuMq1VZuNtYzy6FK8zjcuH5J1Mz2Tzt3Q
5B5pvnxE1dp192/KTJL80JEBrX9og2MV5eiyl6RBhdPl88Sd6jdFT5AlH2kjGbvg0qaQLzAVsdNh
qMmeSSMV7DnV1/RyUlYd0u987QVnLSpu4/JP8cxW9L4dXwwpeltUD0pUfpi//zD8h85iPWlEaAKA
pWmvF7kBexkvWbCj9wLi1dlf04QDBPkhyCK6JK3PEWX4J8eZbF4TcSfnHFY3Ywq+vHO71G9owr1c
Cm9Gyrh9gUjPAGAqICcm1txHdxTv2wB7pSempBJO03RYJx97bihWKLjmy2C8F7hMQpRdExhWrk5Z
MWc41u2DEqnwoAQUv7gwgYMOX73z5/h51JfNMOg2nBjnW0H2o8Xnjd+PAM6mVBtdASwC0Fh05dRq
QqfHq0MDacbT7F4JkW7dogOAOT0U+F24s8Y/UouzEmHYQY+ptp1UTG0NKoEiX7JiRT+ELEbXPGFo
E7xtjlgoQ3RHWNzZFZAJHkBfBG+z/v9h7ShFBwsW/88h9bBm3DPZ2sTtzIiJNuuyQLEaWU+0CDsG
dMVqqsKhAOzW1nHG0EH9vG5Ks4V0vb4GNQjhTK15mJ+Bb/XpaqQo+PkqJkPeuZoAYO8BsphOYwve
KTgyW1S3s4HsydQsvNMZ2X5z3UkkabmcLrEe5RSQi2n6AwwMpoMHqNGV/7WM6Hpkef2vYJQ5jJ9P
blmho1FVzYM3hLsM8aiE3rkole/7JrGaspuXrurSMX6cwVHlyschC5ZPc56SdS6hpTOVfvqJAi6R
d3C/PYi6k6Z32jWYx5Ym5wQ0gyusJXyBeEf3+NKO2uCSUAn+daditnqeLUj40Snc77bxxDrjQEW7
xtebVh3g4CQmuQI3t0kUqn8/P2d+0kB9OFiu78HZwk9vSEJacSgYgLo6wSbZRrIRckSujHcKkQmU
9VnBlRoG2g4s7MMVQ+aq2MGgIYCJHdygpzxSw0On0TrheFs8Xrb/sjGrctMk8aFRYLHhL9SuDv9V
b2dW/io2u7RSREf7UqbG/sKE0AI3naIL971Xt6UDM+IOMQknY/GfQgYk3Aw4R2AyqTrsDiRt2Npe
K8269gQBBP4zxyft2dIo8kOhHStMcMfWxDKEIAeShUp5CHBLTAOepvkc1ecubVQnLX6Ix9Xt+QCh
PLqFfcMIfK3wsO3aIc+M2G8E+a7jfDQgDNq7/7xxQxHdulyndTbm+PLus6C+M3qCROKTuP32JJNF
v7nc8iI9EScNvFByYOByapxO/oEi15UyHGE7iLmfwceWi6RbpC8tm0Q4kBf6GvVN5gW9uTzE4Lzs
yT1Xr23Kx5tNKG9nkKaUyNgF1LKH4yRuWJPjR1986DkBVUzNe5w4eVxWPvPriReNd6qOLt2vaEY+
1k/6KL293fG8FBg17318CU3qsl48FjmYAuy63NwaJgK4UCfGwwP+HL0kdW+FfebnUzZ5Bh0QYA++
tk3WIaQ9VvfaOzgY3PlmPI4PsTvXoMJjAXXUOC6zCcKaXccEf4jTHIBWfPcu0ao9pJ0hEOmms3/a
C837eAt6xGTw7b18h8qY87wSoWwgahcjJWnRFszwKVMX9EmyIqLw5Z7nJJDdxkfjh4s9BnIcTZI4
ZwdDqD8iw3/8R7HUe8Y552f/2Wya4PwpuvEQSo8l+j0ELdDdM8zJGjhwSplcx8m3RFXWrFOUyK+K
c+9HjM/YP5yCDrAEVbKuRubwnnQbmc4z0auf2zre6jO1rlVn8VwYf3lpAc7EkoOUhVCjkFU6h6Y/
ptMrA9hY6LYLdlgryApEq7dV0GxMY9aso1ikNYekBlNeMzPdAHqz9mApBrnktA7eU6KG2UyV2yiy
VxSYG1XIC1jagJUMsJVJou06yzajr/4BMuiSqPHp143wIu1DKs0OXnobId94gGi+WjncR0DFe+vz
MF+s+w2z8AIpO1fcLyZ4aI+ftHapkwdF7FiuX8LvXD1KYlH1kw2aF5tejHVmjHq64ABr7k6P/GEZ
Dz7VlwJ9QzGDk+5GzK0j25Q5ZkqSvdA0jv4+gdfvSYkM7tRNztN64tMD2ptcZLi7g9zw8kBDW9f5
vW/5Yot/gL45RpJEXmmCGb8/L7sSXcJ5o3zk2AAfHJsmgWSVUye1KtqvEAeAqXq+Nvn1kD9iHdxV
w+a3qAE8zDQQzIlkggmMOlvAMOpN/VhovsYI8re4LMf+JQDQK0LRdl9qrZK2uZzRoxaItMGC33Sa
UHNeUT5vMHSb676idQgRGt7x0qtFY0iFVf76qxVyJsr+GqgXkdGKtnZxnYxeMAlVDM7JWIRPwQSM
6V2ciTmtEuBbtdUYkE9YJJcrHmAxFaWyhKEFCOZuHJNtAiLJ6bsMCgMTQ8p/76feocrvheESi0E8
PYVdGzbrWw3iKBNTi330Y3fDkjM6Hw3PrsymVwLRmZMLwdTn4oqjnJRmEG3d39GoIPn5A5nU+c5H
qJ5Np8hIprb0LGVHQJ/LVH0l9xfDD+dniO1G84wGGqIPkSDihA0AY74dYBsky5IN4Ck1z9ZLu4Lj
0UB11GVcJIqf6cHODmr8G9tEOG1JJV9u8Tdi6AmfPOzytWfvkmGEikYr3+npYZ5XHSdm1xxpXorA
wXq1LPZfBtiy2FW5k9KV+wFUogHDc1WLgzOPI5OPocYlximpf4xgDtZCKsjnYiHmsu6dcg4MF/pj
cW1XUe+5WZwWCaa6E6dS4e73DBQb+UggrB0Y5wW5/xL7Hoc1Z9AsqoaQ9rCsNKGj59CM4rd6F0Av
v5w39SOk4XU9AQDGKhstJnYMyCETD/7Es9BPyQu8Ccsonq8bOjUAzzJWjDraRdbefXwhrUe0/EIT
Wwr4AUPnuCfOTgFabZT/9CeaIUmQ7clqAes16GUdaBNPkjJufE1fmxnQkE+P49I7JK0oTGR2inlA
ficxWM+7L07/9149JAc2trtTnh69SBs8dHq4pDwLSP1cNdznWmxVRbX4oHX2L5ZSqD5sDOG8uF0p
UdqQokXyBHRNPi4Gxn1R9gveDrqvVyBYL4h1M3j34OCmvqYGV5esNf/VfiQN+NrBtVdt2ZsfhWY8
8yWy9kNT/Qv7TtGG+eQLzcWk9Wxwhh9I9+dYMO6vsHs9spKiD5yLS1WtLAhYLSAeEivHzJqKJtRa
p/85D5lgKX+yUx9wyZoePVKKy+T08Dv2nNSXx+9nX85Iwf/6SkApjmM4fD8dYgz8ovc6dVz67DNq
CFH3v2wuzBz870IIOlt6ghgyN3tWG933Hj57BYg0ZOjHaOIOQYRZewWKYMwNPRu/RH46uhHeR2ob
O8HW+sp3qXNwotsAvGs2lPTBkK4SRohZ1vh4AbL9lln1KTclnPX285A0riFBkCibK2Q7rgY/p7kG
MD0cuw3/vLWeqJf9UhmnkYqr8NCwvwJbv3NKAFI25d9/0Wi4rSr2eJMwfEWxTUDYk4yPgJiSln/Q
hh3Wt/l1jaxut5GmNdq7pjVrsXuQoVpJ5wmW/UeGyBp6gTVPa1D0pqVAVAttSZKYWBNFjxBzBJGR
9gY4p3TUd8FXCfhRWqV809NxEQ3Vv0K/gEDnaUo5MdSkH0nYg71+3sVTB4hk7UxmT2eIkSirHA1k
MMMbqiCuOg+xIh5pcu1drAoGbwPxGZlU4h+1Ug0qUdU5QamOgS/9hyamXhjiYxOuNLps3acn4ZGX
TNUI9vIWO9zJW+N1Va6d6g+bqjzXkcXG9Zdk18HbUBhfrfFB75tobZ6KvTpvOpaDoVCSfkEoCzaL
V0UEF9Ee/S6tEa+qz0NekFyWzSI19+n5ntScDG/OrLOHinPu0otrQsRVgPphKVdqcI4QlFBiCUmf
DENCkyzi/ENR1xKwk8SLZEi0EyvYFzN+loY5nNvmrK/LSn6weZGv1EUSfoIraOyw41nv921lAyEx
JbXR5LNUBC1BtW1DCQZQDQjaQL1BMBL7la7O8PtMlyx6BXDCIjFXhOZEFqgoMwlbJX0XxBwlz/g1
1yk7j2BfM0iJrw0C7eA+2LuC2xnw906WEebH28DyiGka0Owj4ULxIiIaaDYNVJoKpXz6CwAOxb68
UI8UplBGFNJ0+mIGoe8IIO8Zw7AtmfRnh/hvpRENT7JgI1sjKrYKgORCoHsXtVyNVpkzOxqQD+G7
m1G4f9clMPv7uuOWlBkOWKPbJmcYozaJdvC1oyrxhiP2IzE0Q+8v1BmWHcU5d9E1fW3ilvUDoO77
zUBIUohBUHOJ0Li97J1wFI4b3Bn91Equ/Z3QHBPda2h7cd1oAQIrNTYkkDj8+CsrUVF3N/Zvo45a
O27Nwtgbr/cvNvxMfD9oBqcp0DCGa6MYXuSa6mafQLtSeGydkvq9wQU8h6WzFEEHVw8+9e3ofUbN
2m/HhNvDjsW2Db+TIm7l6Hpo2yoG2BZhZKApAc2OsLzoepSKFWUjqb4X/w3CUkOMklLxR4KYlGXy
DKqN8AYlN4LOQ3fGzRhg2KVfnJKKMISnKt9Jv+4WKF2MUo3Y7LIKCZaOI0BzSNh9sQi+9aMYEm33
ytQeVMHkHOHxViHX6rkfprn8CxgrbeRJPFAnWzfieGf6gnDFtpiAlYcDZ6FnZ6QBSdry9vyZJvoE
1YPESMmZPv3SvHZ/esmBoCSuDgHn3MH6SLAUC2C5tECKTIjZ2UTujceFWtfqufBZDver7avXIiEm
mMHmGrsyi69mMrEvSB+BJ6nvOw2eUh+zqzQyNjkw5PWURuVioAXF1RVn3k0Sq0kSYeBoQOnyunXU
RavhK0uWg69jDeaaekQ7+XqAGfBXIE9v9RUYgnxKKXgyB3e1umze457igRePKK8VP2nWOtcXa81P
KtLcl5P7vdVl1qtUwxeIaa+MYUOHkdvn+sgraNB2T1RzXFqoUD0AGItQ0z5MI3hLjllj2BYHwDoz
gpLESpDAU66MCqVaJ/LLqJ3zoxhWEMBIN/CDnGXYmszJ6+nnGYheKLPzL6FQT526d0QTwnVgXMo8
vN/RQ/1M/1LuSlUmsA31ai82FW+KdRHhpaAIYzqJ1kjNzXYPjgG0CHz8S5Jnvg2ZC5Sn8OusvzEe
TRv2GDLUgUsB60lFABx/ZGVEF/4ccH4LYcxyU63GQSb9sSZxOqy8bM30pvSIeOOHF7Iz+dTFsqv1
WkFpTnNJ/2Nct208OIEQBr72oX89xz0o/7cLhCFEqGoOT0ImHArQJzUuL8JAJOGcneIqmdp/Qs+L
mV82KwY5Th4ATe7vJnmuHYu6JyvDnn89+wndGONv1QriYOY6Mnw8uV93/ATr+rmpQUrOkyn/sj6X
/zzz8MtETJobU1yBL/HoXm8Pv1JT5n9plmgnokWeeOr2VoVO6R/XAA7Qc9T++qae6vabc0KClLiQ
HqNMZc3PeGNDcbVWwlJb8MjR43MDZ9lUI/P0RKG5TWgVRm/3//1DvhpRrJ/yCIhMgsM5vqRWWc1c
cF5yLrY2UD+24MCVlQlhRKUP/gBL7aMDcse5aNpYxabiZKjcfoKHM6CsBwDsedkaJLOmdrh6ZxDt
k42BUek9IPyyyFh/Xtp/6sWN4JtNf7MZ6CrgcQ4OdcpoRlxD60tFa7QSDZYLuyAi0v5Q0DvD3Bap
Z4hrWO+CJ9Wvr3rC1hpIVxQWh3Ku8J1WYelcoVQgAY4vN83wVqJ0HXqIv1mv1/+viBf9kTpFFgy0
/ynbrPxL1dOc6Mjvm5JQ5qvjhP2gawOZ5HJLi2ogjV9ohgSKgayrVonIYzQaTnxyPTIEzF38WVN0
2g4DZi4hFAXsYi6nN3UCLhN73u3aNpFX0KGtm6nW6u8WZuSnanu4d4NhO+L8ugQqnF4raqbBCLRF
7OI1pm4Gp+Lbde0pkXSlC/ZhhVIUcd6St1rojXzVhoXFQfz+64z7TJM7OcvW/UXAhwe7fJM6r86D
xKvM+hLbYomlKEq6owUQIyvAhHzbvYWQXc2wohW1aP0RMeGdF0egPuN+WaDfh5PMTsB8dvJASSn3
sPz9gPGTqDUDnKDfoio1FMvclKdMVmMoN3TZq7nFN+mfwCuRt0Z/wWOWeiGlR8Z2dAcK67fkwUE+
itsdNlWthPsrtmjNCMfyc3aWSAUFWWAwLtYyIMteDPKam6sYPh3UF0k43xp1jTdghy1zbX9bLkVW
JsUdMGjOFleVP8gM4n3Yag4us8aTeXowy9asOdd1RLiz2iRv0j3qJeW8KuF4OMztqrb9W92lmhVo
brsYSSuwS90O6w0v9El7kml9gYqusuF2lclIiPpVRjJLICzRQErujd1cS7t36Y+Q82s/ZpfuNq7s
oVeiS1y2Y+uhlDjc8gG1LH7awEk+b5xlToIrG71dLvX4O3lOAQbqTZl5mUDKf0nl5pfDZ5FlwmKV
F4q9wJHD7R9cPPlR+ydpVzhFU/Osy4JBydW8UkcpAW9AXIk6UTYJ0j1LNzK5JsEb3bMTTmq2clxg
hAyawjZ49uylwvjyle44XF9ZTj2ol8xC7f42A1XIzO6ipjYbDv7IOScUYSQ+LR+olV25SJ5BFZQN
11Z5H7r36PfZ6DXfHNh/9r+5NV0AeUdbCL5XFfwzPcKOZRd2BwAUW5uWdp5C0deBdsR7U59hBlI+
lP+UavKrRlVYDHAbJI0r7F050UQKMltuuGZCJ0TNffK9SLi7FMHum8izhelA9E+j1rgSgzLXU3y0
qIt0M0kJ6TN0H1LITXlF9LV66G2R5Q8A6PS0FkRWYJuOoLbuYuyl9GYFtZAH9IckL23bRssLxc9m
RRUb7pqZdn7T5JTXarUtOraWcBgnfqDv78VtdPya9K9O1TUJSIprg3vnMJRosV97Kn9oOg2jfcUG
iyn2r8xEcTUjhBZSN4+U2L1YAnsFtMXKrlo2eeWjoYVxE9q02JwKtTCK/ll73NU9wO9PYdFpvVB/
Xdx7ICKn8Hnz3pwQkQv9Ooya0iw1gpVHzEcgpkfVHThTCtVbMiN5Q5vdhIY/yBSUWmzrYGTFAC3l
GdLNyPvraxLrZtAedXMBmO9N6SeUdt0QVLh0uBy6zTymaULYb/5j26uQRd2RDhMWgfP7f0JnP2Nm
u+BH3iNTgRtzZgez77Ice0VprZfSVwd6t0WQreJ06fkbTe6Momrexm177RSOto62UilEfwQZAIKI
66DzvI47J+zxJzPxcbpkkPcTbwTEyVGOag/YJ5/h4nsEj2v8r60H0aJHVOcuH/PCJYxG2rYxAaxY
U7n2/bGt8ABFqUZRjN5ROAIcv3fwYLAkE9w07Rz8t0iXqo8R8XKKLddXEgyfA7Ti0Q0CHD3kcYyi
mdXtb3R9ofvly9iM5A8zmVaBy9cCULO5UJIeLTZWr0EQP6KFOhvQ59KnpwBWnYG/7KfYMcULgIMT
JLcjs8tDaN1vq/i0Ph/C9aV92fqWtYzSjEsrNJhl2E1BQO4tGaZeWjXj68/Qpg/sxTdv55ZOFMXR
6+42k6CtTzEFkENwvg1mYC7o/o9xhCsbXEuhV5vQtkH15PqKdibYmMeeLEePtqfBhB0RDKV0F2zz
eW6mDRnyI6U52O5dJvQyOeAqCqF4+3wHHpQx0wTi2nYbOfk240gZMdvs4inq3jSJKlu8r9Wcu2yU
PETN19s2Pxgz/SuIhKTUDH39Gn321io83sW23h7vAmUyZogAPt+M5wAb6hTwJ+XggBxs3SneJHx/
NIHSUIT+lreP1fRmVaC6vFE96uj9KmheEEbNq3Go3sSXOl1iknevHVaDX5q5HIX6W9ZQCUF3bywP
mN4vYEKyKhH8wigxaG1f9t7fO3625VR2VUTW4/V+lYj9zLriGaaVnhfSJs+148m5pVKx8TPhGAN+
L5uF5PHJoPMHg6xcIiLhBSKrZ+oS8Zgq1Kb1qqNgnXUn1zD4lPeLUsjSLA4SJGmRZUgXN5neNTNZ
5G9bq2VZnsv8L0BWD8GUtcn5GdTtjua5aBjN1PBLeOoflfaCqo7FKoQrFpC37r9HYT6kq8Y12ZJd
CCXW69TCjleyb4mKjjwXyuOEClKh+1G1B3WJK09ULjB6PllGp1y7+5rn8nHLFiXGT6oyMjJhGkDs
vyrZCohL+J8NHiZ6Mi9X1QYyrpn++f1SYkdirbZ2oqn7GRizOtZpYuV9LlZ0HzxA3A3QF0/kdyKL
K/WyfDujCZ4q0oEAi7ymILaETfsvPskufPw0b4uraJR3+F2i3I9HG/RPM2uRfr3LopeBFcs1JShO
BEUtIvRChNxV4TNJ3+claNoD5EHZUYBtU9uMKugLeFn17Vg0qYI7Q5Un6pTXYy7YnfvH5nk6Shfb
7W9DTXpdqeCo9uwqIGbCtZpnCD2kihpxPN7/SSsg8Y2INypSBLd8gOdRqILQmUh7SyKcIRH4U+VN
CBmRomnsrtNmAb9WU8q7KztnpV/meLetdXZ/HnnSBpkCyOEgfU7qUyAej83wVKGVF3HLNs1szDzx
mC1gOg1KmqbvyAP9mZTHSPcMIir2fyLkg7TekgCfCiYmwzOIr4nvqCWgP4UZAgNd1ewoG1ia0pmv
cFEIvtDojhgOVdeSuRLsPO7E0U49bKAdlusMsPP+RyDCGGvBsxGxVQf4windKn236XWrtU/1mw65
zZp18rs5Y6TvPE49PsU71L7koQF9HyJw+tftof/Cu+2d3qqr85RiM9OMoJ2jXmlRcZhepQVHOvCD
CbAueqPuFZT57pPKf9qPHkiZkcAGHl7O9e9dZpNngq3MUhwk3WneWyb4JSsqiIC0B606S6HWx3oC
5ka0gopEOzFoUQ3MeLeT1+9lE3bQTb1JdozL7RcIGRMINkcb7iLk9nRpo2FroOa16+UH764ca6Eg
Rgun1iKMo0bo4yDUD0BhaiG+5FeDc3pd4RTj3nEycvIWG6hr3l9gIugXv5iDVFxl7/cgCdh6417y
92mHj5nYAauSQaxpoo4M4JIvTtndKaOby2A71Le9vSJHlGqcnZnt007Hzlihv03N8lbvd2JNrJg4
0DiFPdH5a8efmrTHXS3+iRbILiadbprLc0SXPUMTPsjkwjcPN7lHh5j9TumZ+6PQdGGbldPKrH/H
ZMlLmwdgWZwTGehutKM90tuWYjJWQkDNwnEIhNcqH29TCxHjWoPjgyzJx1V7PcCcJjNySHfqdkmr
8HBUpsvQq6m+rBUZ6jMh0qOEtxzVTSxSHJo6Hx6R/2FqFzLmlUEW1CVJuaM7PyT+Ug+p0X0v//hA
F3II/uhvMU5gYLh20Q8EeAPfAdoDU2vZauUDwAl2/gvMzEm4rJsEq9r5kPyD1ed2F8RJ0ALP/ZgZ
PvEj79YrdNpbigNcioJ9tgmwAZ0y7kYLMU0hRJd7ELWKg4RBG4fzyjWNP/j9G0PeZJGArwjmJslF
mxrVPNueGf0igoAQVrS4YxNT/LtkMkCzfDv8a4qDSMAT4qCKFQ3ruyu5DXjdnDWOybggJbOSy/6c
TH+cZqYzG7w+xzMoZJowenqY4Gwhvp5bJQj6K/dIZi23/kCqMFEFBY3S1gegjomPTlTD3mG/FLkl
EhbX49KAgR236wSpJ4LsAxNM4FJnEQob9N22Q02Gd6fyLJ8K8mtzgTMcYONczg9YU5I2H2Iu2od7
JQxKQVrQSHc81APZfktJFe7/BrxqAKb/dcmFZoh14uV8RRj6vlbmpx3WifCx93mpxJLS35J6x3dU
pfxAeO+IxRWC8VsiXQ6mCpFabn/DLs9cFF1MOD1d/b6TxIwY7wgjyCUBhcZFJ7LpjwoGxXtzgtN2
uBduWPNZljx225RFuLnTJVi8UOLtxXDP1Crr1RN/fnVHp62EwfMetq8IUMNhxbw6Y3RMF3MLsSrI
5wu1K7oUpZhEp4PAMgsk8W2n3n6B3w+v/zg3Lh+a93a4jCU724472RBP1iDza3EuAgGx1A8YG5S6
GQRmthu1ryX92V3a9nLleKssY83cKxxZv531ROEpCd7bqGWe3ysdGyy0AcPwvWRMleRkcL+JSY/n
aTKPPBoSGIQ1ECeHzboIlMxP3zp7jOZECSH+K4d7zr+7/6YFpDeLew7Zc46fU+e0Skpx6bukNn1M
tWFXkEMznvq7+CyrqxsJaUFZSXsqrwO/3Cq33WDU3dZfHdaIAgQf7FSQ1kFTlOotEjp+jwhnQXdn
UP30qUpzUkYh7TU6Atqp+/4me5sJ51eGDHgunuQaHL3DDtuHzJJbCcol+hOFJAOaWmujHMqDm1Vy
vj3OJXLRmYw3TFeXUMnINddCJRyTagYDzalc1Ne2mq1ONLgM9ScXUh+ZWmFaJQZdqLIutAg1o0I/
YDCRFVVszezDbXR6VQDhN9GQF4pNyDZ2rKpGExnUOdW8tCX+u3CN9ytWE866CgLR8G1RVI6r5p0U
ITggq/ATGzl8mmlVaGceWzaDeUFRxM9eE0GPumDsL2H8KlZeuVvfsB957FX0iTQrTocUJH6ZvgIS
TEEDzq+cKkcOThJGtf/OHwSWQ+41ko7YhB5j4t6rPrBSzHiKoM9/poy/ktwfjbd1Mw1VLhgn6Kue
pbdxyXRBeWLYfl5L3cPv7GTjdZsB3q+ARRHYwq+AktYp938FYViwuMn7+C0YExZVuNSSBgK7f1vq
8N5P1iaelmL4lQWsV9xRYNzb3UtY4SulmKQZ3kyujG6dTQXRzm6pVZJEr/m0p0hMQoomUL5zus00
Zw1KaucPPkAFuzL9wgyGVAGzwLSr03ij9jRGYUJogpipPW3VQ3oo4hmo1hT7FrN1y0hJpqTVIUQw
2aXZyq8apdIGGzxpsV170UV1FS7H2Ja3mjD87r73IhXsAwmKJzFTpINm9eFeCjmzLtYNTvxHLQYO
92cfR1El2v155nK5a5yn0gDQioFjAZCd/JB2k1pXE4SbRHRZ7CDl62UXm2ruO2VtP47ICU5/guZY
IVyCaTTcdPnS7tYdEr6gbdGpJ7svb3FEEbrRTBvmpTWihwFx9qxEMuRdnyFQ6dTQssKXFBb4k2OZ
xsQXciyNH1jAAB6o8cASVXEgHbhz6cmrwLUOxfg0liWvDEf+3r5TplXITunlD3HA1oLKO9FiZIm8
wX2xBUNbgs4RTOEc/d49oHL4yR4SpleED3rbbmYnDu/nlcEsThIJ5p95JAq6BD2DWCmYYDAzk/VK
66ldY3wCNxxHRt/ppXzDPQK9u0obvFgY0b7M/mJI4U5twjooaTcwTlJG3JA599TpF9/Sc2zEdPPk
Hz+4DH+D9KA5Nk2FZkem/Y3lABQFj6eWIOIZHRb9Ey+5yqLVaGPCKLfeqsAL9kjFJTzIukiXQn8h
0zIqpbf+mFUbcCJTy8T2XNrTTDG/kwxfLoBtfl6zAPEE1zZUZMIitAk6cADIBrKxlTjyms7Jcror
auor/GyLiSB1nTdKFIocgHySfTW3Pubwo7JTMxdK1hEDNoQ0XdgLvgBLBXD4UZ58Vt7MesZutbOQ
IhMUa37sU3W6VGqCPUw3K3hBcahNXhJSufpWOHRZCj/Bm7+Ov+3uMeKZXHT43DurPxu0fEcu8VLv
kL500Rc5FKFCUTD0KJYI+8+wcHCq6jgqIv8se4Z5M6Q7fAjbyRK4pN7oNQ9gMD1TM/fZDToh88s8
sVdqSpNqIYzCsREOD7y3U/vbbGXM+z61prykciz0p/QteyTq/1qyLLQJtT4r1tqYZBVnti3lGR+L
Xyx098HuLt7/3cTuKF6XqbyQt2KqUfV2gyHaaeuHma/w1lUVlvk2FSAsm1ASqrG3BMOtnqNZpOVC
/nh+tP2zXPJghN24OvBlBy/ey4rzqO5OnNM1byJwqQax59eHH8e8ShHO98piHNgCM863M0n8oCsl
pkdCRJXPFEx26/WLZn6M/NQPpFzJSz5nzAHAHkzFFdvVpr+6JnrfjzEbp9Ex9RMHwMHmBXIJf0sz
CUJ8YLwSJ1wEqoHFBtga+l9opzj1wIDjBctYF48YjEL6co7VX4IBgTvFVsjhvqKUsYN13ltAIaOQ
Bs0b28GglYbMNxcbrBqlD/xU+d/rQS5WRdhYzzSJd4kGeCM2BEINgD3ht8VAHKY1L6CE6TcrPc/R
gbAgFCtZnbUyF6gYasasyJbX4E9l9jE4WeaXIUAc73b3jyif3NxpUV1mn/4KED2fi4aDgN3lmw6V
SJoBNJjRIrBqNTRIRnzqyHouPg//r0DX5QV5r1cobwDW6MGEh70HDbLZCxfqESj0x/0OgEfGznC0
eFFerPjlafY+NijQop0PK/X4ErDisTiKhmhQR2JoDi1u9F/KGUJ2fIY16QeL35fBGYgaFQBlekxA
PZ7+k20Hb7/ixFo6N44jc2ZFylwMKexIvGxdI8gPNjgqwmLbGEcwa3h9YhoxGaZxPXrLuj0Cu05T
MZPX5oJH+cn2bB2ExJLBeqJ1GUi0m1nbo/RqgLRL7SEpVnSyTViuOLk4D5iy/kw/EBfsfrQM+8Qv
CI4PO94HnOiL4vjZ/OHz7j535WtLoolgJINTy+aztFwLCsSo7JGOk/0Y4BGrEyBUgdZYjQC25TWS
RRlUt5yz7iGN40aU8YKT3TCslDFNUTj67iJSC9/TzD81LsfpQQAu9J0YTDQjxVteFoItP7UZZ59q
SHAt2QxyvJlQtBP3vV/FgaMnLITsHhDYolVhBskyMY9x2FNRwCd11qXd8bXZg7X+85jbcOnbGFu0
dViDFwggUz0Ueb+aelWDPMcM+TA0q+VnIoeBJiEyCsGaIvmCTThpcccaWPjUMWE6E+zUdsPq9Apu
0mxLoLIFwNEBn4/pMcnbACsyA1G3J64Ozj+DG5mP22MA7MFqM0C7y1c3PJpyhFIApgMrJ8FJmjKD
azIt6vWOQ4krIY2OQnij2J2m/IuPTsllDJDyNh/kk+/mdV79i9zflQtTJzQ13aBvQD/UVM581/Jc
cr5IHzL53iWtGzbwkxjCjbs5+na5SGhcUNAaZBssAN6jPGQ2V9Os1Qy5JMlqjWIRB1HVxVxQ1YWR
Gs3wCCZzkKum1fjlHP0JzjQi4uXuldzu4s/VSNOUZjK2Jyb6w/E9n8rT6RA0iC3QH1LEP9V+3kjx
QzGv672hA6m0fkIvtu3fjk7DoHp6rFxvZK38QyM1In2U6/aKx/EZ1UNGB7h0peVSlK6vSJXk25eH
zWKguSgb/5cJhmS6jfIwZo3SFSzrx4gkzSrBp3y/XEs8xQrC7RTh4nNApnkEDEtLOHQDOwgufJTZ
AmbWvdpMOR8dGg6CIzIm5ukLhlG25g/7tGP6hNjxkL/dg7DbzajhRRkTtMVW8y5Qux4LChXl03hF
NoCTkXfgwtKW9vQzye6x8DRb1TI9YNLFC4fdoBAN4jY6r7gQ6L47AVGsEgEhps/hqnOMtfN0gPjP
fNP10f6CUENAIHni/xKA5M5lI0Tq/cbloiSn30/abw530g0sz9oS+lD6CveODdKYuA3qLBqeEDYz
/62LsQ5F1A+qRz4L+AyBPF36qWSFgcPyqMzjvyJKfXeAIQFjrBpE9HyhAVaj1QUKjEyTt01+xRKH
AlC3Bhf+iWSjbCj4CaHJDTkcGddeBQbpE/DMWtNVBwi46B34R4aRCUW7iua+mcX37EecioZxMzOU
KRxtWFZCsIR4fCxJSIVQJw6O/4kWx0/DF7xOJZMnKPcGae/1N7m6TwM9V0Btc13ELlIVjsz2ctk4
2S6/2EnD3ESVRXwe824AwNa4+Pu0J6yHMtx1U8TcVmbUIhbbpnt11U81L/yDfuL6O9J/BqN53ErW
Xg+VqlwHUdUKC5u99x3iIM5IQWh/WBxXmPc5ALV0YV6yozZbaPrg9AlGa0FPnNKDrWHDYMzI4jjQ
ykSqIiDzIblK4AaML7XuQmYX6bRQ5AfwM4rfucUpI200nsrnGzP1os3/Raqgc2WGQPuYd6FF2RHv
ieZgpXNGVu5sI0YW23YxkwErvbQngKW4ospFB5zq9kHzq2vllGJmsHX1jMnQaBt60z6py7ehLQUl
mjiZ04jKrdk/3R0TKf1hu5iu+Nooo4EKM10CJQNk9ptyVS/id+fUrR/b9FJGVDthHAfUjHKWCU9W
3AWI/9cdqNxMyX6ShnjNOpLG1pErzZcnbdQRkn4+FBWOv291qFNk6UXInhfL9LUcYP37ZxOfRbWT
Mm3Jv6tu2CPEMzWRIpOiVgmzVOk7pXkTAMQ5/473VbD893lPlPTAkaQEy7wOzkdBNkz1gTcnIkM4
IJM0205O3krv1xI3Ty9V6klaQCJT0i2W1VJxHmFTZOO/UEBIruUeMrCP9R3i/Hv8flul/1Sf/nE6
yv9+QnVAdM/174Lxs8moEfUBZMi2/yfJ4i1NbRzwKeoyL3/25NlCcy49G9LVGlS8tPLGi9nHwApu
gowyhmsdC7i5DeNhW7LxJB4r6NUxYum0eqGuC8J4BILq5KxnH9ylrLqB1d+3VgFtcjzdOO7NixA4
xOsKiXy4TI/wA0weT+oWU3/Dsn3bPbbjJzqVm1B4RKMK1VkjtRH0jRarzaq1upa7S8F5j+PFytk5
IfPSZlNukOQ51+pyz5lyMS3ZSnaK9WG258YxtILHcPYqNtPrII/TUeNTqzLD1Qgr5TcgyUqve0OW
qkEtDcIvcSsqlKeVWfIrZr10jpr8EA1tdreq8pn00xE5q3PxgDLquU3ClEnqsAc/XPbBFUKbO6ti
U0+d1/bLK1grgIEg34m1GYGIOINyaPjD65AI+sIT7JWH2J2vklnJ+aVCKgRx1VmNceKDaK5jjSmS
sjgnQ6a8HFyg2e7d+49IIZv/QjSEuTu2vwHr92VBcVTD4tx8gGRpa7UeVjLFoBKB4xajDw9b1Y4Q
oY+Zyf1hn0iEljHuMMuntL3vyxZWDfUI0ZwZ+DnwWPsxHKtm70CnkcClO8OhtI1SlF6pj8q6m7Lk
WYPeouzNyLlPnwf/mnlD82ViYJO+Ompw+NCGHiw4zaE5iY13LGtekjUhIDm2T4iik6xOsZciuBpe
gXS1xr2FQqnZE4MUZ46dPD/urlKwW1CvQWrr6KgOZYaIfrb3FMOTGIb0CraSxenfAte/4Sv70hJ+
WGF4+dG9fVXE63DPtQiKp0w13KOBEvroL9tlQwEcndMKeE/S5iepS02atd4uOugcDATu2oLRGUHy
5yiD7+zDHhY8Chptu54nNz2FMUamjyyFEH+5gSX4ERNKx6O7/+sJoY9wbid96T7Y330NGwULXKgx
Vr46nd2oqJ5fNpX5fNjSl4nKXAM4Tm02DkIophBAr6a74nCstjZhZ2/xTjsOIjkRQ+G4kR16ZN9l
6ZsNca1jKNsuew1KRKBZsMLyD8R5In3d6Wf1hhdmYC5sjThdo8FhS02l1nZtsJPoJCbYabsY/Z5U
T5bUW/yqokZxbixyGbCE/lyiY2Xm/50souQM/ePo5/r3bIwAvsOUfCpXoZGZQ1dUpdHGT822SgwS
UbKLmBg6rcP7DD7OMtfCkdgN/Unqjyk2UUqIlkXZRv6ULaP/YECoTPFNoMW9CGf2FDtRQkOxOrrF
AF/4m6/1e4rLdD+y8DDdJf3Na7SoHyrVFiTBanzS3bMxWS4ck0xYcyxKRaVqSgNrPORKE+ZAPZ0B
KHeKffMuybtmS+CItjsC7tUOJMa4BZtNpW9PWJjU+LKXPJ9yQWtoTByM3y053GVTuPweGInzD1SD
5hFHvbWEnNvLre4dWsP4k8NnASnH/NRAQaUEV+u2NiCeFA1CJktQ5R0SHwRy87ItLC5AUycSIxUZ
LL9iWxm/nfqMUvc7XlZaTXe9Viy9fPZXuJ6eGA0G3TaP9LZ3W0IeqypvAXk0bYK+ncw0oG7v6kf8
aLA2wlVTWGFVzMjCcXteBmQJ2aeXScCNT9phZt85jClSRh0DS/Fkq/fmFT/l8ut//FW4oxg9ivFh
6BT7zbw/Vo1faRhyx7KpW0tNbRB9VsZSO+as+8blAI0pyr1nRpzyNtyIbobmHXymnbshYMIcVNCN
7TB/0U/3xaaNxVcRBVZTqvMBCBIQlqxDGE5nktsqjoxsgszGeQv0f5+FapDXkVaoWAsn944K57Lh
pT6Hret/y0+EmOi6bYdY5zIX6I33OOXFoMp48ETKpmgSGSZ2vaA2JKUtnlhRdOtbkgRs+nT4QULc
+weoFwlRuri1zKi67tAERXSrE7MovVqdIRo6M3BHyfukNQqbxy7EUvF2ZchyxB7SbuispzaF56TV
LH2dBuo7zOTKsbLZSXtLiMxXD8hV+BK5EBaZWuswRz+IzQ56HjmRihQGcve/9KWIJIAB/6LRtWdn
BvY84lHWoR71UQDCqNqS8Vm/4i7l8pOLeGv3K/ibfYSQuMaRNVs3ne43NQTpgMAAU8RaOEhR9ygB
xu37Pw+QR6hzUzvpNrAC9jgYgJNN6Cru/N5Ow28lhf72AzeogXc+u9jakBCyXLSrBjWeWE6CeXtj
dAXFl4ILSNtNpMpQeKH+8yV+RDOahzyUQGcKWRb/V1UbRYRBy3QRGao1htPq3EnCl7hE2O5T4rwx
6efQKL8rssiSkkhcB37m7kmZWvvCn5n+VH9/lBFSqxK55iUiVN7a69jdtpxCenEUX09KHOMpc6F7
+8TM6qNFKxSiDjTYM/AiMfuVL/rW/jNj90+hJMelfaAlLsKXgqcESVsAphjxxS8qcuy9ifGio/PF
48U+PVIHOGDwXi3goffnJ0xJuASaBLndIN8V+W3t4IKw8acFdpw2XuA8rkCcJsmn64xk+iFwunVz
RCCqZvY+s6DWAf156/mwgsujPVYWg3VRGE3bhxvKqouwI0JjPkeMb8Y+YXAZu6d92s1CLXK0Y1s+
Pdwyqs0vBEaGWbCKgfTOMRvL9d91XqVASeu4SddRsYHLFkiQ+DHwhPL+ehI5qdugSX6PTkwIC3Ma
26dyzJCIE5DnYEZfLGuiIennstS6MF6lUBV6NcryKTD/Mn+goBW5oJ05n10PdMg42sea2Vg4NLV5
DA7Kubbgt7rzhISOOKXZW3MQhCxAZPfCOOZjzXYrL3VG5Uq9AbDYtvX+qzwkjnVhfGlzhLIS80eo
oN0l8zxsSdyFxwEbQAq/OtdL2jHLXVhtG3brbRRNlyxBYH36Wxq5K9k/G049122Hbc0IGTLME0CD
4dpOyVUWlV0dKa9ucNtBEJ65RJGNLthcWp8ui4rHB4B8wHGP4OtxejiO6qfnj3RZQoNVtJILGO9u
e1RK3A5Y3HBX2sUJKOHdQnzui6z7O/avCcG04sVfBPQYJfj0CWc2jvdvlbPUkqRPn5sL9A9LOcTJ
MT1/QJC05t1h1V1WUcir5xUTrHyGbim8VGlqgLAaYkC4YZkxOEV8ICFDVbSlLHds3+5Xxy5pAhV/
j4DW7elapn/YUBwKxVLlrFFPHvM0HIy4i5RnxXseZnc1umesx2G3Q0dlGdgqGr7KcSnr2JG58e+G
/5dadSnYYGQ1hQ8eWrSeSQ+UCpOjyRRBKVoTTAb9ulbu+W59qpm4yZatSVaR1Cgtl6jTkBk7kuX1
V0WrfKIxCixX1C1sL1QyyxMEHTIxwoZ6FStUtmzZ45J8spHyr68+CfMpCvBxW/UK2jQfLLDLE9Ur
H58b8brtkYrdesn0y+7VjWMBZuyslAuSu3+64U9q68aEFHyzHhXf449+kqn+KEqr2R1h+Sa6vdxq
NlXnahuy8TtG8EIcnUemmfYQn6AowyzverOL+ET9WVkq4Ss2AW9i+mlohSgoGl2IQomlbDW61Wk5
1iHUUjuPPFCiM3KIKmT15/bR+XdMSv4wE6HYAmt68ZmXQR0IRMcpcYSeAx+GAgHGcSnvl3VioerV
Sfwq7WY6GsBUcTigWnnvWwkjWwZTpxuBzXHN+odcRd7z4j5cc4NoiOhmRTHtq0nog7onZdbECB1L
9o8GdpOp0iDQ3DfCmjtDm9i1PpNWIIbnvYsXEjpQy6SQl7bCDAuvEX3ikDbErUKHn5Hu8NRPGidT
YggdGt7ecJYcR1Au8T4S7aOMa+gTZ9nCdkeqykkvTHLzsoc73zDMVn1PPEoEjhu7FA+cDtYQfKsh
9A/QfJ6oD5cSrmoNK9wCCcNm2z8dDWH3zJJD+q7UHgLuzTndAEslG7WA0e3P2rQR7PFpddNGMsUj
J9kQyvUvLCG6hnsKRDvWZMDcmQVIYRSkgwHUtHZUbJzfIciVgIhCoAJhlK/WTYlM8jmKwCtSYAk0
wt5uTEqGef8qBm7HyAVrxLPt540MKymT5SDJXJmfdnMgPbaxNBXdvxOTJxRHll3BBRqU0bkGJHsH
mVHdO7wpR0mw27iIRaSAkpE9xI/0qbkuL3abBmFyekRe5B7vt+YNsw3UPQDhvfKaRKhKuAD3TdqF
tF7dY+uyAEr+p4zbZConK/ziyY5eY92llBB37hkwOc7qRY1TN1WIy2Pd8v3/tXTuv1A77qKkrqGG
+fCKGrvR+OOt7M5ZKp/j0SKBbCq9osidv38fKVj+dCMCypsj0ONGcW9kGZ3P258cmHQ7wq3lHVWz
icNR/B9iMxCW9EMKhtbvU/uUDgclK1Cou3qTnoP/0Puqd07L9PNbWdfrM1ZTOrVce+/bFZ7fnQ3O
vA0SXpZ5kCl4X8Mzv9hTOx7c0i6iuVKdJnfHSdVFrDfOvltXti4laCPin7eF/TH2q+W0JfsNjhkH
iBdynIy92B/K5eE7hsf0sMeCwPnyi9HzykTlYKjyeFw0eRGEY9Nw6zQutJI46Qnmwf1w3FB3qelE
p133zmWHJ07J/LR5ve5PkiOoPAidQZBD6BB3ioJVnvma3jEosiQOuH5Kt6Elj5vx0BBSds/Ars5J
Fe60uSJWdy27E+q0Y8tfoIROJ6A8LX/D7ZLXVpU8iqucxp2Sf2lHC07yt38n+CAFvl0xD+tFfQt0
ClxKz3lcrY4G67VyGXTry/HlFN9Va2CpH3SRv51LFDNtHW7Id/x/bu4A1gfPhm57KsN+gkKxtG8y
ANqMkHxalm3NPd/SiITvSsXgzO2guB9t0BZNCgtlsX0yzHOFpal6wMEHU7X0JCEzT/FjFn1knFA0
Of7ccGk9Ir41JuSJ32jgFnXuBZynzphlpLDF7yLKCf8yGatpU7FWAWJHb3io93uytyXV6+0s7C0n
wKddGVtcS7rsabTzFGh+iWYvlu3BEOld56zVdKLUimdcmHkMCJLq/+2Rsxy0dZcQDliX4rgXAP5t
pGK6bpPoAwB+tU1jqS2u+Pa51A+BbG/ZuPuwxgscCao2XRBNLo3Cm9M8D1xwb3fVVdl/xvwLUs/I
O8wYYF3YjYm5qVTMsENwjp45g6F1s7oReeTRHOPwmYHtbaUE5zJLDgblKVGKkc2z/CF2vhpLZu84
6ybrUOsDebeqXmxY4pmKRtbj4sWVgHtOuWduTro0dHq3+6pqpjVe0gFjJPplLB71uCCElgT68O5J
hw2GNC7g31Jgwgk9rgkro35DliL25km2L25Mko8r83lsCMzTXtokw9cY5kkBMU893FFy0d9OkrZ9
06VBKUmX9xRjnu6vjATeS0uJRt6+LChvf7QWNxm0+RHxisWd+rPOS25SJQ0AH8R770Mss2BrnIQg
2fzwXDoDyNvMtnVA85f+XecIMVwuMaS81ciOzl2TB1TrYheBSlcaQrGgBSNJCM6/s3+Ajl3MjeAf
medxDLVtl42klHF9cipxswqGD9VqluUMb5DfIBwG1N2J5SL89YSESRtaODsTJHT9on2ywNsw99dr
WfDbn4HFloHZWGClG7kAXynB41SnGOz2KrFb66AlZQ1ENrfWZuWSBN2/1VB3oWICqWfqSX6jbNHw
b7Vmim4PcJjUD2dpFB7T2VeSEocPdAV7G7CsnelFMPPHRt1OlXRuPuH/tuPUmfw92jp9RGAlVc8Z
FPzIOL7ILcjzTZKj71XpOJGMbYN11uc41XThPdP9pGNzVRKGvTfVhPnOS/3Px4QLdgI9k9Z4E2XO
1XlZ76HtzpW2f0rJORrGS9D9LnS6Q4KD7YQTib4qQxVnXJiujW2QHQTkMjswTQXmsbf7nw0P9SwH
ft8lGpSYujsuvXM7R32cyRjDBnvOkdC/ayTlgPA2YgmH8s45D9TVT/rwky2ziv+sMjmBk3gFFsho
5DTZ6XpEa73DqSuay1o91sYr3efgtHTHgTqvo9eYXCWaTaBlzoBDBfRxIBwpTjPI6sJGTf1U/baI
8dWUZ3D4gOUxRsY8/qo8h5xJsLvnsCkriAluXewJDMHMpoM7OxUi8m59w3DDmu8qSADg/2G5+W9B
UeSSIopxvxZVUCPrvmx9f5EpKUvT+FADkvPwjSlUlBrjnU6ln4sR9oPlrur5cnnrZQIFzw8gBQFw
9nQqilhoYXjTjtWQNcj4XDCWWauf8u0vf7VRWa8Cn+j5DGOJeYLH8B/KHCohh4HoBcPmn48nBh6p
mM2TE90BfxlpMyq5a4i9kK78tGgMneOXeFBvbn+F/7reTyPMagqu3zdVzwgP0V2+YpIJWvF48G2b
KhQKYQO1knKzr+f0mEuiYg+Onu46RB+UAJmAaC4LVh45oXff6oEff96Fc4XxlRFyCwu9+udp0cMY
fxN26RVZge80puLN0eQ1QIPQKBuKX356qc9kBTvTqokUNcTcxh9xqLBG3qM39p7dwquvXrnc+n2z
nsiWH964KqoDnrYYNUKG+692pMHI/4bkTSSUxtofwO8sbKJ7y3FvyrQgYYOoY/EuKX3oJmmpL285
5QW0rcPjVL+cCasgyfDh5yB6qE6hL8m1xy7/ufNFU2380H8HxX9nWvNEDHeJlc/+Kgd1hrPhM93o
IYujQhu9VPxwLVORE11w4dqKa+OJoK1hdhnKN+p2rdxyXh9l9KDbDJkbvSB+7PQl93EPz+zTXglf
Rodn7cCuIv9QwG4GESzW3YXL3WWzPK4uL43a+ivo/7VC7JiNIeisNxIpnDlPlCVzhJJcZYfxoTBr
UeAOwL3aYjJrvInzvOQoM4gNRE+e7hDcUosQ58xefiM8SsfXi2hiLZfWgUpot/YpmEE48uzaMggM
OoOJRK69isEwIFIvUyZCRwi0akPBH0tm3bLH75MzPw6U10gHj66k1j1on0FbFHnDsO7tLslL87cW
VLPLMz7QqDG3v+En5QHgnTU8XW0ZJ52WYFJKIEzh1WS/7RLTUEpQCgtN98ftTDULaQq8tx5w0440
qOTmNz9aJU98xvZHOkPx8zXJpp3rYDGLkbgaDYjzSGmgo+UitfP5PTcvSyyFcETcCCPcf356eL3J
v2WvP7bB3i0I61XC148BrhyCzc0Cyb14s00STniif3/Y48YSWgbcLFNy1BBgt89ZZh264pCjB7Q0
z1PXQoxLDfgdSRiJHVEEeW7laslLc6AGsbwhJwUekViDWtTscKidhEVOQBq1Oj9vh68hTe6WVEw0
Tl98v5oJsG0tIgfOICuxntL1nI+yJatW3YXdtloGdz9Vw7Gig3S4g/TOBIek2/4TF41p+QCowjWw
eY5f3PcYKUr5HtzWmoQ2F+qFRZtapn09RiFeDpFebhChCJvgHqL2vl6ASXOEL3jCwMCG8+3MStkV
rM751CLFwXief7desSPFdFiZ2rHTBywbbaIMeBd9Giry54XZ+AwY4Pxq7/QXQyagoghsQLPjX8nk
woL7/2qFpzXRSt7ekVzpfLgBk3eqiE/1vaTXqRXXPsuSRAEhX7XUuN/Ax6vEOi6fsE7l/mhP1JkQ
hrwXgLm/eOygGhjIWNOqZNdOvbU+NHK7GdbSSjYvlKB7ENV9mnpt2fUISC2pMmNL58IsHCjD1aGZ
mxslBTFfgtZNh68qJwlDs5/uhFdwX+YRhCxzSW5EY5q36EeUjyAR+m6BCaxDaSJggjeHwN7ICnpC
8dGNa4Ot8DYkXD1UVpcegYWZzMw4lGfCt52acGEJDu3iYd7UkwJjotf3UrZjYkWTV2CiZquBKWC6
2Z3Mx8soKkniC5owopPn7uoy4sZNruo3k0NQTgAaKt+bYiaL5F4puTFa9p/i8PfzFyido2vx/alT
Gm0ltY32Sx9JeoP49d4MQ4BRvpv59rpc7/lK5e5tUH8VNL3b3mZezvQIQA5uujwTeZUlB8fNi2p4
qOEJZTcSJQNDyVb6RFPPQkYzYhxMARMghhp91o4jegtzVrJPUHD4vKJaZTpyFZvEa8GajOSmuWU6
okE9TWpGb1GHYgAQqelqJuywBXlem4yGJQagn1gcypZZSqJUt7QEu79P1j+lbaof+6Gc5W8Q/fwY
xX265OMvx5O+ioMqTfehQfOiV1uoxjRPJnfZtHfSRrhD7+gE5JijVTD2lQLUHw9Fb9pk48bJq88P
BWKs7pr458NXH5utwfZsXDPQ2shL6pUyWlGopeLhQqKLjKIrRIWX2G3A0xvDi16Qk3Ki3V3bVb92
hFe5kFr9ld6NSXdhYsa8+OPa6+QIMXWkuWUDhqm+wNFoWW45hdbyHvp/43gbsx7l3fKSQy9Wmv0B
iSzdi9IT3cZB58Sp73WWzuE1DaHxXjT1h47RfxdLar+8+U1sgxx5Zug4puiGCF0DnatAWx51MFPp
SB6WjrsGTnqrf2qPeqOwLzfGDXn39hZQUTvFIPJCsO4rfiyR/0r+Bu9bRCWQwjFL6lZ8CZViH6c5
L8L83UONPk4AjvK6pGxY3EZ7BoWaIjy5tOQZmGD3nZkBQF1q5dqFS+vk7/EJdbd/oXNRWpz+iycK
DLefE1vD/aMczHfH3Byr94jBih0ZiBaimX1EgiLZR0dcZLah7J+FsEsvHTwxRIH0vk1ZP6OL2H6L
fs4tx7P09irDD9WZcS+7CoRFzFbC26vvnHAmgv+BzUp0cN5IhGqYdIRvRxRkJVlj0dqMXN887wUd
WydMqZSLR+sX+BwWikH1YdL/6ZsKzLey5UHEZXinq9tBgWkh0fvckB+7XZtXhGHKXq3F9vntJdDH
txyHdiWkPW74uW8xEOEQy0OMrWhSiZerQ6nbNBfMit6ZOBX7aex7664UpOaVxFtH0lg0xruMLTEK
bKiqhfMnjp09Ub+OkZWuUjjnbEjrahzcvNPe1NvgWJkW2DQavg3TT6Jj5p9W5bKq7H99lNrfGSoq
WgOZjc54Ce9X5aQrW+nawulQvOsIqiZg0wrEmMB0bXuDYVKCXzPXeyV89F8sPCv0K3dLw/GJ5nmK
7f27Ny5p54Li7OqJZQgY4l4nABI0+vNenTpSgtrEifaDViranOKlQjCI8k4UEg7C08nYxLd1xhLX
7LS1vpsLpTq/ZCX1QWawb0utWFB4S0eZy8WzjXZrpbQACsMoNE6vj5eV1EQjeRxIb37dcnjdHp70
pWqERnREW1/O8ifMmIB9pEMuolzsw+CnffgXFEnmEueAMo9cU8iUXK9BNMAMySn8Xt7NxkF/GBPu
ynuIXEfAQPLSzcsNL9Jodb/w3GgUatSbZqx+3DbPIg8MrT72vTfpAeGZVksjSM241Iu8t5rQQMUj
elScUkjn829luSh7UjftPjWLuNNzMg6hhRPOtSV/sfHlskGQtB6etXRzHQ9D5cReSDJgghFD2+GZ
leEkpbyt+co/MIVGI2P2tNfxp3AxnEt/izOOlJ4syYnfzxuG1rOdcRbOSr4QMWHsqSgfLXdUh3ky
tKG5alR/TQ5xxfm1zpNyZcqVp6H4QqkuQ5vQ3iQ9ATvOPFSyMl2kXL5j27O0thy02WJL3Ky4vHou
wvVH00zDs70+01xQgiNjihZICF0bS70rqSXVgV2ZL9PgP6bCdZm/vXUVWgtFkbebhL8UaH9qCuoi
B6Y3fHU7HggH7QpiyXg86Y8OlHx1uBwRjTpeSiO7+u50ZHEtDd0dbK9JiaJKMAFwfeOTOvqnuniw
uYP7KCHao0IDiyaddNTbxwZM90QErZ3wY7VCAv8CJKDKWWVixtNoFeKWqOpZwQZHJdMpvNTyGusP
e8xK/Pt4rV1ioHLIvymB8JAT1H4AfydRk0/3z1cQBod/1OZTi4MJMgggvG4fGFlSWXoWOU9rzmVU
MOSWru3Qa5k5qjcS03TKx4sfX26Bo2TcKCV9ayXaHtOsBj6M2Qfe06Vf3Qzd5qXO5oKeG86y55Oc
p4fk1VvpyOmFUzqyU3Q7sZZ09PYk35pKEPRvFegquNV5PzpGQNsd+I8+pooNM/RDwZyzx9IS/3N0
iAkh5HaGEL2qk05vMBYRW/D0U70wnIcXEZKiJXZpKRwJjI9Nkn8Je4NLkD6v5YYAdba6TieUo6dk
ojmt1U4/EjgQP8wW9Itbeq01JTEe1aGkfIzPhWWz1dr2LRZbnmjbv7fVk6kpkGU0EVsFjMraruh4
hOsd5wuw8lNj2CNdqSGp0p9BF3JD9fImCvN9jHP8dhWhEb9gZ3B7aiO4GGqELLbTc03kqAk/O0a7
FVCX8js8kLFLwsTSrAu6Y952d0Dgfl3JB8CnT9gg+JvBtE2krTG2iiQa6oLvPqhnFlKyrY73SMkZ
mhRe895uwZs/IiTq9b2lEoIhNnHwuhm6Q4o24v0OosEWGuXFBjWUTMT8JDXM+o29iMpd0KzLnIBX
DFr9opB/NOOssbz0TMMXTm2xpnrEzFviNqznbshrPrdRS3NJ651DfQRqs6T6ObSS5fwagcVPiYZT
rsDETHSswDvxXDq/J/5v2ex+B5/0QRTXw/Spo28YS+Xbu3VKmQEZfjyVXhu2Sr1H5U0drinGfLl/
lr/XyEQJHug5v+oTBoDuuZzcf37kU06XptUD/s6m1nn54mKui7AStkfXHEVF5vOr7XH2YOj1Zxwy
RKkMlC0XgwZRExnPYeusjznZM/Qtwb6raEddPay+XjJkR70WFT1pER+hdSDm5QkCyvJ045wecNMl
Gfsz4h5qcN4C5rONl9fLj9ntCIuGJgZq6ua8PSXcOTJpzl1SHZncCuHsAoN77nz3d6cweelIDOiL
krgw6xOZBPegzufG1Box49McUKB8WK9YDxDjzRsomcyMVMV1hyBlePPECKLB7wk3MHyJlJt4tVRY
MXh2u2NqrTGwaafnHLx29K39EsFHbV6VCoaDkKx14nsu4y74Nt2j1zKIA4vWpvqg+k1Q5boGmSce
95wZQtzHVU6RFb1AkcaCZ0H4m+vQXX7Fh7CafPgaNFHGPOx5LphVINKJTewdGBGhSFvRF9BoyKod
yXZX/ETlzOVMo4nh7qlylBNDi5T3iIFG2CwvynBat6am6Y4CsI9mXYN3AUY+grtb/MS0UAt9Chdf
yf/Rut8ukXFTKIJ/LQ1OP2oj7rjIziUE3qlkuaWpPSLpXh2mcmEv9jffizH3AtwLwvoVaAdHTEUi
naQWmJO9tlwoV0KbtBXGcHQAkdOw7aIMRmAZgzsRrmDFr2H31AlAYdTxKyXmQ/3dc5On9oszoQGM
VfKzQZjX3btVrT3eIqCPW9srrEUjh6y0Nsf7U4VmhHcgm3wAxhvSVplLT05H6/7TIhciulVqhIfH
gR6DzJaAtXwYH6Om8gk8uhKb1wrhiO0scucnl62OV+nR11z8KzFc9T9vo/O6/Zke6ci5D2ank35i
abqQ9hhXb6FL5gE4knN0HK1pY56hYp8xHBK/I/XC85l/lsOV0qVzi/R8qkO/NeSbSNoHWaPQakF6
rx9OwCyv4QVSexjuX52DA48d6fH+Ko5+k7G+GXcTpVjodFTAY2VYzRGbZDWxs00HHV7rg8DIobhX
PFTeeNGziPt2LxBO2rpKRvz3Zfj6HtgPsLEWIBnlVBZh2CIHPrMHudjvD8Fl/g2EdhIk3W3WI4bu
m23ejbdLeFXfJ3a+vgYNe6PASQjL8H7bt1g0fLyhU6zwYjc4IjOtneO+/BEKnZvghFv0JNd07lj+
dhpGL2KyYSNLCzrN1RKIrygg4+3WTYeS7T5qZM3G48F8uI2/3v7GwtlNTLvJE4IYO7gZVeW3bP4h
4Np6X51OdbV09lRIMIyqHMfGethRrXud/LSOEv8p9mA4tVwomlmVLSDj224C4YkpN+R37+BriLCG
fUtIExw3Lb5WNjLqkpOcQalBxngZyYFI5n1MqrH9llyfAjKhdviQ+JfkxURBCr1dKVd0BVTlF98c
/sV6X5ZunO/U3p2DB0N9oEsaZewWA0HjrzzEc6/YCGNmT3lfVQFeGGs9SemPhudR4hQHm8k2ZpaO
R71Orqozun0exxmGbQO2NhFd5EUGjR9LMXP2a29M1/rUQZ/TOc9s9buKzb3CVpttYNMBgkf45Noi
C+2EE748jlmWfvXQCu3fr1rBxN4tVJCl0/SkPFLnJngaC602tkPUpAaYw9vP88/gD5mE8+5YjXtf
opcBKIKYVgMMhQRipguIh5pczeP4Jx9iGRWfdXb6ObEBc2dRmMSPnCVkjo+4ssGylxMp0uFnYfF9
70iaXJQlDaAYgp4TpKdJiZ78Pe6ymyV0lbhgu9xLmbIIYU8+lmfVX5h2d+CgPh6LdNq3DwaaKaj2
RTZXknjIR0CpNRIndpzrrh6PwFUsvrvpzNwKIkOqQHBxrfHn/Jhfunxp5kyA3SSypRPYdJAacQQ1
LIVFAwuv170VsYJehMMhMlqrCwwbPUTP+cK5dEcvJKYuBkk9I9ZKlCc7SWEaJRxjpH2qmDjW8cLd
M61rh2QdAA/l/vPfUHi5x5WirPYlKa5ExLl9OtF7i3VaCeFybmTHkKugYUUYadAzS4f6Sk31enc9
I7OgvOVc28BJQx6TFrx5hhscTVBZ1mkVkkPYGONHNYk606YHVg1FVPcJTVqn87JdEmtvc6YVs9lg
RUX6bG0U4c5Q6NE6VFVEsJuMcEElgYb6oyJN+my3H7qSdLxgPnofQzfYXmG+Nm7TGv462xAFrMcB
VHr/Rt449RRYLdZ92gKXikWA/rZQsU55gX2HMZ0N7Pl/DPQwfQPqyPE02Ac8SALC0U3xU2vKzpNW
LP1eX9NlGTpGT/4etBKXlefAGXwQqMnx04DJxLdTE6TJiDVMEdkzL0ZG2rAewSWzoda9g2zfXIwt
v6Kq3VWxcfjdoZePjqO7ssDhtuUYfkcpEqdrAlz8Y7rkCxOxV23DhTjseMZhOvaWuc99u5mfYH9G
jDtQ+7DzyjuOl2DMKZr85PS5gArrpRy1Q8STDyZUzK6LBDTrQEyOIWEYn50+TsDTP9hJ4ywxIj4T
uvIwcpmid5VdL8iYmi3ZTkXZe2MGViyFZk/3JSV9+X0pq7OiXxbcYBTBOWh8R3WH6/HMbTSGeuqh
F74AQsIp2TqReQLBeTOXHIr0HK6jFJFqZ9wRTOcUpWb0/K4RIHk6afQpzmRJ5JNWHUrYO9Xwk0Ih
7AFC8tlF7GmpUsLl2GseRTvPCa6NyYBUjNWl3SHCsZJD3cWT2hS4cIlqyf9X6s1iLPuHRK/5mVhU
lpgOB5iTPVMGn+yj8wUB8nWmZsK0a3tp9sGGP22ihX2Uy2Ifx/1jgLMXwvuJSZa9iBSqE8n+Da29
6BzuQL0qTCxg9AigIh9ctFFK30aTqNeucXJKHPhoaEe2Aqda33ywKAQ8Ty2gGdwf15F0+GAM4szW
ve4pbTd+XXvCpvHOlt++GPhbZz+qllPZmgsGspyFVlx2kx8M4+5qiYFuJuoZJnLFXqzTwvUAepDF
+YMKoUWx+Wf1d71Smll4nyW0VldgZ71wuVKwkmD/L6iUhafMvvyFTTnD+7jPtZ0L+We5PoPmnK23
iGIsobXIppiEUep0WOJchYXP+wgvag+tPWIFmAOU039/mvRRlsMC4NDaLnBOso3ydr4/6JHWErOW
IEpNxhHDpv4OdkfRboNUtjZjHVRnEuldatDcJxcets++AEZVqhzInHtZtrfJimJ/7FbaHROHcTs5
66PBOJaheNiKrhBPYo1LelT3rQ/ShuA5zCKW5E96caKIHo8iJGbjuBDn3u48Lu8sHblteTn71dSh
oje9tx6WPdvOffGS5Kuv+aj7uCDeRGm0gY6EQE+NJ2rksj+jKsY9gW9RgbhaYUrlqjb1BmMUd8m+
R8iq53dv/XPKl7gv6LRKcYCNbUHxHcygUTGroUpGMwGTclEgxy5nfDspuDqh5t6CNnoTIMya2wtO
KI+M8jP/Dqn+8gaqktOHYzvaWYkJKX2HgNBMseHoZy+Fb4iuZlLCD3obgCdRVHmLvskTn+crMVVb
Y2ZQpCKa++IdfoM16wEdIp/xkzD4PEAOoQ31Xf9JFEDvonFSbHz+8NV3jB35/57bhQxUdi6FpEK6
rQiDRtpuSd9jP+oVzO5MIHt5lLFAqRQlLBCsZmQ2EwwFDsK5/DKGgWryMamDHIa5dQS/fZWRD+/2
m9k0Gp1K36s+8Q9uXDTqOG0l91F254PllrnQCWkMzDUIO9jGeLnh/qhSGIKxqAcpCLdWZrYqNlFj
fHGFXQ/fURXNV2BjePHpKU3++lo8IFdMMdOoEM7dktkMW+TTvZLc1M4RjQ9Sp+Y3GDDE4BgguWEj
EX+3r8AHw7nN0nenRei3GJij2ECz9PuroV1Fzzva7ySvh59uK6p7SpPh0zd2zoKCRxS6vRo+TzkJ
rdJdICHOr1uzf9H5r/9Dh5IrrGfoFoqdYDFInOLOViL87s/qHtSyUM837IV/9Z6WaWu5MOvbPPEC
2aJltR9GZa5XyZ5UShqpgWDwxuKrGaTSVwvyT9tv/FOJ7nXiOYWD+0Y7jpCJbYQNWAKtY0I0fDjD
Vdhhk1lE/45AC9GvCxHpPum6Ui7qshZXI4Na5GJqtODjQguCTlM8F2JK25Wxy7klYQYKBGx33wlE
wXEE/t0bUyr1JC+YVDAl/AqSTSCU76QiATmr1Z9P5b26Ua+7X2FlHASew8fgrL2ot2SwGu1Ckiso
+93JBAuvqPDOR5QL/oqsZ5bVC+Krxqw39ny60wA2l2wwds/SWNunIy2gbEhhy+eAyZgJfmE7xwym
5xzLIEZ9WcelUFMxXJbHfjzteshIOeKH0KGL9pmT8q2Vol2bHBZZfExdovxMZO7oXDHkixV75IIv
6z3vnRwWhOnOt2okoYuM0grRGO30dL5V2P2IrWsUpxGMZcbUN0QFMCBAzFijX1N1xHh+Ev5NqDZr
I3iH9fp6lha6csiDfrINPo8I94BXsWG1a14FdFk5RCBoP3hDZDujkijGoXeOSVGxW6SMusObwF4V
IbVarNQzrltUK/ugCB4O63rUlpoZnaWyVDElF8wShgg7exlkMILla8SxSIykhM+9fjb9glR07Xgp
jaCeYuM0nOoT+lzIivxqP3AIUJgtkXjsjeFOJoAmK6VMOoM5fwZQUb4IPbFL63UsgrldMt9FrDa3
/s3JkFqNUu/cw2K32bJElXtVL2I1nAcZTdTB9K//eGnF+Mjr+Hpb+wOR/1zmOfVmR2zqWrJguQop
chv/TJUB0W/5/t49rhByMjmieuNzxBrNOcrg+QbqIVzf+xHDC3nQUkKMycniLxxC35IAN314W3K4
NoFtSrCT37NyBKj0/BItfKR0Td5rwtyWWr9j1atn9hZByfPPj/XJ3p+8LPhG4Ezvcs4f9XriJj5L
O6zFjcIzkzYay4yNDiz/0Z861QkHCZHg0S2nSaURN2wbcMQSmLDzY7qJyc8WN2G7NNHWVtu3tEUO
lN6uY/w++HfdGTqeJq1P55P0VqUep4HReq6z6u9as3F84f4tVKO2TVIHeaofzY2DlH2sXZH8Uzqs
J+/C7bWijcvRUuPpaGTRil57OsOGhEbfqY5CkHiJ6DDMu3ZGdshJly7ZFMm9vcKWatdz8fUitSlR
h2naEgXd8mnfcXfviGwQThYl7O9FZWW0OxMoGhzOrv1kYRmi6zdqawzYclLbRdsTe5C9ldiHknDk
PwJZSEPnmMvgemAy8vsoGmX1oH0Tz6q+6AFYZgSWNCqyFNUi49WRFBjBKOwzgdpAAwPkTnpAZdt1
zuyqEny+VJgYp5CkPrBkvzD3FIAvn44GgqlCDLFCrz5LNvdSdFA2MDygJFqHSUXG6o/5BHt+5MBj
UAfxMAzhaB1lz+voUsSZwgkU3u7NEO6LL+2wfnj6UUhJxckvjIJQPq/ebbkD2clfvVkcb9gbWbIM
FbsGYrdMPPXxdbb1m1c8PAKv9t8kFMNyP/YXaF6pektmtkmDdZDmDOyr8t2rxNWqoBbolylHEHfN
mJxJ+LTWAltFfJsaZOIxKUlK0ZVIbxVdGdNQEs7YtbetnU9bRn/fbqj92FunIT3mGyhyfGZ6J5Gz
25xTI8/h1lYBqihzYTsZpkz9qm8+fm7/O6rQh32HA18RHJ2L8rhmhdjOGp4EOQ+/qRDb9tNTAi7t
T9Zn3y82MsNuLjSI+u6FRp6fokT3Kp9Tv1oEV4sk89lEMexPnl1xyA/atzp0jbK6TpczIhKZ3EVp
fsV/EHWsEI6YrjCNm4ytbzRZZzYk499mqxM9d10dOuC3eQFZ3+GCsVsKx/tAk5ztbRSZqYlUuhR0
WzWRV68DxTPceN9SjjstAnlswpUoDHq1+BZcl0Dh/NVYsyNNmX6JhK4Mn66gZdOh+ANDLA7ZZc27
qspuIVSmgZiC0z4ar6vOFwZ9Lps3T65GHlEMPKn9xe50alO8HvPgmkfvxH4aRkwyCgecljZNG6RY
l0hFV1yDrwYyEQZFaPV8IRuy5sM37gfjaryTeS2R0j1HxinH0BcVY3ghrfx71762Z0bwsVz9Jlwo
f0X8OeFIzUlrx2f9x45Z8yHM0YOeUleSuAx1fxpaOM9my4qYEm+pkqOB3MhQusZZmhV9AbdFIbc3
mkkhlck1UjqJRj1ivzd9rOmAegSySYS21/TYxXejtTERUlY4lix11BCgUVT1TIUdMD8srdamZJna
8v4hs3UfOJOX9vto1uXnVyNtJ990K80TFjVEdmdu/NMS2mZvjZX8ILFQW6akEcVc57LESbyUmJP2
vwF9dWa0Tjo10X06I1L61DaVzpGCRlPR9m8JicBrr5Wx8Xj9DrBLi8pNsrT+CWOIIufdn+x4VZcT
e0lEeuMaYcZYj2QdrWs4wxWTLr6mQDA4Nb9kqj1YroOvnzkqzN3G+xBjRANao37oXGFFHrLcCclQ
uvCCPaHFAGGUUhZmPjZsQbpbLSuXNOhaMiG+jr6X85M5WIDXdX62UjTrBRPwIgP6mGO3Di+JFJZ8
y5e9BsJQIEmQYaHJx/VqpJqP39lOX9Yy0LqMUPDNX5Ji4WG1QCpL0v5QqCFb2bVt+3Z8D0lzWuyp
exTCjaMWQSsJDtT//8Iy8Z2GchwZJgZ54hRJG2AQXOpSouDq3OkgV2N9kKl/7596cuzjXNBlWNmL
BxXUli+ZsC0TmnsdAnbbTjdoHxJ7c4WUwaxySZl1ZSbhhAc2l5E42PlGwU4R/Yfl1VPHVUBIZevW
CBJyQCYb4LVAl0K3KtOG/bKeziEr553Ak0Ap0M+fp7Dm7+SpzfmU6WC+ppFT0C5ZIbqDtPgkTHTg
D3gNABjbS3VMJTdlHrpoEFsywaE2mstxF34L1S7ouIi6jcSksL49flDQTscbZXfX61vkHnnN2ngQ
R8fNxrbU9A608znJOKEOOsQuOKuiqX7/O7XvjPjJkaplvz1Mr5pXeGlnbI/9Tib7d0BQfo8l3cwz
IhS0uGYJvjdWBca6hrx7CtA3FBTDKhosuwhnsLP8WKXifGH2sNxNRXARoiEqEcZqv00XDjhIGwZY
0lTkXsRIb7qF9I1TE9KCqDjnQcr143KIJCiw6irajhlR1DIbI5bFg2RfIXiI7hwstsGs/8O78VQO
N8zYeK7028gUPlaOSurnYmw2SMSP/0L5Pl37v+0SWGxrUDXm4cohaX9oZJkznsu1eYk+X5RaHgys
uNZ3bQUMgwzeu8ihLmdoIQ9D+Q2vx47NdbSp/X1bLu7rX8ZCSKYpOi7TI4g/ZXKYVL0n0uNMHrrq
q5SFl/eRDFrmvSXU7fJRbd6hX8C3ivrNSqsjfbbwqk6pjmkdUvumYyJVwP9DHPZosnifLbeOBnKZ
gHJurJusLLctnFx665lDw8IQv+c3BdMaZhH7bez1W8l1uHFL0nOuQjZHcXEKrAHU17TFtPKJJ+hA
DifBHCALqRASOrVnlXip+eI2GFuQOzC1laDSxoD0KM2tV19joJlbSX1Xrwkx6Gmu3bjMdNHJzW4u
g1FFTf6WegrxQ6GiCd6Xbw49mKFQJQ7/2DLp5G9OjkmAkpsNS4QPp+a5O0JRpME54EqJttHxdna2
NW3zHFIppCX6Qq5SEp5ebw6ihOJjMcYHZw4pNL7vgp2cwdZSgQTBT3wCg4QN8ozxmEQLV/BHyeAR
ok6Lz0kNQ2vcXHcbJMjACeYsVopdmrbwUzX1ZbAlpa53uh0L/O6krQJEbfKkYwNDVhcyrwkzAxAF
N6MD212SIMsqPcreysk9U3Se2QEJ9B2EXGbH8NV2EXIIGVgDDmk4uUYZeQHDEOeLqVZvb5w6XXZ/
FNoPunIHm2pi79z+YdWWuVMzplLlglxLZMg8btrMhyHdZsihA51Agil7fc6aqfNJ3YDtMXYAHyIp
d8FnApBMedJwNcd+NdLPHIoVBAHEc7mOKsk+3ZhYgBbFDZA4F3tX52UIaDOFrp94fzxrQoQvGLGD
au9EgwAQ2LKe7aIOksrJYzEf8/5nRnsq3OBSHsY0y+hpUFEH4+1eoKkTL1GDbmxGILdE72c1Gdpg
MpJs2h2ZOYhvBkbE+Mb+HQ+i7OZTVTiu1OE1is8bICdfbC3K+U9F/8TERetg6leyHo3elF+aAQNn
OPdeYd0aqr2E05FLKK2jvywVjqFm4Uhm4/Ed1chCycAY4sS+iCvgf2H6D3+n0ydOZ6UDm9gFUQ1k
o9oAvf4vPE78x1AXGm5QAoQjZF5TLdXzXI3bca8FoMk1dpeX4IOwG4dprbsOzr1felRV1J72YV0y
lqbK8ytkFWJAlumC4In5Pxbfhu3ILis8tqxGEVy/jMCglX1AlLbRtH/W6XCpZbKLUiYFwDeXRHGf
m1nG6x1aL7b6Hy5bV7stT0ByhISDIQ5y35sThJHyIXZ6tk+V0mIRlQc3bvO+aNC9LhpXFn2l57wQ
uEfbbMAhBKnQ58cKliS1LWYP22NK5t2gu2zn8CWMoBwowYsErH7u6LkQ7GRNHHJ686jcYFAaFxfh
BaQ/HyKvYff2Y6vzeKvfw0TmUYQ6yL3wqOGGddHMyDN646/f56iXx75Sm1xxMRdgEXj9aaBPRnTS
iIWCIsooIM1v2ysvetLTk0fc+VrpViO8GvbTXBGvqGUFK2GASg5YhWQiqLXHAMqEpsaqI/sGv+KR
hC3jv7/KzGggV+OuJD9ofMMUUxAUxG1E32qbRhXd6nMZyAKfKm0avNEGXNSqmEivzr9wUZCi1ZFx
YO4zqTIQfl4wAnAq3LwRhmdK9j/vduEc4YGj8U+zY8r4lXSYlXuvmX/7szUfA3BvZwcqN7lPP/zm
YEPgvLfo0N05dUVRRKigEVoUEydZnbijuIfHNLoptBN0gDo8921DZ6H3D3bDL+r57/Wr8lCLerKl
3QdmfJGkvDQNMXy78PLB/wkGy7Y4zLzbehuV29Ss+5+z/0PoPzvY6J7Z62DcMaoxJV1r09D7mE8G
bRAzcnmLvEf9Ign2MsuZVPVmhwD89ztBsC6Qt3mESrkDnI+4y6z8d1jwC+vZlogGaPdAfqj1vNOQ
017NT/ek7Wa7C9C1JLYWz+bnN3Flpat8JSJGiQsmWnvGnHPj5j4tjGy3qN5XWS0PCVMbqgx++IST
DrftIdsCGiS4pT2QILrxpkMFaSBV3sJtN3QWUIyC6GhaMqLoBt/z3CNZYt/RqZvQqFe/z34CWR1r
4gLmGY/qtHuwB7/CEJS9gnRY32YC/Qm4UcnEa303p8INlrlRI8uY2BT3ke6x0c0uN0XD1A1OA6Hw
v3SYMjTy5kKnfR/THT0PMPuSr/l8XwJ8v4h/8c/VCFQfZ6D/kTn3qF1IM4168vOHPezp3zUAUfMa
p6J25BryNr0DvtGNpiGkzoXA9zkY4r+l0rCQgNIy1mpzQJsgW/LlPTv8REFYzruzoAkzKu+rsDw1
l9jFT/v77wkdZcsEHBZdDy4jw87iXxldExchuZbA/NJFBANs8Loi+m8AoJMX3n/kk5Y8dp1lm3ru
i05fVpScMKFn2eM+dZrORCLs8wSRAqArQunpEi2MPA4d5eAtKIkW37EPFB9hfIMiqiWcR8izY+w+
HN35exnr1gxAd6rHdzwt1eujVeY8WuRSuWEMaXiYUIDX5qa0enZFh/ML3lnQHG9BrPlGAPX1QWz5
kYSSbvpWjKdy2HQ506cowS0mRmlcJ4Rv/1/arz8H28sBCVssX+6j+uu61nxzjUwZDc95kvhhXbaE
s13dU60P2Xcd1/7Ol0U/pIHKXZzR8NytSOPmi+YeKdNJBTZb1n7sjaayBoZmTBOfpISvWoiBOC5f
DO77z8d6av2qYUu6QfLE84cqnxOlhXkGnQbM5BzN05BTF58fm4Nv9p+nJZVH6VFuSFXpTcbUg+Yn
5OBvISoMFGjdm+CpdUnwtb3L/FD9Exbb/qQBpllNRZcrZ+2zGuWLVGONcL7UkQVmacRi0SuB13jr
IqE/NsPyDoDyb6El/tWCO8xHgHPK158M1wPaAlYeck9jyIXcuqmFL9J0kAw8k0LLsspkGQVA/kmG
WuzVCYtsCFVCd+FHsMX8lViZErZWpDKogWfvHcFjdQO/3BIHC8DTbA2utN4OaEShGUl9pgv9njsQ
cmNWbNYrB3NwVN2Wc34ptAXCEgRGGp2IEhCZ8QHhZc3vKytKSsgQfbclMogdMZboeZFziiu/3H95
Mr9KAkKJFmU81UhVWBb0svQwVLMNsDAhFs6I4Sno61m/Xw6YSfckj3SPguYGUdpk7Zm4pBF5Y4Ql
+DOQmthyDurVp56w6A52A+HB2iZ0T2dzTPflGWMlp9/bxioC3+GWspyqyUB00l4fTX8WPITtQnd6
2LUu3sL6kdsGE5yfLkth5prtT3KsY+7gM2QNKTvFVWxQbP4WwZq9y7FhDUW4qaja0irKMdBwS7FB
XaJKhEKXxy9uSNBLS5UoDMghbROt4NIIQ/iN9yJkTy3ChYxiUgziJYH1Rakj6nB4QnMS22YqCPGD
AmP01lmpvAqiApRAvUcU4Hs3S0cueJCZp74vqv1ziPzZfQfw0Gu32+K7mdP2y50Ct1+vMUCfOaK8
2dUUurRpIbZ8C+wy+yqPp9rEshsX9KuQPGwGKTFSmoNl/5jmbCIY5e/EXS2Iq8mfDjv/+1Lmid7V
Hld9u8W2zwjU1RHwVO8mYIwQuFn7cOW9swmPToLBy1fYhSOPh4+MZd9MI7OjhVQ6mx4HZIsUGQTn
qrr1urUbmljPQo1i5kR57iry/4gjGxTQSZl/H7q63BxLJZpbYCH/7tcz8Ow+dgXxjh/SLiw4L3Lc
nkSJulwRNYoPvX00E32llZLvAMxzhvIE5N77oeNN4av/bQa6OeN5iwOrbAJqvYe/zElhtMypEkv+
k/Giz0ceKDUQty/ddIBtXYChnP0qQnb3jIf7EP89H9YwcsAYrZmeAqXFkMNQa/KGMI0TtbKBVfak
6wFZiM6niYr5YclmV1yWqye5PNWhNnre6X6Bar9ML7JJPNHyeMTqceQMKx50upyC4rfJwWmrDmDm
JJGBe1P4TtSN/tq7wlD7W3uuExcSGgHLe3kBKnnBurvNyEAFMVWiRSSOuKifb26k8nmQ4VxxDdw6
LItnNtpa5q4bDN4gH9Z51bgyz/8ToxlUlCB/IJtgoxb6q2FQ4qsDF0C+/GFYP02I+FrOVFrotpKW
Us/GTiL6N+oxT4WhymLMgTzne6QfuerzboIDYHbJ0F/kFyQ4SNYQSHJ5lUkk+Jb/ySpSaWAPBLQ2
s/0icCqboEoOfVR1srRtmC4c+X9uZkTPvXgEfQgHnLgr2/Kb6Pxs1lC1QxxoAPQdEgkhIABrJ6f3
C3T7H/rOAVG9EMlID6MLr3+tPw2HPgFIkpaGhjVbjT0f1EZ+41JEtxgwA0MDcg+HtYdczLe0g13I
VVhFoI0B2JK3U/HMZXGFBvSBwCvzeKnOZ783XDQWcwSdKgs41+dspDEZmFKgntV8iq6fxsFv9/eR
BuH3LA0RsLBDoKmfY7SYXGpVMFZ2BUuFE0WqqMrCqUXZHVPk2pKL17GOl9fp+8s0oLNiM3lUF2W/
gQ70r6ntEn3uQ8ebryHILpoj6S2wVtj1yteIvKMDK+5Y9OglOuBZvkg4E7H4FFhKnI9It+3/C2f3
ahMwlEuVoFCA3kLs1EbWAJ+09VyVOuUrdlN22zSUWS/m2vc+CtMzPAmqD6eSoCZonbHHZT/vyoRn
f773YQUmcHc+vYmS4FnRQ30IVD4rQW3j9MeOsq1KGYXjnc8IfAovaoBgP2GDihfokueFQPEhx5yn
Z/8c4v1vdr/FGAqWB8KwvfNrsDkYyjCR4sx5HXYzF76DFg/TMGPP/1BREOI+TSiiIau6Y3orcrUa
5vRxqCmQZIdcFVemz0RJIafGdaej81aWNI+s47HyQiSTKB3eW++9vVmzumAhWTNTZaMBQPoDKEhk
TwoJ2rZ3hXeYDkjAMUxsi+uaNkkpC5L6wO/tPRFH5JghQQBc5MhvqhfsN4RHxJRoWjJUlM7NDFZn
m/8rYzKzwaxqG8oyVxNxtLO+u6SeSJsXd6SMJPgl3s6kGpmcUOXKZ20673BA2XZPYTUAsgAkOlp5
ZjyOuVEl9v/L8slOf3FKqrhBYzIlq/KqnTUxbEu2X4o8U3W6y3JRfgOV9EnZ315ceFfeWuDKtsl7
ta62Vge2WDatNeVhNat9VSUKBHGdLibHS2BAjJEN1CPZgzcUIXSO848Z5HCyFoXfnfWZ7VNYE2ea
W3SvhyE3Oi0wQc+c71ntNi0gWCC+XguTbI0iwo2vDlW3vugH9PP6ZBhaB9LWn3ZyhwGQmiMYsHJm
DZ7qtDPKDStRLOx2CwFvvq6wSCnkzZSlv2NfMGqVC7CP0TIzU+KP27ml6vUh/tkbgBozLfRqxsQS
RtrpxDwx4wixQq6Pbnd5JZDgLM06IdxCPST2AP/HmsxFFqBW85b96pFSf012GZRfgZrCO/bYHXn+
I1vU4FgM+KC42nJ5akKfLPDnURbyL9cCghVmBtUlVAlE6DcYUwxDORMcuzksR2EhRsTTX1+Fp7Iw
UiAXphM/Mv68L07pXoe1fCSJaWpGgV+3pFQf9bDj9Snbj2l6fpNfKd5pEWn3ue9Dt8aNVrhIo5aN
6cvSHOTOR5gr5S5QG3VC5lPyCloSYzax/CzNHZ90TBgoHBHfpiqDCfnFm4/yVdC0RQsDmD4XqSae
ZM0L/gxUqzRLGz2ohaBsMkSfcOo3h9FtYTNWzOFf6RQo7nU4eHcOBPvFjdr6Yba5NHsSPc9zPjTN
FUmse20KAmGVFlxnkMRT4w2ZLrfyjLNNzq5kdrGUgkUjl7BlWhuYBsosdYWBXZ6lYr0hygDnlsgl
KRajY5ZfVACKajdXsJuqwrI+h3uTXFApkQM4hB/WFsYD3bFRn/GV3ZubVC03nn5JNYdWQnpsXpEa
dD8sThaauNnh6j7OqEWtQ8zUm4zfZU4pcwGgGbUUrh+siZhXe9qntIZsPChYDVcDbXaXkGy+QOdE
lrZjVJkJhZHMWfG2O3R29b3vLvSKi7pV+WRON5CliRIw0wzXJncB6dgbaO6YJGzxqrskM1Jn6kZa
OvlehtaocOj0o8nfhCYbRVOuDQF3qVaiVWSJmThiewM+j8ADq74b4wsNVPmBdsirsnFRsFWGL5ny
0B3eKYJ8Mz/ro41LKNmSxfi1w4FdmRyJ5WE0qNB735rw5UKXXfTUTJq4ci+se+DAO2oHU9KBxD2u
bbHQlwI6URGH5nVx/vWA6JlI0U67VZXEBOhN6RyEt3Fwfrx+frzVp5OuaxPzj2Hq6XIibLzSeP5c
Xuah0z3KUfWyY120l0fGtn43gV1/mYXnl+j5dogv3gsdrB/od/efWlPwcgm/m6HB3OVsWeX1B9b4
OgZCg7hGEerpfpfqTIVnC6xIeW1FG3ygJJZ+qvWZw95crx2307/5JT/pWw9Uwt52GPneMYTwp7cH
0sD2B6Push1DuHhe/cbM7C+HJLkmlSPo3JFYF8qIDuM0UvuQnK4D1WMhv9xCTt0nQw5RefuyLBaB
S1rXuBeXvNNvhACa53lyghds5ThestDA77WLsYvQWnh92yj9CNzgiLQW+xyI4h/5R+lPVs6qHMjf
Ae+mIv/IM+1qvoWTr/i0gkHnxDQ0fPs2sNT4cN/hs4M/zRTJeW39ri3/CVLtrbMeSbazwbRZKFpT
jVbusuuE6Bp+5o4JP0C9rlTUxxBEyD6zn48LMEjVQ19YZUwzh8rJR66j6fxMdaFniAghZSKG1709
f6HoWoKs3+JpqoKDl7m8cnJSzPJyE4HDggNmTBTyr6MEl8Lw2ln3bbTf/Cb9wZLCbh0AdtfYR0xG
O+/ZQpBRlPWdls1JC0PGablOKmvWyWW0oS3K+uxO83Arcg5X/rvDSCTCdyKLm4Dmvw0l1ajRLaw4
ZJHouGiwVC0epW6UlM6mZzSipieJ3KMXvenzjt15Az9e0PaeB3YDzhrfxGSGQgk+g/RMTojb6D00
coXF97+8njhLjwUjtyZftdB2bicPMBJAGwJhS/iNvkJaS2REnE7I+bNGGwgSVLDX/kGQ1hvxT6nd
G+iVazskm8oTewvXIuT5akCjO/wcYiaeusIUomf+oM3GDpG9bsgDHba1Uy7MvEytmm2oRioxAI1f
OSdVPpbbP7ASmUWkRAH4Yx+UFseSzHtF+yjBWmouAabQy0mPhylaWBNuMSFbCgH0jP0M7pJxnodG
RdMhHIrtCn5vSMWT7r+EqD7V5bYTomDFrZN6A31ZtE8lzhzy4W9JVpgq32gIFngJiA1WN+N0S9Eb
dbIkTm6iclYK/cu7TUyditgRDBsPyovuP+zEo0TAAAN1+pZDfE109/Ga3Ut6Q+mACWPnESen/N7l
apKvp7iw5zje+UEpmIS7BzCgALb+s3zmgAVnH3c+B1IwOcdd4Rh4A4dcUFQsSGAi1KLX1I58nlmB
pf1cOaszAj6JRkXIswXwfnDRU8dln3BVdfLgkol8hKDd7Q1dZS0tIY9NbBh4vvyd+cU6I3VAkj2+
IXSjlwW7MCIKUoa2ichqLj0M2DZqzVhUQgDpSzak9V9xkmYiCz1TM7VbY+cP4BDs85DRr4cNdbpI
shd5Rwzbj6BWr/V/E2TnAGV905Ms2LVMs72w97JGkm8hsWRnFawJHs7NobChAp5el8e5bRzEX5pb
+DEYXdPL6khI3j02dGmaY+3aDIpsGNoke2PjGNbDv7s0nWugtR5H7RN81GNPapnIeb6D4DQHdzD9
cPQYwgMU4T/5MKJqu9BH+LmiQr+WukYeUJgNKjn9vy5s7iZ/VCt5QGtCX6r2x95qswKrj77H9LLT
qUJ+pajAJxP32nyaoSJdWBsexSoX0e9bw4+oBAxJkPLGCGQiGrGMnmxW+VzJlMCyyHWOIPIVeAPA
vOrs75ZUh6CONp1//+8je0L/tM67PQNWds4aMMtOKjXYRvM3nLe66AICnYL0gnYoiqbjk8Luv5d/
IjMu7DLFeIOTnU9z2sazLWioeRhn3rOUs5aAt3N+0zosem7/HqYWKSQKz4SgO96WF0l6HbuIHVA5
Uvt+vCUDnDxVUiyfkSG6uVSpjLKecYFs5/0JB+j/bZeg4PjGEM0J/sTSQae6lV0Qk8izRfW/sUO9
Z1qo9HD8tFYitvM8vJOOcWyUeBfgXTsBNTFxb9mX8sXLMJtLJeqtZe/38i5GKnW/1MBvpV/qd2ZU
Xy6nPVUuX03OnE7reOw6XDb4pNtF4YKGnRevq7eKAnqz0RLjHe4xhTx1KUfc+yi8y5YescwQri/z
AfuhMAXzLH9uA4zDUWKgTVDTmVi2eRfsrZmrWY3FGBzgfRXIk83yPgX2EtLseqrRFz9T7omHYzYO
+N1X/aA7s6cBxqHeFNDXON33+av+UuyQ2znpip2N5M4O7+Rv53Ab9iykav5jM/sIjd8mB+pJ/1Ce
DdsbZH4JzSZCNEyp0VAZ0dlmnbgeH3Il22DLe/9o7OE46oUxJV1v2sWmYHC71cK/faYDGeP0JM0D
nljtONn4Pb9hpPPRUcjS8pk06utUw+ZVDUiORY/M5M4y581nTBkQqMenWWLiXV3LWohxL+itX8bg
6ZBglyZkoUyH+8BAKWz+KQgHez7kyKb2ytyjm9z14E9zucqTn1HoFJ3OLaajDvkjP2MUgX1PL4XA
rMR5gSO6j/6278yPoHngjhYvww97wLCtJ3A4k2f8CslQYpXH4yM3yBsSRqaG/08xC9EhsLvCFWl/
AAm0MjlZCDW9725IUveGKeIQU1xEwCPPzHQGivP4nWVlsRf47X7z63PIHayNskKaIJqH/MRZRFQ6
F2Qn87FO3AFfg0Rpmarh6lXQI6NC003FUUT7aBzwVT+WvmojLfidr6mEDxr+i6IKFwQ0JO1PJiYb
2Tw70Xlb7sJcaQB+HpXQ6I3hToTVmOwaqo77Ajwc2+4MTjWbj6lYyqxYwby+tj4ILcDbaHCl3J3y
jZ1WnrU6dysL0jSO1kxVOtVm03LSuY5KQYxnD3sMpfxPq84RyYiSQxKFF7jH06kSdk3q94YgJjA7
QSJfY0j3VlwghPGszlmLUz5spX6TsvSs6rllmvSHm76jkjBDK5DWIQw9KAANU4kfbAWCVkYMY1pL
pE+/TsDQs6qbMXTLqEgFuNqhrWCe9wXAA1gbpE0SoRhVZ1++UZGN4VTSJtB/Nw1KIfirVZJuflrC
1jeuLC9+/0iW3tRxCCD7W1DCkIFn88g74zltq/Za77XPY6A/WfJiSf3fc/+FaOCRi+4t4Oc4IV6D
qwT5lQ1FMOyOIym2RUGXvZ5ZzWnWuK3BQ/GOq5IxniqipNK5Sr4cFAfvEdAtqMrowgCui0jXZn6o
OUgqkzrekkeom1fzClvi+KUZLt2zE7unojtru5nMy9WnWQ4rx4CkFYBVvjNO8T5UlclkzHDZWNpb
zKdd4IQ32i2jgjBPH2nca/E9yOgzolnvHQVAgaH8R8KZOWlWq5dvYS465FiKZU5sLIU/B19DIPjC
/0u4vIqUenCg7iA1j+Wo+QTmagflHi75YXrXzusbh6A+5gwb/s47U9Bw4q9NmkNBQ10PNah+xgFm
WBDW4lf/oTcCzZgk8GVraf9xVi52mBlm8I1DAU76URrJFQjuTcBBlxnXkLWkrooCMewwnL7MQvX1
v00+ITSRi1j3ZyVdF0/CUxNyiCwTnpAzwHySL426leaLmMeZbhbMzvmWe+q3w6CHW/RxHSVa4uj6
XcKSXVmoM4binQkfrnVbxmAR53xZEnDYX/v29s8ucHX+aWfuAuL4cDn6W1Dw/hMiS4QNTRM3bL+q
AICGurscfGPLzOUTf4hnB3I8C/pYMAXVY29dfsM7blMNsoFzXh+MVenboLNIBHceGdpPJO292fk1
w9Oik+Qevz+OxJjNo3x9+TwQdf8jwCJokBZBj2RXxFrFKkv7bcxxZIoZdGtfRwKy70NOspRlor2L
Zo/S9hpiM9HpUB9A9kbPDtKwpVP41/FQUOGRTZxIvz8lYF7h4q4CcXesCFnI6hiACyIBhikA8xkI
a9hvhOxDDdpGv891zXPKR0LHAC+IDODL94VZ5ky0ykM5vnyhQvPXsJuxkl2q43qZ2e+WTZgFHlYY
eXVtsPMZM1dWKU4rF2lrKeH0+s8NJpxM/LCdxEVs08pSch8/qNNbN9m/fJEBSrSU0E+S+bG+K20h
ZHXbM3L98rT92nXyVbbzBQ8nVXUS/Y5Sq929gQW+NiEVIjURyr59c4GmQOkucLdyREdQqxQAySH/
CfPCREAlszs5nYoIM36gi54qldbp04mZ2lGwjGgiwoN67buFZn+JuDQJKUYNyTX6WhgDhY8W0WIi
mMXo4J1rzMsdJRWCsqZlFSOomglxpsAz8Zq6BVbAxYTn923Yu75006TBeY1EHaHeaFNWAzrvxE+A
6csSOvGcGoy1188aSAH0mFepmunlJwHUddAmNJlxmVf7QMC8FOnLEO4nSjTlnPJ2xQi03/KwnL07
H9hn9dN/msCibxfuiGxIzkXgv61N2IdNAYmM8G7Xl3N7dmHlAYAsv7qowJTQWIdKP1EPVeiszLXr
X11nKnj4YX8q8aNz3oGK5iF7LgRQOjA1dNJAaj7jI43usBn3WYVFAaTGofPf2yXD49FPGiLlpN9g
D0ojVm6FnguQXTkuD3gNn9tU4NgJfEuNQeKkBxrq8w5QwnNAuU86gohokdCeaBP+wTPgkETXhnuQ
3iVh9CKx+vKvqMVdR3OoRpiki1fOD0ll9lddpY6R56VMXcgvtV2fil5LI/fPaOjn5lPsI03o8kU6
V1Ra1IDeCamqpHD1cLiLwtDvdMShw4ag5lHemVu2N14dsFsLB4JADS/pKZYt2+JdSRA49liLSeQ9
HS+OhnFQOwAGW3uP4w03r9/CMHzTftWwiqaMSMsCKwe8BF4kgZN5B2nFho8KqCbuHLtH6RFN62S9
LPgqPTuCYKAgueob5A6pO8JU1KzQbun3Wvhc7lkQcr0/VvOxuQNypbJn+Rw7QU+iFKODsKXIZmDP
ypqi4YMQ4t5bNOU1pivAogeZocBzGUzXPVe9jnXvxEY9PEyPg3/eWAIyWd633dZI7+kHWNUkdetF
R7kYRy4WaqPz73SdppPqRqqa+KRP0sveqPs933Dm4oSp0KpdOQAmvSnsg403VEhrT9Kl/WanYO5F
lmQGUvrI68z2xtifKFC4QJevseVy90XOjV+h5b8m+7sElMqei8CPGddP4K05hz2LuLmCfaO0fljA
gMb5R5xdIdcBbd5WVeGbOK7/EjP3q+vqoCsq1zkr6puzrZYoqeIEZYf1V3qIHl+7L1VsMv91B3OF
JSD24TslB4mBLJe6JMgRQgW9o6HV2unAEeDCJwDZYjoCDD10QlgaGCarCCY6jPcxzF+oaClyJLhc
ny+ghMSebOYmAX4r0Huf/l7bdg1YtaUZlnGd2NreomLwX7fVyMXWUeWboPsAodGF71AroKxOUyEe
fVFQompzeDEIbF+3YUtgBH+qKCz/CQZrbTZbkpp3TAJjrVXC4EwoI9hB2DdRfREgWtMqDGpVaCRz
s9DNHG/mWxl2AFqZr/CvbmVe5EH05aPgx6itAfJCRpGswl5IhiIayhQvuElBP5h3U9a4WZg+Zrei
rTH8w+9qhGz27OJhvKMYz24OSUru6/8t/USs6HhShCYhXOn0V3gza5I1+dg8QfF4GcUUrm3TDSNS
5Pvolinx50+6m5dRgA7sBnZi+2j8KzAjvlGKR4EtWnj4C5/IDLnF6FD+Nyr/IZMG+Q6JHCT8lnuZ
VbOsAGjjF92MCNq4ZSI+k8ewUk1NmCj2VMg/SF58AC5atRZqLb26Zdc4gUAj2NGrV2oOEnL0p+0W
RoE0Ivn5ZjKCgwSap4q5jo8rr9+o763fKCoLHse7+jruZ1PRnbkyN2OQYNxrCVD7s4q7S0JM7i1o
NOaBT5oy2wPQfh4TQxAFQODfUXkhv2iLK/L5wwzSBnz/nezMN28Nm+cSZ1lSpWVa368x4f1gSgS0
dW8rjC96TyfswF3jPz2ISsAVWlUAFbTGVyHBalvdXQKYVO+yVlVOOz6s6n/VF9eGZaREzMQ4b8hj
0xl+OY2ZmIPJYfv2WVw4LUXmfpwFGHt7rVocu/LjX/uhp0ZJoPV4oY60kijib/IWqGbpswuzq5LN
NGqk+dD67NCRsG4qr7q/0mfvSB9+E+3cPag/4IyzFwxdto/FeUgNXHIM+J+xI+sltnQmuLTf1KkM
NZL5WECV01vmvFh9DIRx4mV+yAPPn43kAULqdy4YAeZvP7Ay+zAYRd+3Y3QHlho0Rldh1il1vYo5
5ri8CCCT3lRF/pttPDRLRmi7DoMmr8GeUdeHWnGCdi8pbDa2qkDLMs0cdCeEPysG7go1DTHop0l9
jtOjF/VJfb72tBkD3UR4vOJ+m3YFfmEq+6LCKAnArtvdK8Wbd3hSjTiW1gIB+5KdpuoWNdMXVyAW
lvTdLmrRmyDGzfBqgFkrQx2B1dfrxdKT9dD9RHX2Yw4w3slqvtJajQqDwoDIlm6NgYA0kTqUitjN
ahx8v48IhkSbfHKMyLxI1vzYKRgEukf/BWcflfZPhHb2iXnYkjq95IXF29flsidJnQiP85YfRxPn
k3SaWeb3CJ7UP/51FU8S7ExzoT1C/8r3Mfof4f0Ab7BTDYcAJLtuWnuesNbZi0W0a9t2vzdqowss
h2XlFySiyZqVHwgGlgPziBmmfYye66DdpVihnortBtKxLtK8Pr7nED1R+DzEFca5rWZoV6QFMxzx
JqL24OBoPnxLUKF3RPZ0Tg1Fud7pTu6o21T6HH0cKQldfvDorDONylyKhXmBv4xN/PYIsyur6PKf
8iDJ+LHDFgcjrrR9DqdkbPf+aqKlXLrxMT+yHUtmRrTpMjov9WF/rrPa5NG3LgiqPBHuk+u7XgTn
QSLpfVpj6d52Vr6GfMQfpyW5WxBHPuJnb/NIOLFNJqUN67NwlJQ4Sqah0FnaNJ6mWBqZavs0T3k0
Fsb63oWPKFuk5O21RTM24Ox4j20eKWUrCkJ7YQhuRaOnjinwHfSA+P62GqWxfGviurieGe7cgl0M
lLn5/949TQ5CthYFGzTTptkM8G8katU/RQ1q1dwigX+spe2tLNyl5bvwdjBmUYjaHBOjWkVatLLw
AA9sMuMsg5SgdlyhTk1aCl5GqKzKCLvEzLyzxg78sPjCm7aQ3xlVxRJq/g4mvigcP2DUlvSHcdok
c9D2BEtiDCubg/g82IMdqM/DmpUa2Nbkd1UkZ9WmQsBEwrr4l27wznMmJ5QXURVyhJQeaZGfjqRP
GdwsXPfEJYMz5q97P6NOowCSsaLojfTEBJVUpnB3Wz5qfbsp9Fw+gdvvBdSdJVawStKyQ9zeNHZM
d2m9ogYwK8acEP7PpeKb76jaKUU1Lr86NrzMh4fcBIYodq6zYT+XamhBzK3yEOaAMYMg6jF91yav
u0YPdN041SzuiAnem41e9a6YmzVbu47S4JmMusPwksO2In3ec8RxULlKFwyWJ8+BKdyy5mZadnA4
iao1XNnaX0I3wFeggI2jARQyAEqDs7smJO0PyGTnGwOwMCWpIlM6LvOG0+E9P8vVNxuTOcOvF4Z9
7QrLQhBGKcjE4HQwEPF8NY9IsqQX8+92sm9T2GY+Vl+yBmJnbXWXhAQLE6Dv4cqHD2qml8c8gE76
zgsZgUzM4ZHwxxrKrYyL8gPX6va6lBXZHH49BnckzsPyqVjyM29K3Yxqz7w3arq3Q9e3hSMIDlzo
DjbbFz26kZvARB4mc/WCzSaBTVMNCCHVsZUfenCtOaouQC48U6th+ZpVzXybeDIh4QqrLLHImdkD
HOjuqi3bI5Gp/TEurD4zRxQ35kv2XMfNI16sfvda998lOyALsneSQ1xewWirVHUttYG7wFo5zysS
qm8l0HrkdOnqpPdbZLtyXgnwaGZUYCwYdsfJLfjssBh3UVt7765GwrL2nXZwcsfw7cR9/lmBxpsJ
wxXb9oCDiYqEK/N/WJVPmFFdO0WtV+uW3QsoflaJ3B+eNFKCurfMWPnujopxO6vUfGlLtTA3N5l/
CJoSw50r0vipvFk3glwokOHH4LuZc1kvF6hn1Enb51GIddNgIzl3xOwynHg3nQv4V2kM8DuuCQ/q
R/aO4bgSeInD95Fql2Hk0OaYPRsRs2btHyUwBT12y4a4x66q8NcmmATsEb4ruRJdHZ41tKpkRAlK
FQ3n3AEcz7uQFEzSQcneQVKUa4njU2YO3FDyUF06gYVZx9NABEdyGg6sq8PIqvU1Mp6fb+0W8B7i
7rABz3SQDIDIRovBrAlC+1jOpyLW9bungYe9U8qkvN5HwdVhDMTcVkwfaEbmEEXxVHe3NHMrsVvS
ATMaeyjAehAtIzPfcuAhkj7+b+RXj3bLa0QJuj6rzs19Xz7megXU8ac+fEoZXgMOZfgvvT/uNDOn
kAUXqXCvXJm9lNwL7JCTO3iBVSWooXbDVhvTyg+vqyY1PmdgnJLdYRkVkeWZhRuYrqq+3LovLl/0
M7uB54R9QMolf0JDy61VapuTkCyGq+oKgpNwg6Cno7lRNIMQ/aJYCTqrc9wgYM4bnYfZQp+OnNoR
vnxQodohgQ07mXs0WDznKxn2l67hbv5mCMFd27iEAQtW0FujqEfD8heDrLJRtM1ciANj1mR3lg3a
bwJYyuQcoPUeXYeQx+fWkSA+EIIMmH/GTLd2VV+LuHfxzzkHoAlrmwt0wS1oP4PT23s+LXBlg4kb
HwS9YEsoueeeSzk4DOi2HJm3YleJmWzCCD69EMPT4k0p1bnV9P2nFxjuCLKebXArXo8rTAiFgSEn
ozxVH8MNSg82+hZPpc0/iGm5ZPsu9gfF0/chJYXPi/Tfgpp3fDLYePS3HttT459Zrc1q+ksnDv2Y
wJ0vMvfJDd/xhMYP1jpNISgAA/TJrz5QybtQ/Hbdsj0OnRXKvfo5AAd8cqACxvSyza0XUKwVD4Db
udalTw22DMW4KIwMqBKaNRYkrUwwo28AVK3iwh2HZN4pI9pF6+YZwwVsLHMKAQjVxBFs6pi+jG1J
Du8Yah+rlApmKlPMGmFXKgx2nM45S7jeAGasvusyeu+gMJ4p1pkPMXlWcBdPHs5ve7aeNVfArwh1
2RaQ4iYuQjCadEaDIxNZMJ9DilMSoJOsJyR3/LKY/9q7JzWsXYMr8AvYldRyQ0BzbEa1T40mNIpT
rlI2vt9LA/o4dXj9oGM2ghFUJlxDoewkzp75tc7cE8MURpvaNjDuBgKPEh0rdQ2WK/mDO2lzAWcx
Rm+GbUBOzmDU0GtFo8djfPDe+DgA/aFnabaEQbBnx0AnGV93a9h2OjE/sWVCl3PUHJBoBYVuyb2S
Hqv0Ck0rlz91XAiVSL/zVoB3KmVJLKEamLBPtx6cjSUw6zCyq3Ep0yy4VbFMWNBrvknulc8VuhB5
CNGMUaI3RB1a+5IzhZ+vyg2yienaTtONDqSmLRDBKSj0/izIE2TS2AafOkOAk+Crss00fvigAy+i
6iMBlg/MYEb4hhDQ51NYGyoRpOtus+TJFc6zbsBYFKd7Oa3ENrn2cjxwS0cOgbdRfVKWZr310Omz
3zj6GADiBwigCwuTFxh5YxNmLEN0YpVynI5mfNQlPSaEemUNJymNq+Xzhf/xi49tJaOWqZURhbLM
uuHpQRWm/dVLjL22Z+zUTk2wZVz6LRYsNUfn6uQ1HgjLD96AWTCeLFq/kevSOe1aJDQhpBQgutKu
Y6UC8C1W2T91fb7Jh2xXyuKTS6eeeSPkw7bFPtk92W57gItqSH6bv6k0s8gPONm7vacs491ebd91
J98DrEaB8ftGZBT0/i+f3zsEMnEtPUZGT1fWlDD+V2QSrlGJAso16l/5iQNuuaj5kcIAfpD/hMxe
oXYp+iq2VySD9ybvoLWVGBjGM/AmCuhoK2T3iSrC31Ef2BjMLeAs1aRNehILtJdTEq3FHSUuMK3G
qyenUxyxCzAE3HIT8ng1p/oO1S+zQ2/Ed4QrlnG5gZt3o4KRQzvcThR4/Hgy/bdYc4JMIFA1ZMAe
9M1vjda10oa6sUXFYRygfn3lz/px1NyT7cQhUUjuX8GChkvU6nlX/kOqjrjl5NbBt91olM3NLDaT
zjQbARmCIaJgHdekHTO64KHupDpLZs4SbiHJ6v9lwbausvPQqvA0Lqv96n64+9K5pc73klw0CzUJ
zwJVN/n9DzNKX/nxWBlYtr1mhw25AfeSp75m3q3+X0yKn31vwkRCOenGEb05ZwSPikavTfTNp23H
/7u+Y8BTmV51BiJoYQfRJmjcxGWYearyd+51UN47cej2kUDnjYQ3ELlPAFxnqWUwcujHcox2GfBX
OpZvWlvcwfRwPYJ4BxxFmetOq2LlElePZfpmua6APn6mzva4ADBoXsNjdf5xiJ2FQsr9m+tDPA2g
MPrdlOUBsfu91HNgPYjLd9bCMo/ApGCPKpD12Ug1WmoKBihKnxBdSM6YNesIJqjjT+2JQYyOaiyx
yxeJS6dotSj1KcpCZxGuEanO9+S5NImQTVwiKWPp5z3PZJdADpL36sJfNOd4a8blgNhZefTW4g2A
TtZWKdrHqxXY1b0PdZTgkrHKZriswncTDTNmtc6uFdyZ5dtqmDE4OUjHpaEETOr07VvoSt8tJV7V
gOT+whrqrohGGLJLYjQh1G0P7aB9xWVl9Lolp0O30+WYMW5koMzYG/gv1NVMGLkbG5nIjjRzISvv
gjWQ0K5bB7IgpHpvWeQfYjsvJ69MsEjCtq16QHZs7i9RDDySfva428CxErTlPVndrqhLC03kTFqe
VTwkAE073xq/fYSt6R9vVYpgOfGGicXneie7BautRpNgFNIzbO2RcX5TcNgR2wwdq7lf/W/zN7VA
nRhX89GXx159zRxVHb+DLajp7MmWztIoDRnrRAdws7fe1NZmZJtt5o/SFiv/JodC/Jx5j83HaQrs
KsqaK/RIuNOpwce8WUTxtH9JW4NPfe3R3L9+WCMWE2COjUIMNuPWR674afgeD17VdY73aeOHF+iI
pE6pI8z7pIGZf4a5bpwFSp0Z7fspYuWmolQ1KSVdamq7F1xKGNrzc8rWgX5c+UzpcFKNi8/cEnjL
1DFWt6vRU3SQ+SC1iGRhHxYgblH8e3CiiHHnsf7jsEaYF1R34/uRGyntMkheKvG22X77k7bSBXDU
3yyrnMZgOMBxAuMwHkzEOXO28mkUH3wV4FWPeNivnuXj7bAT1mLop/00bZAp7H54pYB3bthvL4hw
ks0AlDUI7mcPXN1aQ0J98VfbIF2Gw+2OYKb8OrZKZ4ELiFRlbyPROrokyPTvEyKd/6NJ9sDKp74j
qI29O6ZRaqT2rdq1vL3XlnGdWIxN/tm9RXTVg8D9dOwzNFIv4+CQieBQaaiFypXEdx49SLj9YlFu
t+1YKF5LWgcRGMRrwZGJJI0P8f3K840+wx/hTFcaCbq4xlFXIXBKXDPzyNt7MsAXz9Nca27ccmhx
dd/Ec+fMAhYkijTze5+fpF21TMI1xAeDXMUvu7FV9U5mQiGT5lz3HyZpa9Y/uqsNU2UWy5TtsAHi
Zngl987DfTD7Q+b0MMhZOG/Tnh7/3dthMy7gadlgsguu6qyks9oih3m9pKNllMucpt/vu5goQNPL
lOo3isjhGfOY2amYFxE+zxbNnNnIAbKE21yPmsC4lZCSzbDcmOZJrhDRiM8drJq+92yeHts9ohq6
Rgtwy+PX4mZ9gOT/cEH1T8kbRL+TqwQ68E/dd3bWL0dLtNcYtgx7iZP/JJxGdKjUidievtiGo3nK
sf/2HHmUYCD6p5tQd7eRLBQBrhJM1toAIi2hWGLDHordHpq1oYGP72uimUwMpNDK+uBUnRbWPBfs
FIos8lUUCkcX0y4JJXLKgWNWraobPMrRu3IhCvVb3xrJfBsTw7jDrTaDCk9CUOkcDd0Jq7uKOu3k
sVnouNajOXbsOnFqBpwVC4pfZtDcVvl6seojtDFlN0XNtZzewqJ30bqg6u+pq6sc8kjRt0SOU6st
d1hM+Jv00E1jYFwTi5bXrzkd32kkKBwMpPd8fNaSG5guI6FGROJ3xB9jcju0X8WTCwKyBjCXV6JC
8exSIoweqENZYi1VYuzhLuZuSZg+tiPEaruui4/ysZwrpTgwDBls+moXrXMccdvsWdLgTp0ZG8Tz
WBvXlzSpl5l/Xnqkahpl+OowQ43k2KS35rIxHdp8K4TRegdOqvMauExDeHuz+e0Gh75p+tCC3LMg
933dQq0X6iCPySRNBZQEx/XF0tw4Zr/ieBWy7VyhyU646WXEqJ9EVByUsh68i4Ng2RqYzJ99O8hh
V+OfSWvRRRehg30Gxd3riI5xs9HcnVvY0e+Fc65n/JR+Twtf/MW6dZp6h0ERQGVnfzwJ1588dJiw
I54utkT8DQrwotLjYcwilRveJLjGVyGM6aduur7XdyPaB2vYXjmQ1MlqseFjSDX4A7m0JJAVsH2Z
GubzuciACIh5Ja5N/kjoIm6NF6VDUViTpYyXyXPyNweoSrHEIo67QxlWrhRigWvfN4QueuHpMPJH
jeevr9q5kLk+SB2YxvqoDZ+0fr8ndcTF2WZBR4xovRkL/6lTJ/kdX9AoU7fpyLR+OAfYe8QXSg7h
LADVEZr4SVTz+Dqec5kE+en9qM40zZZA2B6ordijgmU3wi9WelGLtkjcMZEEBuOKy68NWBbTk+Gg
nYpjQtM8IaK6dWZ0Y44paE1V39TiA1bHSNtYXbXyaw40N8x0igJJKKfoMW0OgOsB//Z5EbF1cMHV
5UYXKdv1886QdxA5EkfPaTUAZXOCdNpDaIBWvFNP4m2OGLg189uYM50ykwdkcw+ftyF36ves239k
mCNRgi3sj2jX4h0h31RtDbrE9eXARWVQIij3TKz5q3qvhTHlIZMFM0S81yXvbhCTT/1c4mOcTJyM
sg6JVhnWkPwxCCQjBk3m1pqfE7cTaCMIBF2dP2J157P1Ks7jwatE6+w4lA/6iCoKC7VUdhUDjLY4
yHJ/9vQXaWrIDisF3gm8zqQURAJb0WsVZ0QFam9NC1DIfJhm2lKXnJnKc8WCdkbmbXoGmWjxbJOW
YqknjviLHT4HsKafZxXTRawCO3I+Shu5jkyuspFxC2D8IgXYphSGKZweh5UhcRyV/7QTC18LtHxU
RnWexNc6o9/eZx8ZGyCDw5Y1KYcxS2OT3JqlFclj5v1l219TM1ZQnPMy+r8pCdDgkSVnYbLP6EP+
CBW0Qh5Yrba7tMUgjYvGkZP2zNDn4Axj6d83I+FPLgPJvjQvH8fDHCoa7ViztyXU9PAX59Z2FNLR
GQjweVaig9x3y+lBeJubhMW2aMP3gaG/x1EOaoHGRgUI2zvYZ2rHifwpdzA6cAyVrQJMBfDxTvVP
9JLH6oHlMHjJJ88ArR8XJJ4p3CoSQznFZq6pG0DT9adXAkMTm4TtJmYoqeSrSPK4IRWp2mAVtEQP
KfRQJk0iJrp+5ZUX5BIPsuETOFav8NqLnDR5uYXR3toFilRbXy/k2UaPo/aaBusGaCrn6maPVSlM
/tItXKZMuZ/F1NuByre+qH9wl9Lj7gxqJMeZNPrpyG5rqEUmpsoBe9bJPKpp0vSD+J/1Ax3rGsZP
Kfzbi/8oudEQKm4qFpEHecz2wUeIcnr0UCzqqxbyQ1ZbS2FJ4ezN011q9EROk1V1l31M3j6piwQp
BU5D0cbZSUPOeVGcVW21wwUdUT9/cx+3yfQItlgku05NSCX/QP+dk2k0SemSArSnifQamQS6Q7HK
PabpS9UQfQvmRmHsp1tAYYx9qrz+/2L4wqiNCjkCb814I62CqO9imOiJ5cRy8jaGk6Dq0iPhpRL3
joipdiK1ALgaTP+3Eli2JDKOleCS7qNxVy1w7n/vqI+/GTI4aRcaEjCJLH/Ohwgev4BRFLfs6JLy
86EwxbRtLQASbFEY/mg43Gg9tfbWQJChl7mDim8lcwwlqNi3uPxdT5OysoliRst77JW7HRXwOy+m
fYU7l1ggOxuKRNn4x7nTlrOLHVXEVBLYshWFZYoKSPJmIUQqyrZnEMGknNOO1O9K2vG9irWpXxlO
a5zI0se2Zr4amVzF/RYXpVenJ2le+FLSk/GtfbCs6xu7Vtkk9fw1aaCJHWa9xiVou/CXVAn5mGXr
kEx6iAzpKjgcQcF5638gjLRePI3vLBG9HpLkpeSQt40L5sTlVyxSkt/b8DbISLDFoTAFse3uDliE
bXqmkxDT4qtRhAAiMTnp3qz2gPmnD3hL4LQPQ+yZnR+myu9CZIsyyRpc3xMRCiLXQJW46FMi10O8
0SOvY3OaInBAxHAlhGOHm2ilHxn9THA8QSbjHwINk/LeOw/fFb/7xHOEcmv1hEGYpBq5vJPZrnzz
oPxjBa+6RIDlAJgFHW2o919WaFIk/bzeZxCldObnO/igY7qsoltj9Ygs2ccOVITvwFUFIjarnKig
Z8wcxbOHxY9aFBzf0bss/4P1eBQNABoQAXXjl8BfY3BWhvfhT0za396UNta5oQiFgya8paEb5QXU
WWfAG4mDeTIY4EZrwRTmtosuKdgcr1mZJAJOA07dtYMuXv3D+On9+55VOcl2TlqjIeI7BwYIqHY6
hY05RGiS2fUkfzlJB1Inm958AZrO4LPQI/cmqfq9JUCEXrAcEH4wzgbQIY7UgHkrdQyzfOsumv8/
RiCh3j8HUcXcoMDfkRHEZLQ+ZTnA7WfV0OaYUmfQxxNVhtqLx1SgihPpP54ppqY9fwiOw33E0h8k
0gEYFZY9i4yuhcHOYAQd51ytCuE1KCRfye+vc60eKJtbaRhmNmFHrYRL9jpoKgD3m1W66/pGBgcZ
YRE1FDlog9ZLYMrK7dqPRkfsn3z9ssGH77veCyzDOGKtCk+B5c86+UAuIdgoGbGxzKQA5IPmIJ3C
Ns5WL81/IJNdOfwsVmeb+AFfq1tC4oW27M3K5bLPJHid1rS58NRFBPVTZOT0By7vfDvbfv3NBUVs
HpG6rPUMiSAonx1EU2l36Yhhb2Jcnl1yF5r3WGxcbpnWm7Mkt9bumb3cIOzpvg2gClbfi4/h58e3
7tikmlueinJlx5/CnFv4AQ+kDDePzjFmuUsVhr8Q1yFdt/DmgGRkAhdI+3gVLrx3xc/c9qbFQf0e
6C3mnH3Jq9bwBsyjglYzcQHWW6ywhSjf9z23rBMyuTjg1rgYq+i0JyZpj+cHbZ+QFnRMg6E2nDdR
0bdzn3FEpuWuMV9vcqGcL3+nMbSLi0h1zIa07RU7M/RAGewEO6uOO0WYx59B0qGfsa8fERj87jpK
DxoDhizvVkaqjdg2ZMVewG9Ic+8F1T38gJb5vHGWsxZthtQl31usEVZWFLx+6+lGDOr/4EyEmeDV
U/JWe4nU0onO6Uz+NXpPDLQPSVzwWyelIacOJUHK5gvmUKoiHymFlxnH6kw5qJoEjo5VTe6t0Ij7
TedaFRwBYd+i86fT3X44I58jPa1HPrtFR1ZBij7NCCSSKxmiCBYujvtc2ymLrud963Zo9QBCG4e4
OeggKed131z7aQ+EvfWCQ/1qNxzbXWPH5nG/2gEls649s7mnWGcJOZlXcLiuLLKXthrUKOV9P3Vd
5tA1Pc3jLLQaAm6J2+D2khyORqRe4wHHoigCepnBnhTZ26PrnPaf+gKcjU33lAECOTG0zt/rr/Zg
ewFQYSLKsx2ZJrcE3dquPToGDbGZ6gBxkQbz8yXLiZkE31VaEtSo3v94Qi+KfZAy12tu7WItesRb
uyp7o+YLMSZ32dgu4cHQ4wN73DPhPSl/ZqmYhffCouvnyXisCpwUQQId1CEzJ9Al2HYAwDthiHKU
03x1989np5K3GxIzuGwxhUr8mh6XPU+ivzi+QH1gZuDDGtDUBH/xScc6cE012E8seY2QP++U+rUR
mvlWNiFhFeU8Yyk6AU2V65TirkQPK0q7Ne6CC9YLCxbmykaRYrUza1TUsCX1xaKn/Kj/C1Zei4H8
A6fyo50qsD/ovVLUf5iMFNV3leDSQJrhS+P6qInIovEqQ0XItUgJk7EquIVfmYqYPYxhvc1HRRHP
NAz8+D++U4ue2ZLn4VN8KBv+fDA7KXx0XhKCd8OAGpisxbXckbwbozhEbCCx3+JvBMLg3pJhVMFz
dBIoUp13ipkVPSV+bHNHWSkzWQqXg0H3N68D5ObWCKEdw5VUI9Y7ngzVoxO+kQNju0yx+i6BTsuN
W7o0FOshMf6DRK4FGUahqbz6foi1gpUl65Ve2nHnt0HzxlNAdbsvfiGRM31dcikncUPxPcU8veSi
MzhRpKGSKXXSPo64GjoPLIGy6VkPxvHsrU3rwDGWBXB56FA5c+K+pTDfvd351UL8rXL0+5asd8F2
tn7SGmAW1inGsr1uYKvShlVWjFcY4szpKbnTsMe1rlVjijWmoI30n1nary/Z9Y4yq06IugGuNg56
kYOtQatoKRGRs3pA6oGngEHddZgBNpQvKX1O/S4Nb+ysTZ4AA/LY0nkr83uvtzhrVaePfONKAlID
MT+7uvZzYwZPPXGG7+zYmI5g+7aE5HPIXP4vOE+hfD9uzrb6O5ODPQ98RZjoddIrS48n6zzIh0cr
wMOX6Iv/ByM/0Cr1XoRSrlJggNv/o7m0ZUCrOgm+//qihHI8ZIUf2AiIs8x7g9Q8tQc6NykSFpKu
JdtqdlV0DdFFztrVMCKdFfnid7aM9wn0r6+c5NAnCvMiDipyILFTjaNEZQGEXylfa5bHdf1u2h47
F3fzZ99N6fnIwk4hXXDEinPd4wAIVWmT9Oikd3mjLi20R1BQEUo2Lhbl9XHYNAE5/UNl2KZinjZ2
uRWkb3tNyfMbQViXzhLBgK6ky+DwQkvcqAQAgbbrsRk/tQfpc/ZKb3cU54ofQGN6D2e3UcpjWGt/
QHwan3oYgb3yDzRomXrkuSjcpWf8wjoVC0Sa5z3/+ogAh6wLeHnMfCt4Rh73CGB0SbXwJfyTBqjV
jW/R9a95OOHWu5quOxlmhYdhr42C/MbZ+aJumrmDXskhUK96U4YRnYq6eLuNrdQ5lkRYGApPl7/O
OaCPzEa3k4GXOHr7PWU5OVOllUbbHMfsNAsdMhLWSvn7nqPqlbWX1q7wuuHf6mIMAOnCuHT5NJY9
eSX811N4KpQ+RUJkVE3pZdpq9smudPL7Uy/rmXm/cTOUkfrRvc73GxwDYJc2CdXamaFc6dPFUI0t
D4sLFitbZtENcN4x3+h5nYj/4vodZ7NI50P3H4nXcWYznULZJuSsp7JOIPXUCi+80hdQp/Ws9P/K
xNYQvlFBjjekDQrra32z8sd9I8+4BnI+pR9PQmaPSRwJcEOUpjWmF3qM8cVcZ2ahdJCtPYaPc2JY
Oz+5NAauSCu7rLbWy245Yk5bRjAHkhc+4dR8/5bkTEIGABt2LgMWXwS4IMa3R0jqavJP8XDS2Y7t
Ihv40ZB5DSGgUQX/eDNGimT/x7LaFIuDbcxCVVoT6W69f7Qv2fG0D40SsxBmT8vvtqq7eqN7h5D/
bwGLtudPcsaZPbZtYBuUSibgFSjUSspLMxP7rEwZ40YYLwX2M/v0XDJ5ZL1F6athoPlVBGeMhTTt
6/8wu5dH3QTattrpif6ip/JDkSMErZ5xp68CffR2x21pEdPAxJffwu02kkM9Y3I35C6JC6+MLbbQ
hV1uB5I992XnL/FQBYwRXMGwAoestsUVdTwoHdGlw3rpUkZFwiN7FG7wts9eUuoJFRJBMob1y8n8
+2mOzamctmbeAyRWk50j04G3nFl07TlRvDqsqo7wp/WNmzZ0tzm6fENpjkNdaPYSTtwo8ITrcC34
CarSMMWzZQ2vPlm/wBD6mCMJW5BhLtAsOQOlvvIqdQ64zRhSHgSB+mw4jEuiUqsdh9gU5TgOqs/E
GneGspiIzrgy0IUICylPhzlGTK6Ww1icb5wue9GwJ6R2eavL0HW12vzsVpMWZP0by/PPuhdoDCzj
zEX8g46k3GlVAB0dVnrcrmPlFQr3zdVi8iKs7H3cBgW3IMiJ2q88dv2v+n4MTpjLaH7pZZ4QedzJ
HZBPvXet/+gZX4qdF/W+uafFcqCEsI5MLCY+NtHba5WX206hvr06mOPDkcg8MLVtI86WyHGCNqgQ
TUgCTguQdA2lvHmHjhex3eHsXz5cKBVjYunpjAnMMHUW9rWKHHtQ/1vIA4CI+ssHnq6WoR+NEfgH
vE7scTJiiBhCVo3wphHnP+qjxm2uFZlG2GixjbIEOLnPvPghnuW2zT5+gpQt9w29U9ujJMMoO4C4
9uJysLYYzYVqlQ2YNMVD58tjmhzTSfNZgvJ6RZVOcqKxQRVKguffbY1ILR0VSERtl+b8NNO/2m2G
DWazcwApt5OBUWgJF5bUEUq5HF9R/nLbhbYdnh525xqvK8Zub1R8nCKlAlGzJ2cuR6HPs0pbLQ0F
gQ8tyEruFnG6lwTav/sqo0MNjlubr506afZf15dbbhLmNmbd8O+nfDQhZNfT0F5M9MoWG4fVvZpu
8lJHaNKFyOLcsm2I/ZIfBJhT0rxO0ovgQPGdMPnGPzLohz2mVZpB9mkr/ivaW73eiHzaK2Ix7jhJ
wGKbQn9fnMhE5XseHVk2d2qJaPKl8EHYTw5B9p+Ur2yLRZq3isZcmy/N/z/f6gImFguzQ/Rtep+T
iDk2r4pVUzYn92STucmwU+cRDIrNeWIT4KhgufisRLuoAkT+gmUVYmoTZude8b7utiEwbeSo7glE
qT4OH2jGo8+FCgm4fEhymzrv7+LlRw0UOaEL1oCmbUxp2M31r8AhNUA6dSGvY9FOoBoCSb6J12vx
+G7z0nL3dUE9tgUXuQB8DUoHrTNWOGSrRL9g6cIyw0huAHxyH2mBrQuryMrix+jo3YSJBE5XwAD/
i+E1hSWSjXofoZAGlU5yMnLS00sXzBy4QENtVNXwZ1j66dpl/WQTLikE3Sxob78I/d6cUb8LuwOc
kuFZLwahnr8tCwY81FaW1Q4wuZbbfHr7AU82KtIhjoVRjYWXKo+ugtNl2Nyy6gpAtQpfytJdg93Z
XoyxZ9SLto2xFpdTWbU2uFEHv4FtYXrbhO6iF3371OUpP5CwhcWalO5Jx47ujhYdxoxls7oNl+xv
WoXe4uwQUIWdIAv76JdByGuuk2dg0veoQntBwJSSYeYFi01yh3fMxzXpppcMEpIhGFRmTzHDYbT3
W9f9+5aOxnZAQZOuX7oe7aGuQQzuXWmH01NtlhGgUldr+iw91ssBqRIh2Ar3OI79GFu+L09jJLVo
9Orq9b0xFr6tgZ7P7Hcfxh170jJj8ewy3TOKkZfziaQeL6wMs6xhdEQ3a2oj8N1TDUjRTGpUv/Yo
93lK+UZETEXmHoHOW1Jo/yQA3cczeRMFlYE8jqQcMIGTKZVn6KsKqDRDeZVozWZ1Htf4gnh6QsQX
6/2l5+2992mHDQsmp8VoiVHmZYoQ6MihcNNri2XoEaDeG7IlQi8a1tG4jXehgTUQWFAhzho16d6A
NuBumjosPvtCIWRxzxxUBkDqhXmRm8XZx11lRNi7eUe+Psi8US3bRQarDk1v1MBthBMaMLXP76PL
Zh1ZmaU/lJvSj/bpSaJ2LEBqI4KFvdd6GeHJ3IVCl8JXsFNLPuJH8jxdqVkLKU2lozmr+zYOdTJg
Q4+GoSUD8ZlHkHqI2Nv528VyVHLEsFRFdn9C9AXiywZ1ko0K0CGLdnG7T8Iq172W1cytA4rJVkBh
+ZwGkvc8Fl669eVMu6Q97VWKIiS+l9fZVDwxY3y+TTPSWuJk6Xai2U4PoIRCuwjWr1yIghmzfosS
oDyBGGUIYBh1jME648aZYMdwmBrOOv8u6YDwxeA9YP+MOdL/EBw3VoWmHNL988z8F9Wmn1s4ELwd
iP5MLlPXlrLoamBswa47n2+JoRxk1Sp7eIK6IS6g+bOiHNjS6Zxvv3PMMSZx3bKMTYU9dimbj6gS
WMc8cppNVfyKKXsB2EVKulwkj0ffLwntlVaxhqkhtDOEM+WCOBU9RE/Ta1LxVwylblbHNZ+aigPo
OsgkqCB/iQp2Cb9LbBHYD3+Cfq1gZXf4bf7ZXYse1AoJTG9M5WqqIrUbl4QSI1BFBOjGiN2adkUz
8I0aXo/Fsx8lCqjPgyoCE8N0bq4wFJQnUUkP8M487EQVZQHJTH2AvC7imeV/U9RwmFjF9NnQP3v8
vW0KKi4FZP7p45fV5jukWcGSQnc8FykQ3s5tuSuxvjN2LMQJl9yadnuMoCN84fUE82RLQRJrN3Ba
WBBtTl7+UUu829hLwevNlZVsZRI2stSiopMoO1h5xz2C3bpfQzWgenrw97yzskr4F/cVooj77f4i
Q6bDZdGFZ4rOWZ1pUGrPxu+vfeLo63M8Ghew+58e9fIh4dERvkZVYnxj0PYMELW44JmVAd0xNq1L
Z3MaO+wpEckfThiiV4OFmIB1sF53OKrqFt7CyPa5GsbB+ufeHH1ovBJhoXfk4Xl3pAmB0jiYB8d2
DjL41g4cWx8oUYdUJ4MmtX/XbskD+kDUIDB+w4SDMUXrA5yisgXehkLdTZ9FiUM0hRNjB2Vj0Chw
YxEQuQwt933uAJs9lEAeB4alb+TiDmKsyVsPPIK5jn32W7f9eFJm+LbyO8ecldDVzi5zqWYnbf+Z
ewkQm8j3nJ8nvbWkQ+2twkXQni457dwfaNFsyQWJCOyE7WGdpOBrdrYTKY6ZQHOG75LTi5P0TiaI
J0WnMgKjRNHeitaNHKaakcLjWE8wiwAuRmItW941nartRjRGT/m3W+9T5yV6vO5cN/g0PvYxhxod
1XA639UD3tdaDs9pxP61wHain6PLCUwuA+oeNQPNoB/n4PrCQ62a/3wx+kIGFa+VvbaXv7QlT05G
xPw+qZ5mUmN0hHfSDdATLJP4JGyb3D8WNj9an1oCzfzqeNJw73gxPded8CFjN6Wl9xGPYoq5dY2j
Kp98tjK/1xlIohuEneRGFVfwFNDzT7ljomJUJrQWQTFPeLL/Y+VLL+mJsiNEY0fZY/LZTnRouM5d
TnUyqbV7mEboZMhy9MwZpApHUA3CZLEzoczzWHtkDrG+O+Fi4kuud1MLmCtACk3Bvrk+7ugGtB6W
kcBmHZ1Ltbo6+2TTZXFySxE8DpKeB72GG39O/6mSwmtmn2hUQrg4Ad7sOKN/HzWzlmvIp0jb9N1q
TpMBqL4PfGNjbonjL6fAp4SflkXJli4nU4YR76VTUScp8wU282gG8iH2oLUHJ5yN6BDR86VosDgE
cfD+C9fPIVsZm2gTYiqAOfU8Cgb3OL48iB7zJPLzihPradry0Zg5Tg0iYlbe9wTpTPasZ4saDDRf
OIBlG8y29f3fMORWySbyJbUPSliAalw7mfcXeO4gQPQLmLkrig77Hjb0gKGPfIZsjKyk4fNFlnyO
72fOI24W45/rVS84gh9RofRWgw6Paed0whfF3LJO5vf0E7Y2Vclly7a/ixxFwK8ZsXZjveHcBAUC
p0CAM/C13Rl3PTXgEjfQ8vuoiTRVD7mre/I0cnpP1IN6gbHJTkcNQmIvsF//X0jq2EXIwW9N3Nfs
POAK6GMDycEaZevOoujP29o+EHVWg5w5cqR7MQZ3LGc5KgqB8OBoUmbMeZr7Dt6OPoFWb5lOE643
HFrekZQctScAgdgUOL2qzmgxEvUGRohhMlFI1K3a9p9hWDqeR+2g7Rq+MusPnid1VQVRYA3DDPTl
VWhDouFJg2kZZYh88CDYpBT2wn7BG/xgWBjvqj+K76mED6umr/UnmJB/oeKjH4mJIC+m2O0BOwXj
ooCtrDQenSfTaLh2xUgHDuoy9dlFbwj1W8CtByTtsEMOZaE+lRciKk8UwoJd3IM82Dg8zRMsG3qD
026Tf6KR68fLEqgISyBmpXQJCTHWc6u0ADBipSSwavi9HvkoS0RE1lCpO47tdagxY87USWxuzZPB
QRuYO28+5gSToN/nJjcE23qG9R4KeBcaMl32pwmyGAwgos7QHGA4+x7wFL59JQ2oD/GtjmHpmVOm
zLetrToqiMustSkuWWcTzidrOfLspyf+Sv5BpgTPQQo9JX2oBRnLjwpuw22UiV/4D0c/He38DKde
9+UzILUutA2dkjDqTjaCnLi9tmTflLoEr2Bh6kXxwFkZVVsg9yA6VIpWj172QcirgODM99WAwN1v
1w1dRiW26ZJWF2MD5tEdoYsLMD/Be9V2KWti7jWR798TN9IREp6TGRiomJ4BX3wrY1LnO029W1Ep
kJvxjsgqHGFWk3V8z63XQUW193uojo1taONeDf53Ly5J9xq9JiW5Z2ZNCUa1gk7c1/LXxdb/iV7o
20TP0N+Rhm2fjae2SmO3RlQcLUBFUrLNVJDv3a9O4Vpr/ODVf9xyWVGq0cZdSzPg28pZFC/m4p7G
psoZixUo8bdgHN5QUcR/ZA4A8uUfzYps0dqJ3ZsAZ/UNBAk0pvzC7Q0nnKF4hkYajuiiszVjZRqT
fUHBtvudVLKtZUGLk58AtM18A0Lp8i7BTonMQPcvOSYbIk1rPgx/2OGzF4WUsgdIWhu17zN8FzfS
0EUj9A9TANjo/TYGyLSJsMDZM4w4KSljfJQFpLr/vXQyvhCjw+WI8hx1WeEHoaQaQqnod/w2MKzt
unlEF5+qiD/Wsg4pmNaqWuozyuqkWQz5mH43NETBT+N64vznVgeuU7SeKMCI9auAK3UGkFE/5fyi
KB2Li9VkVR1xv+MBjOYpCF0tsF65BRUVAk9C7fRMY/ExIu0aV7tUy7NXorlJNJeJ9PAl8MsRGx8R
hNhqbkyTFc90a3+8dyNJODGv0TgRQkGuLZviYQHJwsujwPS0c6cooXGNstHGv9WWRLBRpnk+ceNr
7D30UrpyHDcFUw7aTMwf2ONxU73/hcxmJ0a8XXjmpyHfp+yAa8zo8A8ttkiJILUyrXdhG9brVcqu
Qw8ppwievxlsDuvHskTjuHb8ELY8QdSLJuB7UHDF+w5EQNigQDCTpIE9Z9AsUNStiibEmEKv0nNU
hVjPoHKGnKBKo0bccmZVpPMi4p3FxcLdoD+jQ+Au8y2NSUu8TfYNVsNnFpYE1xy5aJeQFWOEwzZz
Yj6+VYFWktAQAr7ubosWy7AR98P7IMHI/a2aRRQ6hrAD2pz2n1cPjnK3zs47xYbAtkM0bQEFHb/u
nUwpu2PEtCEro3wfhpybco64VfjfLoCcRB9KMbwhPpsYTnsnnVNOmtV5JXHDmF49cDi+goqnR7SH
BqVk21BrJ5hMaSuEHTLbqpAceMUdpJZmpLkcXPEciis8fKErnCfJFEuROwSi/DvFv2LhR2ifxw5d
Zy/JR+dfQ8K3PiWx81ArMW2ifRUWiVpM5XLqUE4McvxD1N2l+51Pv7DZMjt74+Q7Zsaqi77/bmJx
l//tqZXJWsVHVt9hlW4DhSlpIQufHun+7X8umODSCAqePb4Rfj+6UQs2S//Q3BCE3UL60rzI5wp0
haMAdDhWvzwdtQRv92k3KMjAotbSGhCgXJiDGpbQblVGfef4q0aucGg7G143SftUoalt/erwWGqB
1YBd2ZS6r3Qg6DDGWqOWVMXUkNsO8FFXKhVzlfRb2gKA6ovsatnfmhG4WQzXiDQkcJ431auQ3GSZ
+FjbMsjcu5n0Z7eeAkn14B9TcQicxpYmPv+c6kE9OkvOFowZP7bk46J2hSLzXvOcmK6lPWzihzkr
D9dHOhxPjDvSWn0EhKnwMNe6EsnWVTTW8UOL6u+EJpanY+xFrr8lfM+VQumvgG8Y6+ob5zdapqAi
r1jh3P7i8u6o/a6AxeQg7DcRNgCiJGENYoQIMSHPdrcmhvuhzAtb9kEkonZSrUKcXprEI/k1Zi39
k7R+vXS6Nu1qPfFfsqj1C/gVCxFqlYShEHpB2CWkiYRyIg59kWmwkMaejLvLwoizHN6yEqFMst5P
EUP3h1JVXkz5JHCcaaUdiCAkuUqZKdQKESY9/F8r1Jn6Vl8uPjN80oGw4gez0SgAlqHXevQI0Sxi
jAUaqmYtjxB4ID9PGsuzb8lIPhrxN0QqXw8pJalgJdFpuezAkKcOoTZ4XDzpgQeLJmPxp48GK2yb
PZ7TXa7uZinOZAmQDXmrG19eGclnVdJptPEiFZaS+XdVPVKu0QqtVU2nUhH/cOnXhufqfLSqpT8V
Y6Ds2TE7RnEAYHFDkMoOJkoU5wXxo5UnbMBeUQGJrV3Dvp33y4RyaJi/osz483Hj/xgKQOG2dk6L
BA6rN9fdN0RHTu5Wdg4F2XR6MSMEXa3fni3r359oWs+pvDks/iTGJ28hhEdaGdwRu31xY5a4/gfZ
y6gjR4aSnmiafca0/y2LJLSuDVwoa5n8/iQbDRY1MvClrn04+zalkiOiOV8oyoLjVcB7KRrAI5pj
DRyrwxz77EIJmPakofJzy47/3oHF4G32TCLUxEjnEiJVEiryw/oilU+oS+lLDg982MFg8nMq4Lik
XOhfMNQFvlo/4G4EX4xMtTgfff3rwxmBR+a8oP5ryklJVAdmAbhMAIYOFkEfNWJ9oCt6zrhnPQSj
InuvKPd2+V2SQZGreAz1hhg81KYbRA/L8KrIbb+DIjOiJ61s83WkcBiuTRW4aMrxYqTcm1D6Y0jV
Cf++/cor8NnRZLFC+GwBJSBLnB2EX50hgFwLWQIjV/y6sajWlJbEFauBsYu9ItlDpMCkVjh1XPuV
nRoUJo1xOUuO7WLamlz0e034bl2O7nDxkm25p+90urM1gLxuAFAhPL7bNOyeBQJkptXIWM0aAPdH
rD2YwxD7m1nnApuuni8PM9banNagfjcxpTvyxRAst2k5fSzm4MWUuMb+lgVcD7ZMNpFnvE3ThSUq
naKzhMFhzkGGlxHl0ZHnCJh/JAkZE338gYnxXD1TfPHCeruYSR5SqdN9XNWQXLnSmecmI89mqwer
VpFJ7Ba+5wOvMeeQDj2EQQcZ8JL4OgkfBHbd580LxlKUF00Xcr/A9IwgTlGoM+RZt/YgLkm7TCD0
HeYmi2RJFirH73hZZlRhkfBXoBvIOi2ebtEDV1jLEruTm8iEEev1lT7w64bsxKGF3M8ZVKkT1sJS
FBEvv+cY22Fz2zVtYnwCQv9Cz1XNsy0l7nA7b7uWdHOSlIAKM92AX3OrcatKB1ugCFtzrHI7EAoD
0BXmAHLLHZXY0961iYFHxk0qVLwoAhvtEFP/L3d3z7JgdXGoqyXg4zqjEz3WHAUvHkkkOrcQyDQy
ufhuA32bab0/F66pSkOQJTCOMTGWFSLDzAPqP8WTbc1/wrMdOHo+hITijPSqmTFQd2l6e04xCMko
Coij5X6gPzqxeAhsmaQidIfQWHq828D8PODZ4HKiHD/4bRuPWYiq7bE9peS994Y1nvnOZov/HpLf
hG3F5tRj0n2l7ySUBGxyEXo8vwJ3s/P3z/mg2KBxJZ8No0HTc0R4t5xyOMa7zDHd+6fRx9qWXQYb
HW9/4lSNUEGRQeSgKT0OsQeZvYXhBs5D/cTV37LEK9AmWhW0R8Yd8cszOZ4DmZGy9Qi9Ar7RmJ5o
XO2OTg8lYoPjJA3kdpLPqKzvJBTqbPOcML/5mn/ef3Yq08r4t1EuUaZPQ3TmZc65UvPOM6OiuAWU
xSrM45TzQ+h+liWPpH7D2SfzmCJTcy91CRxchMfKo+IsN0gvNMh8jn6Po10EZHPAwfshHQ33YVVY
xTIcfVi8VVKacBnegfLYfKzKixd59y/EMZM8GXvBoKHsi8ex7UR9uKYb27x9MLjXW4cc0rheZKvc
NTalA4Xsa0ZQVx1Ciy/RZ50MjXl6RLRTFx86JeXbbNw2NAJdJqr7G2N2IP/4wvvxP0vddsR6Pu7p
ex8jxiY+fSk2HXSaRrJ3Di/oZlkj+vZjUWBMzECq7abVK9cvpfX4ConKDNPdtIda0lFisYpvJC9l
LN+oeupmCx+JFbR6hx597H/0e1HYdAprAC57rPCH7SAaP+36wLUNJEpKPXGUqSjNvRLlw8lnS1/+
CQNgnLH/FM3LrIpU9WVdiL8794ItPcA6J9n7MuN8rPj2lWvXW14A2qdDXkW39/6iAd3L/2D2kYeR
tM2E7ZrapoXnH6nTVbmmIowKfaAFz8hdwkcPYlRhhCouvTUSrBEZFdOTJA8aMDvuudM5kMMFqGj2
ppZln6caE0OBSmYxGBqNQMasgW5IiWVpnQqpmK0lLaP3OJJvWQuNMKW9VCpNzqqoNXg2UBlG8N3f
qDOEmZn4xVkNZXvxnPnu1pdXr+/II2KN+S7dHTm/ih07pBl8tZg1gqCU+IleoFDfc+3AYuWuH4QN
AOtytMZBmOisuSgjIDsoFhoZFNKTp9vTrjIJv7YYeBkraXmfSd1KY1Qo7i70TOKF/VHbyBTRjnLU
tlVLSRNQ+ahtxUorneqXdD9+omqF0SjkUSQbaSZj3b/3uTJ2smV2sEzLHAz/bh7kqw9JXgSii9ZH
YXUaw46Mq1DFxMebHIT4UINyOxX7oAdhqTg1hGEHzosnMMITm8zhAIAsoCxpDVjqSP6tAykoO7ZL
jMrbZhHULPvo1mdFPuBMu67cpzhFZ1eWHOmPxNrXNz51PLSiCtnzPjwa6aw6lmdcHUjnBrLKjuCX
uN2yCg2keD/J/QRWgNDEUckrFN/C/sSZ/JHB7a8+JIh2NtFSOwXPnZ6oTZig45GMu4IrBDB/DBPz
Ovxxy1eJeOQbEdXmUssUeEfbnIOrgBeoplyXFGzVdbwtmeEYY987L2BFEdCZ62H3E/iBWIWofvdT
ARLxx5xsZtm74wJt1YT6DweuoMOlKnFhK7yFkW8EhkjWTNhEedv/vfCUbEJ58/kib2QxhEFxl3B3
wHy24LzybsSXQuO/RS/iFevbIvEaL6AW9jFnW9ykbQsrkAHzp1HjGzcZZwKGreyjfHevQDWy7g9C
COV/C3EKdKtuMb1XlC58Uvc75rPZ4tr0LSB7KpJiY2zKHcO1jJrYZjZ3L1Xz401XGFFKhqQAS4MB
Q6PBewpFGw92m6EGYWmK8O8sLp8/f+zPp8uizaxp1+JGAOHwgOjjXEnDSKg8uxjhhRYTsGahapXS
U0BZM76nHahXks0TIPKXhgumYjOo+p2FvWjmvZsq4dhPgVKVG9Gcq1ksc+7XJWqJpUl9AXDqd/C0
Q/6KKYbKoHo6Gau4825w2bXK8w/U1uEk8/4t691euheI9XhcN6aEQGewgoc9ocF0N4T1hAQUuHsL
zYYjtwVqexLPVfhzvUEX2zvWpV6533wAPFy3FalhBAXaJi1mk0Tslc6JTAdTJS6583NGxy/ciZE0
0P9TONXipwXrtW397AJ0lAoOHViL1M9XmSZy+SpzARFXRVBTUwczx0hRiogpCdNqBQOMObTFKjoX
WJp5MvmdlbVlPvNxjRki9mujDwg8yIEuOPT7DgjEYQuDGrjqYLuA05bbPGm7vBlOU0cNal0COmhI
aT3i3GbYd54EaUaJWt+q3Z8dn38/6NV50og79z95QkL+ekjWooa7Jm1EJOFil620BNur+JezQ8hQ
XR7fdDW/gIUCost08BfyrcOtyzkr5a7AWCxhtj11uPKdti8V2VeCBiY8jL1+bznCihnda9y0plda
TowniIF4wI+e6yHZYT2zr8zNfzuHzvLnpVA9QAISfNNO0ama1j37GzL80eJv089gOR03M1LRn0/a
PQSjH3xKi2KHgAMzl6eHuXsrSSSa7OYGZgrMLs1wCzAITpAgQHXf2c3T4HeUAkO8HMEPW29GJ/Hj
8/HpvllhT3xPh8H/TO0XSL9dg8WcMXuFssAggCU+doIbcXZivoWYRdyJ+ZvCYQ+OmKluH4GonZsg
1T/QqBL/Isv5uvBqAjHq5EcR7Bl81YSZX1TdUPfMQJzar0PF6MN9xr6KbpbAFmNEKcH9yG5rzYLm
dfTUzYbxqKRPCqu6Ej3zMG6dQwvb/zLCk+HZHNam0dm88RcBC1Sr3FywKAVv1x0z5Dg/HMQiIpma
Ir0pxqQiT8uGwi5vsFEC8azbsNcy875F+Ku5mcSUrFPOlQVrm1iEDAIMJTUBwv10dO2shxWxsESH
XqUyenc4dh02ObWPmKZmQpdxroGr9xy+ZmQnNvNdKXm4cqeEa0tqZuWC1HQYvTSVNIlDkkrJLXWz
uTsm+LP7oPZ4aDAJhllxMdQqQNOJ7SQST1BQO8pChm4i5N7Wn1fEPGbCo2L+mFVxCqQSele9S48W
2Spp3IJUJOMJdiy2yhyvJpNinJG/U1AxTplRLjs50JPOaODPqQiyyVNxi5U3SCsjgGlUadUz3prp
BZhUoulnaQjd7KGsXxy2DO91vlYVL/jH5T6ieaqt/ELWiR/fGwUdLw6otigHUD4xET3Hgnxq9gmk
JMSvlkuG2iz3sxQ1zpi+PwjyLQiWxIXQE3G4VEzYes7jzoZ0pI66Qrs3BOdxr2M+mmw/s6G57jsg
HGVM0004Z3vAapHeCpebDr39+jOb/1Ypm0H6a5+mhJ/PNUZViQOOGnjr25mbBZjaKMcZ0ZfWtu33
+hDrKr2v453CZx2PWZG5nCLJN6oVz5zUVLlHBX4oXiHQYOditq6hBZ0lwMXHbjzgqjbdN3/tJcpo
aw+Z/STcUfg9AfIydNc69QIdYsPwAKQ8ZJOcWXcpJLQ4DlSxLEfEobJfMvZHseLYiueoPw8CCxgE
x6AewYn3flSL4BIf6HK80iBiXVpx2NYlLsn9B6/Fl1QGwhrbA2xeLMuJ4qLg1gy4ZG5QcCEJzzA6
qvOEX0C//97P2rMGyIJNrX41yrmM9yKTE1qacPR4pEFnm/LoHEtez9oHHi8J/ZMo+ziY180CZ00/
hSd0D+wjMhH7DwVAAgeflY6rWDbRjcU0iO6LDORo8AnHIaIJB1wNKv9CQ3lQ5txeRFLKpBwiQcPl
1En/0dYjHhLuINSzrvH71zSQVwBDtBrQrn8Y3Qhok15oKF16gDrNc3hi66P2UeyTVBK2LbrAj6kj
NMeDIq4YNfrRm7BglIrzmUx3w33a+CXIxtqCectu43+mYD5s/HoUjqJHEULuSHRw//a+2597HMZt
M+wV9a4TGFNHQWOJD7iXHbv0uMRcfRxZCBVT89+dNNFsNVjSH7PiwzY67g3iV8HAuw6+1zCr/+sb
5CNON8hbwgP86GVzJWJLEKSW+y59/v9GscicMfFuwUZnp/i1eJpJduDBEpOelJW6OzPVBio20gfZ
dxVDosqHxzbDl71aelMhpTUsbLqPdugvxgnBXSSCfdzC7kaZiExWgzAhncqCwx14+jcYeQiqh/Y6
f4N7u06PSv9IBtTSkoyPKgE4vMpy4C2FE5BObD9ktx2slYutyJTi1NuFJpfSf8TNdTMFzGu05IWP
fuRncFSVMIanc5RoWC2Ws39Lqc9yk1ZFYCo/qLciVm5EClDtQBaYeksPWDxq45gk/JNQ5fMOBqKg
JkcGXoK2PbXd230XRDIWXSseoor4mLjaOxPGamNO2DqfqpWeEoQo4uHZuuS6T7i6p51+f7w5Sdn8
SCztBdtaeDt3ywTyMbYQeVi5Ovxo1dZAsp5+39tvxjVAr+cMNyiBc8CEK+9k8Ya9i4JwwckwEI/q
lsm768wyCyZ9UTbYvb19oT4RFCsX5N/eI2HU7J8f2l5dYBKrkfrys1/xmPyfT8Rwa1sgaqzUg1zX
AXO5hTnx4zhI/tU0fzOhCgKLsw2TNnuraHsYRtnsPC0i6L6S6ka91CoqlVQmcqE4rAc+emJxHhJy
Rc/eK5HBwTPcQQh0q9VGcnVt1FgLLkWNIPK4judj1vWvubC5AOQZiduJwjxKFOUuwyo0esKsDByQ
SUDNcVWvKtTQjs8BbN4HgnGe9oLlEsyvSy8p1wnKf34VfU9lTUgR8ZFBlqorXgnjE+m9D8Xn4w1k
7yWlzazFqjYKSb6yLdJ9H1bpONZYRkKISwPiU7MkupY+Z//Hoxs8gYS4Xwn6TFwEHjGb/3hcpzR3
/WRcU6+Hxm9dh88O3gELTah4l6x0R8tjn9s+nK+vi+IYSiyVPK4bXd/6szsvjfkjTJ0D5mpLDEHj
LFaN5RxIGHXbMj20CwgN/AhvEbBvzlp5z1O2pRiviU7teNlAmtkC69opto+4+RoFvHdGc1qtYmt3
ytC5Rx0Ab/hBjFQjLVEs3BHp2fK6bRAZQOyLdcPvGY+S8aM1GtMUqtXAjN7XPYEuFlR4I9eSL08F
O8ei76SMiKij9RBIOwjuPp83dYJboUvA7/vyEFijLWSGUhm2h1SZiu+lJux3iqk/bZGbWOJvz8KB
fCtV5lw03kdTkVJrujh01qCHZad938GGTlBCg25iCM4I5Fi4hGr7v4RqYZpKoaCIS00VCGaZ6KCf
Go1v4Z1jxCqomfEFWujADiRqmcbJ70ktRgTkbbHfd3DLe9Y1Ye6hdlUdN78G7sv4FEfg+WnBDtbk
DQGHZMyJX5ZvKBA3nWFf/z0tZC0yaOI8r0lUte/t+nZ6Azbt5uXWwwgg/4Us9fLicST+hSwLbwKi
mEXYXFYRoAvSPy3w33FjdULlE/hyvN2BXpjIjCDZY0fqDxJwe4CH0vL3n0PWIUL8U9KDVYrqEytO
8gdEwV6HngcG7ThQaN29kVPPMP54Jfx512yOXmKRQ5G9XTU8kAD5swh225yDWe71vTRP21C5N4Mh
uLmwXUEWtbm0aXro/qbmwKkgK/lTH+yP3HNFrzc8aqahCU9i+fdBvsg/tfpzlFO5d2JiuZKrlN87
POqNgDfodcgKi0tJuNJ8wl7lz/LSNoJcMqitYF40RoRrEoq4/CvO/ivGsxCHPON0FLV40EdImZhP
mcOBAth2GO9WydmMe/u8jz+IerUCPL9aYhKEGIyIHPZ84n4WKTgO7EIx8qN+Z6VSmJAYwVEV28W8
oD9IyXL+bYXjaIfZkyQksQGFnisVPmI3owOTIimuvw/uHC1jjpuNReJ9/AKzjDwfqJK9CtV9M1TE
y85rHm/7bXCRFdrUZJ3F2y8hs4CMEWgELTt/WNvDo/KE/WP1XgSWk/ihgPxhD1synHJ9lkdRYfk/
KXhZHhHgeF5q84TQcBht72ixPKSGBvmYZ+OqfsyyD5X7pJWT3bYKmx1ZZswRQF9zyQgu18e1ULY8
I5mjRUQAmm9d1iQAaR+JnIhCdkDbkHo8+0+04DREM1mLeknwwP/WM6o6TEY5e1yYf84v3m3VqkoW
3X7IM9sKdVwgSxlE6WMS3XjiDIt6VY0uRTpuiDCSSabaC1zTK62aHww2n2bDzdC8+wYYgJjHMHtC
TMJ/bvsyed/PCjSG48HXAZkavNReMshC87Efa5DM+zNZSk/RYE+7xizy6mCO3jhGb71wRDJ+sbHb
eKaXBlVkV0pq/AaJz+fivzGKJeT/QC6ozF1BfnhFReg0STk3I0DF40OhQPYDksgNCx8zzgb0OpO7
L4awRjPbK/HX9lUYt/7MhP0hlmBtSsry5aHD02ZK7DIGcDngY2f0u400NGYdTGUYIzyYXegMcRkq
1LC8LXEnudeo19Ty93cEaA4XOtLYWUmEZNwRy5hQWRKeQe2N95VQgtB1kAm877eCDkD5nXDk7cwb
5oyaBJ4sHxTifpGo51syiKZZ8mNd0J4e6B4RWK6R4wCmQ0BdnNwW0uAq6PmvaVqW+Bt2Ijs9I0p3
8QuF0cC+Mg4TU9zEfuBg0Qvmx0K7SvZ9FsB9vgTVqw/JBp8RvLKlRtE3Yy+AT7k6COv3gImaoQ0Z
lQHR3bGSC7fBp1caODOtK1fUVmse4K2ltuH8mifUKyKMwbHqu9zAHR62z0GcJWOEWBWQPMgTiDP3
kG1hS7G0GAzQoR8RM3rjTviNWkV8ZslsujobNaiqBPZbBaLghmLMrETuBKPD6wsHaffafTYpvlna
urgxpdfv5Y/xRkKgq9UjUUfHg9UznZYEGYPM6OWjOk7oqYwKX3jI52YtA+pCOBPr2EhLYAJMFJJB
vieZyjvXefiYVFsvc9fblmq2Z+MZD8/1w3bhvQiFx6B/AhD/ETUjpS1wfcPRoG1NLfNlGh0ga4YO
O2jfgv+fw/cgQa+YI29cCRPe/jGevucxZzqL5WlnwsqcsYP0kkIxcJYDanc0k72/CzZHA+B0NMPt
RqM4fsXcxcGaAhMkF3/yR9W35BmYlBGg98sgYWOMG1sCFudRwIsTfzoROstWtWSck852RxNU73vh
/R7dNMFUc0jPt0VAXGw52l0DRHhUuIKaKeldq6yI1gzDiIzuwtQjSuN98jDBnZt2qHurfCKuaSVU
/ZGVIkp2SwqjCv6r2US9+DuP/bPjib6yAFaNFMlGG2BeI1j8q7EJvAjUnvjLsPEnCeo8eGdnPO/W
S1gVXxJdfv1PRI+MH60CaIEiVFW4plyuCtrplDIwTc7+JYpyrRlXOt/imPstZ3uxQxBpOOJbEToM
siAB0/Hwej3Cpl3s2C/wQfSqPxiTmd9INRd2CFAvt/ahK6XYTi01h+RM366fK9P+2rxXWOLlfRq+
iMzDEXbcMYqnb3a+Ib0/iTrTA8xrOaQZ+JFemJI+L8ONnKn0QD4J+xv/rGkmlQLfXuLN7lq+cxIZ
yWu1xNofWNUO+XbgWiXm9bz6j6bKUmaJCH9d6c3vAQcNxveZut3EQtImqYNF+9du8iABzBdAuMTi
1onZig5Ut6t8i4NWSyBq72NHsPDiI0jngOlf1u/ZSfrXb26Fhy66Mf+HTJ2GNC4vKbUGc8pWA8I8
zBgncIt7lJj8AYJAE+7pNWDLAFmp022deUPEfZtP7Uh1+o2aNulPB9inn28M9w+CEpzdA4bozrVC
5Ku0Bik1vK5DddJawxOndGHVge+42FWwwEQSW2WeG53iwAgJ/RKAtCOpkv80HnTuiYygCKCFVy2f
iev4VoZdJeaFc6oeZ4biob3w1FfFOsoym9dmSMMHR/UZsBHZvyrJO1V9KAPRY9Tn2XbMsLLmalx1
tBCSwBvzI5IVFc/9SPL7cw39yhDVOzIGlVuHRBzHbkxXd6TgKVqJ3xtKkRRFfzCO0ml1pfNn7X2y
41J6E9PD1cfIu+YDpKBkeTUeJi5yzkITKB09eU+D3kT4sD8WLG56ZUFHZRyAOEUtV5IfaQOU5qaH
/xM3AAioedngnqQ/Wj4TQ/j+a7bp1TJVHoFv7+Gprzkm71Gdy0BkDDZOk63GDm5uzFpRme4lYR/5
ckY9kpB0Efn+yMD407rPoJKIWcITJLLT3hEFx4jKRI5tJ3SAuFXnOt/3wx2OXfYfaKv12bNYf6dv
dd7XTOlruQtlC9ZlhqA+yFZfL7W7JHFksyHC6xGs7JiD8lGRjoI9n4lh8TYBPtcw/HynnrnTfsPa
+I7+YTT8pMutts8e97IgGNLPrHvOrXvtIpEz0PiQoI9B5CxMxCVG77cKtNYi0952TyIgSZ9eQpwH
BVNo9Dna5F2NKR8vRJu53zalBv+zFVDKyrtr9muS5Z9eVAKR0cVhqpjTgxJ5a08ytc9urOBPeBmm
jlxZAKinkaCq3QZphH5gzf96TIUcj4SewrRUfaB8R3lz88XCIBfCiJhULU0Op6Nj9V2bRzwLKNpv
yqMqbD0HQgQZhbYChgq/vsci/8YH+1vgsrd0ZSPDYJEjv2EF1oIZ4sa8XAkgeZ3C9qgaAOYhuoP1
A3hgc5rl5Lz87P+v9qE8oYI6SmWzRDe3+PaaamziXE2/O+TF/nFJkSq3qra608ZtHX5dMfZbIQV0
zFIHfGpNTUbBQOXaay4fG6hhKWAXETDpSDc5zea0IhzmcHyntznHQ78U+2HrFlMIGLMOPj5jldbq
xIMFbpKTtqfG52NkQ9oDlK5eApcFU6OuQK+ya5hkfk0/+NkjZBeEw7aGftYA9uc8NL2O5Qxs7tna
dFcAn9UzLKhnKj2dbfxrRlZRzz1+G7p4Qffo/CN/1Hh3iIZ4/mEJQzhBaaFXf2ZYRcams0uyxksx
DJHwa1SzAakgzKTM9AdU5r/TnXH4GRjMim1/ae2CkxZyIg3f000LPqolJwlHDYCJb00C+wWpCFHd
j0EM7rqXUmgnCnJ6a5cAItaY4SZD5gf0b1MuctH382cgIVZSqn3PIeCO/eER4NLndi34GKMLk7mB
ibQTZ3OgDq0OgtAuNlLsR/F84TjVYiucjrcku/fDcaQd9Nv1iSRP1/fouviS2nmvinB7oISCF9ki
+0k6T+Ws4j5YovU5YEppbjG/xp+QKqptHfROh0LQJICOsquS3f/CnaB/xxFiysPNWh0LcgRmP6GL
pb7JsUyIdTVs+Q8+Q5gp1g0iLjUbE2RT+1NmDnM2GOvO1XitS5/FwKlWLgIlsiP3KAAUP1e1Be1s
8/C/Rej+U7PrH+mLNLOlvMrjNS8moUhUY+EAbHM2+u/DJRjfJCGMilyky+jrI+EHnvXewXkTG7vf
YTExfuHr7eCKhBJUgyjcxdj/h6Z9LEMX/rlrsx8mDSInuJKreI/BIHEHDOgW4rIcBX4L0cqH0FYf
oqXG9nMIvF70BqiQFiFNqVq1OT4YFjOKWbmHfMpRvwhQUWKTdJJc0P19rrg4QZZUsTrrt50DECut
LBEp7eH86GIrCbXS68LxfUy7iVxOfc3oRRV+oxIeqZYUT4wlOfcqQOY7tRKKDjqk9PISckeD8ogX
4nhNC7jpqxozYrUogN4CQjdTuXntN5QKVkTSWoTKlCo+y1TU+lJTWljVK1XXY+xMVirbtKrGkaiD
CCDAeeBA2w+9Psu8PVUgv7x2Ym1uW7jhrKUAtkBDRgE7vmFGiXS/SWbhhof07cOk90HPb0GBcLIv
763hKkDp34UaT30mQcV+0/eYQdjGxmrmsgV9NOQ3nbhzkC8+qzAQONA8jErpTSSRDSNl5LifqRVc
/o2g7XL9PJZzt8FDfViq9TGUq89muHacCBRjoQL0U2KfLSPpnwu0Y3pYOUGpHQqasyeY07538bHf
T1MrXGO8aUtOxlBZRqPgn3drO/pG2/amtqdJ3SxOUl4pJUzS7DpeWReWPhqZ7IRgL9Ut/dTKvpzb
I4nXaKHymJeGhtpZXfLF7nr/pHCEAVC+hnZBEeaJ+CcolUmnhmv0cVg/g8HT8b8HT4BgT9typ5AV
R+lHPoYNTqXTT+dXxwJnBdo9MWonstvVA0Tzah4soumQ0KHJULYHfxtTcdZdhCqTdvM7b0yngIR+
q66F01vSwW56ISLFjnK/nlTbeDDFt+/Y1sojqxVQLIg1l2HVdzGXZabeNjMwwOqKbXFSK4MFAXL7
nY6HYgvnLDk00ZKfvGVBN7ciwsBCNRfTYSa1V6RiU5/kIy9pGz3GWtF9avkKWpIk+AIZk0Hu2Y6Y
jbvk7dR8y4aR10CVwqJVJ0LHRl1j/dX+Twrt7U2Ok8lOVAngdO8ZQ2zeEe+utoE9eQEWCAlooE7G
yMFbv/uuYs6TPXVUGFlelsWREt18ZzDFgk8qqzwh+QHMaATF0qk9aRBf10FvD1cW7JXH7bv4d3XS
hXa96owu453c1dd4jx55Ke508iHEPhk5IPHmUG+0QN6/tQHN8sMnczYS9ImDsPzYLv7fvSoWOS3s
/GMbl2W4E+SutFM9jkuBW+CzGJhtgR/yfTCvuczLZqXL44Ogim4ge3mx5Pc7v6Ia+e+Ezzjk08cp
BTVidg6unrisy4RmQqSbatEEgxMdTtHETUf3RTr5J7M/bgJh3nE3SIj6bFPWM7OYOVxbVPOD8mUi
v1Q40aROdkmZaGZ/jRLRNHaHYZ9PgU0Za2QE4AZ0sRWBrXuBdBtJunhi5Ze1LPTAmen1vp1Ru7o+
MfGb+bhoab++NPRS+GsBUilpxYATdlDdHDlKAoMhwZ8SuXPEOCzQiLmDiX/1qzaPWsgRqjCRxF2g
8hu1ro66oTs5mXJB7ozVd5+kvnAIrNBl++GMyYzipd9zFoqsYFPKzeNb+4lpavx2MbqrRQc4VmON
99IL052FAcm3UPzddWuHykBH1c+drD51EYLpC9H6xm9AqeePv2nqyiGpOAlKfMJ4cUUwuiO75Y8k
rJqXMgXxKBZH0p6ja4iIqA/bEMoSMckYSa/KgSaSa7w6wi+kaaz502/cAQ+9wZAWbU/MA2dV1CJ0
5iNQgq5n9PO+900c53Avi6aJogF4dPslp+kEsgqiEPLnRKJNzGruZNGYT414u3TutAs+q5J6nucv
BMnhP5DjunZLV2bVy8LwFly+4xLvPxTNxUqlRw6GJAyvhhF5uzT6SPCDR2ZXkvDl61rrvFSoQJ+N
3K6l3bLV7sfUBy8GEBsRRaC7yEqxpF+ZGBhyEe7NG4m0ZDJC8R3tbxO/88osIMUGnsBpdaHpWKrQ
4ehu0JwK3F3FEqx/qg7rfRR3IlOIy/qsqLOHD+yXpCjgyDfGR7cn+R2npddGGhiQMU045YxT9K0p
WOam4y1eZxTpdEU3Oj5W6SpI20FRnROLLOq9wGXry5AwmbFtTLeHTJeC6jV6pLNmuocmM3sqbOJi
PSLsuw2ovw6JCrrk2PIbA6uIBHB7NCjRNYSmRAACbAJjJgWBnQLxdnRO/bU1vgGWcAK8W35QWYHd
SmDnAi4//273VM+1u1rwSFrbIE5+Ko3oaRk3y1bN+4lHZht8ZFnJImhN18Lno9zrLuSTn0utSFNh
ECBVCDWlWYNWnmDIxXSw4erUZzIBRlc0I61C1AxoMjxfjRGmIShIk4CXVw7JRZrhc3h56DdT9Gsq
Y2As0u1Hg3kLZao7OW1y9k9YZHR9fMi8zpCsIvbwINZdAkNCDJoSPclJsC4x5NRso5tZemsI4VGJ
JLCvPoN9sjKqCJ/3iYrkB7pJ7eDKmYnCXMaQftekaQy4qca6NmZD/p5If2+nHnYFoMe2n/GIQBEn
3fVYLeq5S5lUqaJgXmnDVlDsQEQxAx+BK9JsE/pxQFi6YX01Y6YoRzVuPT8uGjMOZFMJy0P6Ediy
nCWK9wchv3Zi20k1G4Jyn+Gp9UPEyh3tmvqypnVw/7Erm/+uIseiGFBTCqgdmsANZGVc8W4toEWL
X1ModCFXqGUgF6XqEqZUWhaNRI+EOpiJYDL6rLJIZ52mZYj1gGqhI21DlW08yIDqQHme81kG18HC
NngAWsadvFUm69ERXM5E1e6QKN6el4wBE7bSynLn8QmQDqdWf506ClnyY5LDX5c2ZXSN4Xn12umj
RunkfOd73z4jRt+iu35V4QM6FAuwtdVsUpynAYf6eGNc78OSg0KpkKcIbBVNOaWi+ULzP4tflqy0
qAJIjPYrJTE/7fsZhXrLIvj2Qim+6j9BQX7VqnVY98Ku480TUIfPouyJ7hQUSS45ZecMdFeicexq
miI4XUzYqFCLKa2XoABLBVeSZFFHu+G+s90VKsoDt5J4+1w1zJZS00HkkOVvaq0I24ddzx4fu8U5
ZLgBSg9aiuNT/GieHhSwaQvqQKMe3lDmnjoPSLHBNTn50sQPpGEdVdlH5k/NEJ7+CLfZBDqhjNaF
LAL1TXZNbPfpe3dp7bluoN4lPH7LpS96+tbUtXM39XVj10Bxij6kCd/tUb2+pwxrtxnpYuRjh4h6
3ZGVZlsEqiT6EI4JXTuUaezpK089x3YForL5xR3w7XDGxZKwGdofT69tyQzGD9v0HnMK0oQIDcrI
C9EDBp1fghNUMfniXJ3QuraJBb03BdTxqDNEqolchqVHzaLjhkwzcsPuh0Ono/CDz/E5H1aZW/14
LGzcqyKmif7v56kdlsOZT5Q0vq0R/qflNJC2eB0uuq9Sh7zn/5sfEcmgT2ltP/yQYjeSRgEdvXte
CO4HhNffdey6AqaX9HUQvFrvG0/bq/8unGXAVXCkZTaUDBQ8aaBqW1uiTQx75A/DgB5d2uL5tfo4
uwwZt/IkoAOJDEnvYdj3SOzjeZbculZEUE5KF/T08EKweOVK/RQjcotcHh8uPP/frdMCScbDeyoP
43BG1gO312DIvd23dCFsno41PNcJJ/hyIImEA8EmM1pdevZBhgnE27pjprEElNmJ8Pn6HnjT3T6r
D8jvdYMPpfRau3kYJXeDN0myxrgUttjcaErNfA6oeAyjImIzRkqJzV/KmU8w5UbLWgWXol5OKiEw
wOkw9Ai8LnAKyfmQya8acaGBeEIoP2SCKohsY+wO8AnRtLv3/Y+Pwv+SFgbaq5K39OcY0AvJG3J0
MYn8JC1eunUU758Ls3YLa4SAHmJYqAFCQcWWUNCCu4mEF4mSXVpEhx6UD3SGaNJZwO7vCAKhWgHz
91y8kKJu+Hk+bqIR19Xl9/t+DEYvcjv+1+FzdzbNefBYcZA91qnXn4kC9WRP6Iy18a7qBH+FGw/e
izGR6k9XizfTZlG0wTa89Re7QWkAUb8B5lQvXoBoIbpiLHOUeQ6pji8VKX92T+Pv5x+Wxid4PLhe
9GRZ+Zt7i0FFXE0rNur0TPyRTzTZJnjRBToN4GN5FY9tnw/x72S8HATMZBgdK6ub1abUcUCm4+wh
Bc4e//P/Qi0+lenyCs4a7XZYpiBXijNaWeMVqdf1xbOu6zc4YnQKXyEl/wIHLorLMcZvBLmEuvMK
B6mF4+Nm1xaQ9jcNEZLiS41ciFwbNzL3oCea8afsIIYQ9CRyhgPlbfIVcCBke13OBXIEXpYSp5le
W/bR+W4CFjkg/ApEPrqqLf8jGl3zxu0aRwZpnDM50oW9AnrIaKw+JvyZq2+Mrw5QtDelRgkOFyb5
aENVjDUzpzorXLvMGsquulEgqsfUQjXjzYwl77bC6/ilEXEMRMSVGjNspX5alf457M7qFXV0v0gL
9guWzYcK/BvlobTk2hS5b+y3UZrfj8ck3C45EG0wyseqU441RI8FoRyH+l8IppZa2QgYYxiKXkG4
FjRdrULgvyRxdRup27S1KRmCYXzywaoJKh82xjFJojai0LZDcPoM1XH4Ii6mXcP1F4bhYRvX/mie
jwqWLfIYsN53S04Atldv0GED2FKOvI11ARQJg6EWqynXJgKT4/K1lRxjHZtyXKAgNfzRKZyty+Pr
otoXuII9NrRyAYgkxUcyW8Q/gGdfxXTJE+Wciq06tmud5gQNsTT/7Ue1l2If9hOpR21M4qdCWC97
/Pf/fgCtmUrhbjhp11BJxeJwpNLz7xWT/kYF+sivY5RNDnHXDBcPQf372iIhpXzL4hhOIC7ihqqG
EnAnRfwUMWNoKzOS7MgC4o30qbV4nN7CI3cJnQrb8gH+hIDycsDoY4bCacrpz74Lp4CJlu7vPZ+5
W64XW9VGHYJUXzNXn4ly2iAaqYEJ65Nk1+y8GD8W0AMZfpvZqiCt5gglHEgzbV4Rd2IRkvjQqi7s
nl/firXxITbmfGC5P7cKEghxJxdlZQShh4GFW0cFNhc1WP9UzBMlw3F87CFoXaDYpe1c7KJ+jxc3
J1Cnri1v8pbTNufjARQxhq4wVvCgxUn/+L7HE9pxcOX/GVsVc+hgQgkfFWH6aQ8zL/2J29rzLtEp
rcWR+GhGPvIHGzjCGQe1Qt+kxspn+EaR6NocBKZOMYFgo8tZgtgiq1AU1Qno5sHqjgdhMxNc213z
uB1FLHXEFYhEvggN9Jv3rrvgHmwqJGBq0/L1RtJWRVK4U6bFYRtp9jemZqWnAGXy3Oi3FtbsQOeZ
Cm292PgmEHA6qhwnRD9SqWpYZg0s9zmKKXuEVDFIlozQiP3oaETIIBZcJxzS+nOP5vTSGkhQsrfA
+QWfCmiQHZuusbsGgFIKLyPwuMcOUpifidJj3vh93Rwh4QseoRxMDsJKbRnSX+blyPXH42qkjmk0
j6wX1Q0AGplnZQRdVwsp4/NLtfAPsavXLEOCPWb83+v9/MBzBMRXHuPjQlPe3ro6VQ3V5HyvnWAX
aKniE/BgPK0tqoGtBU4VBlyOLmw5ExOjA78ozCUIx2klSwRp8XFvrgfL2rzanRxly3+0KFOVeEQP
bhPM6dsEUgX0luUPwLW2XEBXAwgYUU+F3spfhV4Q/1MEWrgl8+qTW4XkvNxudioxJWjBeXCn+2R/
6wALrZDPOoL+hj2XXeJvXqs1WHVoqd8/NMQ8Uo0J4XY3qzatHCdkZBwLMMHogJTVb1hYx72PDaeU
k5gNph1NR/qOTYNt1UAWIV1Jk4KhYa8T6clyLfiuedGQSW87AioYlfFym7VdIdY7bbUfCSGA3G8n
ewUnfslPeP+tKxOONmvlJS8GrtAwywQns+7DvaHg6zwm7QO4RJjvZ8OkQtfaHHu4qLYs7kpJsMTw
VOWRGj8c4ujZeAZ4vnkxnmBW1QN0RgCveEtLUaN+AkI1icWB7YF76D8f4xAz9d9jGA/SGRmxchHQ
cKyNDVhE4kela8y1mAbJpg+wHioCyznElJQEDxLtax1iapsl9wr0ZbNc++0f1uZc3DYVqB8kRcMk
TvbhDu4txK3y6Flz56ZtN0j1fJbjSV8Jbps6thIIIkDS5aQcCU0+sM5zX52kW4BInkf3JtgjkZrf
szBfXPINQExnlTtYfAY0e3bCYvYQLFRuVPOZPENrlfF51LLfdqYdGuHH8YTjfeznuqaW1ov4C4fT
KQUxY2kux0w/dXa5dvFZbCWiczv7r7yMRimNgtcW27hagxe2RRNTnOu/gBP4d2MMOvlgV6opqB8u
ZrCtRr9VgCoLGjLNi6X78twVEKItnVDyQ/s16/6aJWxJ66fi7Gmq1HjaX82O5byiAmulrcVJ6T1s
rMUdfr0oNAKAlvgrtXe7FERS/YLK6c/IvU5580spBjT9fl4+nXVY1C26bApdXM5qcRYrrrP1XqM0
CjKOtlePNHov3/K3EfPoYMu0Sk8b/b5JjJningKjTJ6XoYx4u+iR7J1L9x8YOULNhPNgMXcCLpsw
eqfBRyDTWnaZBUISno5mfOlzHcQKQ3tNqtDSPpNuImQBn1fv++sYhIFwATpajnA3G1PtovTC9Qd+
/rXTz75Ew0ab8cJQGQtwrkug1+OwmgKwmFaadkTreodZc3HJb16G81D5+EtMakUSyEiW3SIR7k66
sSfIbVNE/fjh5hGR6JPBumZYX1WNHxldSx58mnsRQYhcHT7kM0Oy5GSnCC7HvnDdyufpO4aKEj1k
mzp4Vh/fVRuyyx6ltx+/3XOLF0q8j8Uy8s4P4LE66AiOTSpG52iToUxBdVMWavN9N1QlG4an5Djy
jLwbF5xOw42oW1tTem9ZTh6TPLqCiF4bg3DSBbYkWjzWNwatD7E0hXNHcTjDVKWg2JOxI3H3l/ZI
v3Q+c8npHsJWu1tQNonVF5o5xWmCIMgS9W3kqWou7eQMaHYi/XgZA6I9oJ45umw/qaUbcnm4MSoX
ht8USxtOPFEdTnuwtXjQ0GpJtHk4FC6Whpog8SA0kREX7zQbrRGDppzcF6YXppuBoacHiiHe4HZF
O8T3DfvhlgnGKoNwPtQ1t3A8gpjX4tB0X0RXwV5pyDWM0yMfU3LXGSCl5PH9CDZTFiB35JitkEYB
oOTkjIymMGm4rTjbejkiDgr+e1DfOIP14lWr5okxTQEg62C/b6tORVPQCwn/fbUlKnI8qJ7UCjFM
yR61pjbjnPoZYQPwkFF9aoBbgq9weanCgWIii3mq3yGRR3LLCI3RUKTEsdkDVBOd8IDzPGrx8Ed1
Yc/ppt2K99XZBF+dHQiE4eeJsrbl2K4+RClu6C0d+57y0lqAW7sOQlUNw2HPN3rD2HkYvbUHQTCZ
g4k/gY5x1mSNvhlnM4RVs4lxV5boHfUmJnSxI/gbf84Uf0gQaqBwWZw0mjEIhUmljnvLsS1gz/XB
1ggYsOzCglGeSlKuAPwfaV++hNuoKhYSwCnLB83x350sq0VgPwpGn1QpEqSbjNSDhY16K09zrRNh
J6aUT7MCvTMxQrikatDpeb9WRNUJRbjeHKr9oYvibDfCb4+4GgsmHreWqgr7bq/hi3QyPekAcrDq
RfImCBbXguXmE5T8U0Y5bo09EUOXFMh5f4iZ3ECFbUbaxjDVY4fHqmrIyFqyf+Xt2FdR1dgJhced
H2SjHASEFFdRB51/v3eb7O2YZTFpBu/tFHrZg2e1I7KS+SHxZ6Osw/PyKA1cMu5ACqpW3OTv0yEU
bRRQbphd0/PeFCCgQRV/bLY4o91xQUJH36jiZrlDAsUZe1ZjNPEjvrR/fJLdP70X2PLr/cuB/idS
8gvlp9GShPCxxel/ftEC4vD00z010Jg+fwqfnCnVySdDBz8zyhFxc23L7dQDI7ECubPwlSJQlKfV
11IJE7uAIzt8YiUDIO9XlZLI8Z8bMypUZsp1Hknk2w3kDZyKDmgXYVuPjJq3LebtkpwP7vzbk+Ne
OpobSArZlrL6xb4BU7RpmVFx2eIWJb2IwJWXnX4uVO41XmMpIPFFX9e6qcjn5q7zsXVnKit8Up47
hNinyNE9fUuv6iBee08Oofgpf9MT4y3Rw3EucdpuRfEVFyAR8bXJy4txUvpPSr29idVut3rI5Asj
OuTkEpuVMldozMIokhLEx2+5DuUr/nAFJk7r6OD/r3MTPFRiKVhjhwLxdZuZOscImEfC49L1yx6f
1POKPwjdiut7Wy0FdgQJ/iE2/qLoo0+8d6C1ELSbGZ0PBxvIS2gdPKjzSHBhx61OwMYF1zww8Am0
kPHIV/FNpmpHxcMQGHrURuJW95Vswl8ehXhT3Kv69o4cUhJPIIk8oC6BdT0ZslP9zTNTmJHFeIlN
h9MjOt6OyStL+UxCRoL+Vp0XGa9S7Bb/oBXshHkdmrTnK9W3y+yYhuTrbapFgZZRjk/nswJapPaD
bZ1IATVNY7TrEJ0COGrI6P5QHD/4VDDAWSv1C2OCh7WY+fBRGkUOOZfYvxHFeFl0hBgYLa6E44Sg
olt89mD1KoFs4thD8KdeA93yFWiBy80fWfJ23/xzsDSn1qnnXza9FwpznqVgbGuLLUA0fRrIt2lS
S88uTim7dQwZdbp9F79deeh69wflPP2G7cM1fHQBe+0syRAamIGyNlT6QxmpCjoI9bjbHE8E9AlA
JO3bhC0EyRqaYnARt/3czlsfh7tmDMOuhtFAGUbfWi+syKI6KIAK2wGFi2M28IxehVLWuESDtM6G
kfzSwMH6XR6D74fcVAvcb8+OzoQckzwFHHRkjhfFQeQNvNppL33vpYv0gJdc/cLJQYXk0z/75qJY
x+SJvQnDdXS5FQ6XjXt0awJwd8d/AVlzsf/b049icM3K5dQ8zuYCAE518kFM+yzXtcS+Tdoh6Nyd
Idq2c/DSK4FuYy7Eoc/DR6F60DdQeS4Dqlw2GdoCnBP39brrivTg4aI+mok20Esq3Pv2FtkNuPWd
DVwCcayjm2RRzbKxu42gKKFL6kYof80YLXz8UhtS4EP0EAup+8RYV8HoQaXC1UU+eQ3zAJzLFiV/
CMYMWz2OTDJBDFor5cjfbKDDJItmn+Ay9VjSWi1LdX06J0ZvjFjh+HPbpucrebScTKaGXlYX/2FV
BX25R3E/c+tUUifEWfXjLmOWtzwEc3Do4uBeJvvEr9ovxxGciCOvQ5ztxL2UoC5FOa1/Kug9Tn4E
VBUpUbbJkMzj1RRXUu5z7buoGtf1IkZvVvO7i3zMdnKgkVo3pFY06fqZQlrVVXpwObun89vECteO
LbMJ6AoDrMsGmv9DAayXiyNsR92kfSFbYDwNw2FpWCnelcayoAGKf0yJC6Cd95RvitS1UZLIxsHq
nj+LwMiOLMauypSQRiX4s3Mm8CfmpQJMSix6mCs57g3vYh5eedU0qNYMmBT1EPSQaapOYxK6HMnp
8SYEhg+ZrN4o4mOnwGcMzFLWjL2dx03KVADwxPE/KqoQLJktyN3oT3/OquCcPxaM8a1ogUSr3v+Z
Y+WCvq0VjOdvWquMfxEVQ2nIz6NP1hU0s3ihCKXORMQiu2IGFJPUWSS0iqhslKH/IwFmOyA7uIod
ECASnBXfPj4dusJGrvUxzPGLfhCX9A8ZW1f3oaoRjeDLPDv4keniNDdpKM+dJ2mhBT/dSbZAMqII
BJEZK2tLTKYlMs7KWUegJLAzG8Vfz6JHX8CdqxPMb6VixYMhpoz/0wSLWTi5vX4cH4qn62ayehRU
OTjf1kSL+HRRZeLYu71SPSkn9nbnZ17XEqBBK7pMcNzGNRkNUImHatgDPCfMHAURlpzoaKsl9JbW
FYt0MzHtRbQtz4NRqJsps4zFQYxhRXUSSnVo62OsTUl5ZmcnLGtOxg/roECO0mEtqGda95aWnr/w
3dz8UNB/N+1+RrMK7vS8ZNcQa5wyNNE829mykFWPIDkoI3Srv7jli50K2cyKvb0U20DeXSoYvO+U
rzdYMnb08sbmMgfLCgOHw2xK63mYQD0RQIR4U6zuF+ey9DKst6+P32l5mIgTRnYZZ5+NskSSM43r
XHFBlmgLroKaoHwmqD8k8XT1iD/aN7/msEDRwy2AcQztDxp98KyoeG5545piUneSOe2sm7eHiENs
Qc+ckbMTKJK8jwFvqqIPO1PwjlZPbspbl3spKZB6yHUkZcbl0ox10/oBzHByuui46tojuXNzQePx
4F9rYZcBqKxa2bnaxS9AEgM5fVUVJ+RsI4wsWzW7FeUq+UanZUZBh5qZqKsSz3A/D7UKqt9q5t/Q
C5hJHq4DIrNxK82yYPVrtA2GU9g2NPNR9dYrz3xOODvVn6VYwHxdVWxBehR4B7J+Vd5O0RyKrAax
USyOQWYdERjmuTpIq7q+ueSTKu6Gw2ZQzoZLjwaD9x02CZasEDJUnpAgMYbQeIZAS4r+bJ4BMuax
NA7hlCDOkAh8N39PphxA+W3Q401HY+izc8NlDIXBAdGZp3L3tWQzB80H9AkCnmD8oN/k7ewmj29O
N690MEtyy/VVIHD2UjZ8M3rVsPo206mLvG1j6YL2ky4msFu7DKqP3pWgIF9qoCFsTiJEh4bDk0g0
hJ0vZ5TdsuOaffOiDZvs/w4gkMv5rSsIrIZc2i7i9esOSFoXxRP2wS6RCdOwmA5e8fEGC1SFYX1u
SZIxVAJy2Ylgj6PYInQH9C0crMaIPTYXq8gkd9pcJbuTc1hY30OIvWJxj+buv2PSQAH8VUBv2W1Q
/lHy6Z5n0zTq2P4arC9NLvBbQbjOf0ujyNVw4ySfJEkw6u/szcBhS8PVLOMvh/K6NO5f73veDVCk
9zKHto5fvpaoEENM5Sglzivt8fYVBIiQBRfFNjBUCG8Tl44nh+gClER1c3GGnkga0TIjxJFyio4u
gyqeqoNqhKOBkUXIAfjfZa73rVXwtohDDM0vjUYJ4bgPc/SKk0XAABKpQjPik8cUaUI8bEIn4K24
Qj4oKC5/oXbKRGPpVim9esm9MRZMbu+O9AecmasTc0Sjk+coZXpbNhrreFy3bKdufatBnHmXpfpU
x/M6e7mzuZ+6QI3O1bGxIFPxAklaFEcwoz/bQb2UWVqQ9OugyA8uUKl7btWnfrf/F8fpAo8qZfGj
TAliZN3wNKalGNNIS0XpacCxAWbIy4fh/5MV2ucL3ZMg1eooWM/TPvfRdYr2+mqHyqqFqZbHwRnU
4xUYTubxJBuePBsZu8aftnVz98X1uVYZa2AF6KmjSRbCNww9rMWVx+9q6oOWmw3hLBDPFFIQQpH7
tocK88rewvVnTQafqylG2l59UHPPM7d5aPXEKYNjuu+Glw5tJ1j3LEGqxlXYO1hbqoBjOVGOpa3f
02eiwyldUXb8RR2WuL7U7IU2lrCSKLlcBu1kX8ockzJqfC7RyrpMO1+U+agUiDwVxscmDeASKwfT
dUTPBe1OTqJFTTHmCLvG4Lblu4hyoxVTny9O7lAxeee89d2IOQucehcMgzYWXRlqh3fxCMt+kPPP
DutIf9ZOUJbyEezQWQgyOsM47c/VN47efvdhYxMuciMJeSknsqpz+o4Hn1vNghP79AjxGrJhXpT6
u2ZcZw4cDxmnoPqA9+16sEDOxkqgSs209MqwFXUkWcqflYtdK5+tgB1iIdA3YaQdCLDXmLyxyzGN
29LSu3I0bVRSfzrbXZwgd1IeV7C6Uh2J6hi1RW/HCv2Znl5FIxrl2z/K9UPiDBSmTssQ9wZx3P1S
yizkUpFcm7rRUiz+4prLSU4vGA4/UPwE4kbGQc4Fw7X4dWmwcWCR1AH//c+GLUJ6j06VT2gUEWY/
WVqsVo22C+elIzDCBgbeRjr0V+de5qL5izGhjjFi5Aqk64YO/c1mU6UiIfWnU+ttDJ5Bkj0ftlf0
JNOOLX06SXwRvrInwubPJ8uQvH+4b7m6ZIDEE6IZTCOJ15xT/6RUp1PBiF4xd5mVtGghQvgExesS
rK60+6F+t3nYJnfZqsK53NKSegHD9LLzTowGrq/f7Fd2YAaMVg+OECbhptnVTIArDKYdOhskMcpN
yfeUnHrHwjfO+vnwxpNsKUk52gbtS7Apg25XZupimZNZsG6ooFi95G/NVuSqdlDEssOV5eLsRyzH
wGBXNtFoozaj6rfCUVSKzhAlzhDsWPqwQnCBKhOiee08i0fGnkWNfJgbbMSJPZAgwpiXoFJT+GDM
Th4bq8Rw45izEzUJr+6jjuKA8khnvgVwJyseYLkOoOdmgu5rYKYPYLxZxChLyUBp7O0BEoXDPfg8
2GPPCEF76Gzsxe9Ai9n9sG5E/NKK+jKDO5m7RpNs49/Ruu196NwzH3gLJnxC37UtS/sBntm4Q7Z6
ORpm6DSc1vRo8zgmgRtpzx7H7K21KEZxgyKrj7PoJTctFxZhDcKNgUGsY+w18Zy3scITDgDpgYvl
fIlEHFtMfL1pWpxw4hem78RptGKbp9EKOVl212bZh/SqEHpCkXcYZm6Nqms5bGAZ916cUu6mm51j
odJRlBXkbSRgCjYWfSVIE7a4BUMD87JUEA2IksznZYVxXLgSkHe46z25PUt5e8auLJeZ1oBpjUX1
J6yNtqMn9ZznOcLsKkxiJbqb7EwYxu7KxaSlVyIetYMY1SziMxD9S8Sp2dwSTurMLhmxXImP87Os
Iy1TbwXIY4zwRr67esRdTtbOo1El2IL81BIi9Tu8tD02HCE+VELj/tYcT5rLomIQQxqa9gSFxPVN
JInlrIJvtMYjDsd9YrRtW5awN7vE3aFbNGyjDZI5MV/xIhu2+G7xSekirssnBFzAybgYCuvdcCp0
+JejtL7sT3E3Bd5EjYrQ3zmfkkyXKB3p+NcWmq2HSniS3KYs4EZsyOXIO6ZFhi2m9zZx4tBygaEO
TYO8papSrmPBP/A/+mRXGe9Z1mFl/Lhi35+G1YD9Ug0Fetn3cHfqpG25bbLTp7LC6hAvPXxuiiiQ
OwEbzAe5uoQgYmcJb//UuUus9zE8b/rOM8RBHWDzZ1ouvrHHp+CS0KaQsDK+q2IuztvHCKA7iWs6
0Ew1oszs+xrTsT9uZxBvVjYbfeLjMb307BukeQSKf7guo4MNL1cQ3YIFz9wl/b1HubgaeiM/fxda
vLtq0VDqO9ErnvC93UEnYfH5GHuBQ5kvRvAL6Mx5otcj2VVe0icE1yolzUvwt2WERBHYMV0k74Ss
Jtj315d/AeJXlIMGF/gW5w/NCVS9rgAKpGDRT03R8Sa6Dn/oXUQwShA4vPGIsC3O+15sCIKOPWPZ
+sAbTCEquXvoQVwAvc3X8kPbDaOx9ffitIBPr7R/nmEP3ts51r4SXd9JzO5XLzJYh0ue6k5qVMbF
ZlttlB/O/BkNZiVSaI8jiNPJQz7RfHB/Z1L9h3KnPmd3Pp1JhDuM9O1fvYQUZrAEZd0F7ZZBIpDI
TgOlwU7rueOmoQ3UuPWyqhcknpmMAXBObtTd2We0tA65JRVfmCLXuSgcGXa1081KwFGc0DTJBYPs
FEoefe+4c3AR+IUDuVb13CT96XEVTLNSXUuy3k27KvOOioNkUy8HObx2tGBqNPq+JPqd4EzBklW8
bnOB/lmTnJ+x/acfQQh6nrt5nr9P4/F9XuRWQXm9O7gkoYYAoZgU1V5M2+XgJr9dbchZZxr5V6rD
mypOrDCdWD3MFdxA8+9aUBK390c/GArLjqkJEZU6hx0lIrq7qbGAmaImJNVSd7EDt8bOBvrQ6hoh
uG8flgjjFG61pkGD8mAXaaxUaizec9/OCtGtduu58q+W3Ud38NMLGZiWGMynhpl75Q+5w5oSuf/3
idx1prsJyfXNpL8JNS2GGJ14SbkenhB1IL8m3Y3P4bPYZzWiTz7Au2Ne7ApgzvU/76gA+iPTl088
IlVWlqXtbMDcdJv9w61JoChEK8wQxd4OSdQiT6HiPSBiUe94D7KjSmeuGD8XefDV4NPjDmAH3tKF
M85xFWoy5Nwu3PVG7leOHK5LSjkg2TR7yguXxs5R8hzIsXkhIVoTMqww+LBBbxfbpVEbfCiVP1Rf
iAj7BPykxX/Oevdlo5RGjrj6Cg5/a/1tDcE8bK0gFBtQeMtX4uInjsspdGgPY9I0Bvqfn0tsKW8i
P50W4F5bu/clvBxr6/K8bSYF6MaGdsLcrp5soEBTCcR5stxogbYsROW/005qjAZkxSttQzPrWdDP
Smmln8Ni+pNNrGT6SC5OCCndGvm4P6hTqS9VCFHl/XAvrc+NW2DT09CdVkOUpl7uIKnjnBIzaG2d
KlAWSMfdNFGElC1WdEtorwSj/OCfPBuEsk6SsI1LU0h9A/tFv7jsB2KE36e3JdetZu07q9KAMqPg
KUmfiUq3QrdDAFKpBTVtqezzJC6A8PPLgWZHa4BTpWM4Zw4GccQ/+gZl8A+BQ4nOYAcVFGnqBiPE
bG5KIzKE9iulI7nhe3KEbhwPW/TfF2LVxjtTezArt85ne5GilfRd5GhzoyH6FfbgJKnuHVZO1RcV
bifkTjEh2OhX1eVykzbPQ/Zc4wzzlXJDs/I05ASe7v5Sj3kOUs1acG3sSAMNv087JuYs/cwvm8rW
9egcwprFTySwMyJc/idyd5Df+BcYg7sI3YMvl7rc72Vf+CWFnyj0hz7JYsxOvTTm+unBA8t67Ec8
cYzJt/IINmvt17rlmmeQHVHU+F6KvzbKM8nFMtYR/DEw2Cat0/08hGRiPb+qxlI4aUdZWr9d7D/H
0slLEikmDlXYSksTtsks6GBaomkEyqVT9enk0tJhPsP45D0VgLcgsiE9+dciqGFI1EV8UZv2SqOM
EOtJEzq2Lu93Dz/Z9lbnqPN1VL3Z2lrKAlxtYRfMaBILibusST7+MzF4REjjvy5H9n9OXT5alUcD
rP4fCoY2x/r3P2cFanxsfnNC1a4TCq4jeTlOX4adYUjmLBLaYUjMEYUNXqu/sbqZRIruK7pUO8F3
dYrbxkw77QH8iJzSRt+WrvrPoGypgPbGmlwhGUG71D1oiMHRTOaJ1FdamM7o5AF9iAZNa7TO0VLx
vvzLx213O/SmHycEKNPSEnBYZw4srJQv3jYSrZZIt5P0T6CxsLkKRzqL8qUAmYaXlCrMia/1ISWr
xzo3HkZzji8OyQTpURuv5pdKWOt9ef+XIH7FnQjxGMyvz5hsKFflOlUbliKu8Y/+oGqrRq328QVr
xUJH2nMEqN+4JTeDBjYapn441ylZ/V24oSVRchK8HC55xjw4r1b4qS/GBrTHIHPNrOqO7RVL8A0S
KDtSVZP9V/flLR3Fyz3BLMxRlUQ0J8vfh3sExjLg/BDYt8w8HlbV2j/MEuaxIeY8vKGpVWCeSmhD
IJXtPh4gHaudK5c/SDo+ESFd0J1fO61lya90jyjA5ZLk8eca5N/f9cPqtFobVIWWvQIXyc1WRZum
Fqnpa6GpsiOinkkU7iRvuFj2Z2/qBtWBvdd/VV/fh1Bz7u6tyj8p8wO/iui3VueyLQ9g4RTPT0Fz
QIQ3vVYwc/fksuRthDIcOLXWBqNsgtc3MBIdPCHPkIySyV/ady2Gcr6MOxzi94CFXSIIwczNmEnq
XEs2G7GCAdQgclP0fBbTkQQbgPokFXihivUIHwUM4lTG7af2aaL7IdITSChiCLMzbKZ0JJAim50G
Tt6vgbSzTu5f8Dmn1U9GjGspOxl1gkKlGVDepqtFSme7RTeRcqBcbozHNeRtSYqty+ojK5SnbBD+
vEv0GspuB8GGN7mQRyvFjiT/O+dQZ0pf1QKW+2vWiol/vjpd7uOm7/wjzGxUj171bsuZGIKdWRXS
3MDg7HElYQI1FgfIZAEeuaSCdZRsspChsTnPrNSgbsemldztF4QfDJ6CsKVNORpBg7H1Ef5Y8arR
TD6dX0G4/W5RNfWbYi626Au26i1kmySzMw/oWydm5Ig6rFRGl8TWulOM2ly3FrIH6jA0U0X1lAo6
kg7Ec58gt2FC8Mb8wMveR9AlGRdm95XcNOPcOICDU4d3FWyNris3l86c9fO7sb6spkXn/bvSznkN
6uL92xVk2IplOfubkxoAGtNlQhH79tSnFDucI8lF8smY0j7JWYLiSHgCdAJ5Zn5CrmzYfZWIAHxI
cf9i7r8X7t94Czg1lVsfmj6gSPbzBYfXnyrLzlrUnupJDwtnvQS4B4NqmYtOufZ75rzroHcQihni
+7/jN7iOKQ6OyQZwPMsimHD69QdhN7L8fAVENeu0HHsGAuIlZ+8ttGqcnDmi2CwoiDMj+36+Xqd/
RArrsJNq7+Zc5F5x40NH+iXFJQwmSIJqQTnrpD76Im/Tr8LGqo2roJ0g+NvC5NiJpP1zVUf5nxeY
SqNhRPkeVpNUbgelgE/vz4tguL+ON4B2X51eMVP5qUeD3KlHZLcKKH2KnBOfkUFuN4iHN4PXiZab
xDXqrgVyIyM0H/d67ryzmcgSn1Tb+AmRQl/HXope2pAfvl3rgpj3EaMuR+UPn0GCuBCe+WcUPtal
Dy2SftbUeFu+Z6KuylkoyK7IX5NysZDFGHPWqWwW+Wquh1BpymTPvEsT0ZVPycJe3g2LgHzQkQGn
eaK23XHTwU9UH//1bWVcUqGxYe5NuCVD+S7xqPJ4RfYb8Ossi7gm4bGaqQJbtbX7TVA7FBiZJCjO
y9RqdHv97yC8zCFwgCzsXjDUCXrzwzU3qVHODx/goGrLLdMZEU48dKYZyiI1+aU8md0aksbOQcxG
4rhG1c5gBG9Ss446tTgiSbLttWh5dDBDlV7TSeNGgbi2wIGcy+kHYIwD9aQABNwh8im7ZI2VL3NN
ol0Q85a8IpzNxaMWp+BONut5BKyu0NNnWPDLsQlWPNMILRjKa5k4gf+gvCRYvaVxUQD/xMvsnJW3
/PgrU2xetXztTyPW7Oirk4sTfMDY7mqLFUEvAvQdl5Fk0fTtzXBcXKwZByQRBEZFYOViIqGvk+4Z
N+fxMd8qliHdh3I0pa86JU470S1kNIRcubTUjI1X9f1fWoZ0Z7hNL89oSDp70/8ZNR3hHOqHttOC
ny3BNHhfectsKktf4uUuNOTYSJRq87caLbpxybUi56MZUd+XswZZ8mbHrUIaU+iPHJSTH4sa/+1B
AM8zoWYicdCo5EDguTe7FtnOPFgBOxNgeQvVsFeSyVHxXHD49tiUUQ7uAs4Zmn0UcO25VM553+E8
RURYPTRlIz363XoJVXssQXq4AIHJ/FSqpmg50eqLCdKYx3b45/wYWhlAEg+N+h217c7F+mCc+VCY
qwYWSYJ6YeVvOzsVekqlV2mPwl+d6rs0V5kEG4yIJZFy1f2vPyYaHf4r6bOAux5ADLnFL2eet3Fu
Uh6AgptBSbpgDn/M0pZbJIO3uNqnG0wAAqSx1Ye1BIJ4khYLx1hGGURXOtwlIb5SvxIBiPZY6dsH
BqKLLi64dAtYji1wCBYSQvXiUvn4yrtn/wS1kwsmLRirgAYcfFAJEQC4P6ikiRXner+LFUxnPJMj
mSuwWhgjfV/uDWjJAQJxoerz1MhyyNDr/dzKPlKF650DqgEDhYWL22GhtFkdOtfbhbnK+3FUYvx/
AKPtKNrR8NC1WdpDGXHnzIPUSUQ9X1jNAHAqq4h0JWjcICXqpdOXoak/4N/xEnFStFOvmdt1KyU6
kv7zKJzFcjpQwY0y4UChZDnBKB2EhuNVy3vGD28SR1C8XGP4x4069+tU5hNmhjA3ih9bjoqaT6Ih
wuLwSXBs4UYcJ6yanGc3yWVQOZ8XqrkVJ33t4H0fZu4tDiwWijkJovEWYMcJdrsrTqnNp8wm232b
BdRh9KqctSPd2/SPJrYbu3oJTG8vSdesguELmqJwjwqBVjguEpM0+dFB/wDxNOll/bigQaPQI6du
dqJV0srX8T6lkqTTq2RiFtEhasNoxZ8pVNFfp6iXnqwPRaFrKwW9UpAayZIkszsllu5X+IWD5gBB
vcicpdvXL5h4Ht8K+muhPAbbHEIF2x2mnNj2Gsp0T+yYl0o+Ln5NnR15yVuo9hfqi7fTigAaNhm/
ZAJpuCQ5kETBjJwhCosm6F9b0JgQmuKHgKjf+523ANM6pvGRDm52FwrEatgOAfwquUAojJQvGjh0
IXoCP80OqmJpbRnqB5eQIckg+mrtVZLRigPXnInGeuN84RfVgNjvpj6XCQ4xtJLtOqphpwv+aHcr
Nyvgno7P4LUM5RXeOfUAr1EnbCRm66GIW0t/OmHRLN3hWAavQl8bmhVxWGtAXdmV8oVoxi4UYApf
QxtWFIYWk0CFvuA6LY1KnjvcfQGaQRwjjIhsqzfmZwmI+QrstvJ9CdFPGK4htHTTB9OVscDg80mG
D+crnmKjQYlFHyaXXuDY1ZuG94yCVEmiW40hkXkO+x945vv2FvJGcP7vn+xy3QiAuYB4FWev7PP0
Ji35gUCfXrT+BDguRmpIjpkvT3DmrQRd1PKcM2Ai82nkXU3fLl3ztYrM2J92Sm/bMqESaK+pXkW1
Lkq8AuANxm2Kh7n1NKkPXorw1vbBUGVz8dLOyl87sdwRnXgqwn9NIXHcBWaOe3IgLoBefz66N4Ij
fjkyIm64Gr5k7hToPJWZK4HrwpWnT3zAtCsJKtOSe6YiKhfXC9N/0fRdplhOdPaxd1VnTKlCKdQb
KyQFUjeFiII+itQ2UFWBtafQN72JegOX29MoHqIgIIdsjZnpactTIamo0qDdgGnzswy0hyVflwtk
AdnMrtVbX974D35hZtSuWWL0I0acFX4SUwmPaJceIhgvE+wVIyw4SY0HOT1Bmsu0t0nh2VcSR8aK
NuL+RodSbQeaFf9aT1ebpvIx5H9TekX3Ikw7FqUYe+Hv0VkgmFcLN4Wz13VVvuQfXBFxNjw7mF+H
NYMdA3TozQODdjQb4vSyn2uWpmp+b5JW2/TQdSyvWyC02ViwKL2xiwaQmeNR8b8RxnNvsL5DSxWV
zUPV/NtfE1vja1lMt4JDKBDbJacE5qsOdv92QEuyBUQMAbDdle1uBXc2sOzTNDw91nSMlISNtPHo
BLJJKiFC0yFtbBN3wAjuRjz1XQdTaYoG27kBXcqrMkng/FALd63OGc1E24KnsYM3mjk0xdc7XUFC
5ykn/dT9HKbZZKLkvZqPpTQfTq1q5hpCheFCJ9RTxTHuzToH7muTv6Vfypm1VuJgNPBSI7liNp5Z
gQUJr39ezdwcf3cbxlGDRNC1lVuC1elSjL2Ss4zr6cnuRxWvTr76F3p+Gj6B4pFQTFEhEz6BsYp+
qdoycW5Q6xWkhElNrkLKAagYxunw1N+pRc17ranrexAAvYDC00281cKdwB1I2vUtP/Y5TQkzRAbu
lvKEeS45potkO/ZIzXeKxFVi2eTfW3X6Rv9MrSsCpeR6DcuGjFjIA3VAptFDlhdvDerfhLEeZ4dr
pkrf0sn1dmcOoNMoVqHYzLrVRq0Xw+YNxYBIe1lZTVaIkQJsfctT3tgToGx0O/GDzmCplQ5OMSfY
SYKT6BIACZsKTHm9Q9na2GY6Zlg5wdaV2iC/EF/P1ywlqHd8nc+WXNABKDKFLH3sdQO3LLYIYIUz
4pjJR0RHuCcLrNLQairDuy/G2gqePa/Pl9rakQ99cFQ+NdKJ/7s6CBB6ps7Vx4No7mfd2rScb2Py
Z9HWrAmva4UC5V8hAOVlZTg5u6zMzNAfwuql5VcQVi/1eMLgkYeSA3onhwogtCyaIUfhcDMTNozM
a5A7PRmh8f5pLeAloaVhOdW5Z3mRyyt6xw+2gt5/2VK27ANwHtOoPS080Ti+dyQrTKsJHEk5SHl+
CR83l7BrCBgGfZJf3O3p6cGRjcB/7vo4cpqf/x8o17u/Z2jheXHBmD1oOZf58Rrf4CJpIqydTY9j
x5zp9iVVamp3Vi3/y8CZI8lMiif2fBcwh/gWFTJF709+Lbm2MHakFwryQJj94OyOFOTzHfEn+haI
ZsJw6FJPjui3qlQLDbjFttxHgeGa/mFuWgnJjM3T5rCEarIDbn2UhoEJ9X5GJ4cye4w8uQDpy7tf
wNeA+703ve7VLNTEcsJpw7lQsvuzqbkaLTAFgNB4nEFQ1ephZ2ZInxdN3IXshcHd27Iof0+w+sFA
BzJv1+we7kEm0Z6r/CB4HDviZO5bFPUxx6vG1KFwmuzfg/aWVUf0lvav3jdZWTzL262XgX/yBxtA
efcvx3uquXv7g5Lz47togwrEdkA72PTyGydw2IgzctVn0SZl3mGv4P0anM2wdIc5jU8FJF8zWUHu
qoEo+H9zPTAjIRnRmLeFB2mnHDLG8wNYCShHNjRpcXcCZcAnt4lvJgy6HJ3p5sm19F/zH4qkNIc5
0nJzhgUduTuM1rAfLB8VmQzH+eN4Fg4awyzdfxMvPw3ZWW8HfPvUijJVcWkt8r8WX/zPAWD0w1Fz
woifs39yS9m9H5Ha1TDU7wYBrZDb12hp4e+VGhTJwF0PzZ3CUmm5QGCDU+QS7VFQr678mlu/vpVV
fDElAxsSrP4UeLVi2U7EtVbnazdemsoMhbqwlM0I6vnv2ErFDDuYrRm3LTsj7ZPPKWMgyNUQwDud
lmnomMROZ2LAvvGahir1+P51c5f7bV34RSAOsy4ZPpyNaCZdlabXBmhbXf9DsIM/krxGxFZISB61
9gW4EpQkk88rm71AdVQmsyWi8woQZrpnmQniDZGMpUwQ40GNYEQa72KZf4f3LxTipYtwdVT3EMG8
kIpb2IXA+OoSzALuO4tuTbRVpG4mHjGrw2vPxx0Go1Qt750VZK3g9qgXedQbvItvL6Jhtglo+ngh
IEKXu+IAJH4bGbqarFf+1EpZpeNDmlmpfFXC48BcDUXjuQrdfnCbZgURrQ4uBW9xgBcbxJGdFzuE
ucWoTZ6L/IFos2eewvkQQJL/Pr+5GmoGAuJEbwRR06RSzm0DNwOzI4/7Zc+0L0K82suVKaQ/pSbs
QNeZVWaLnjMDL0qc6aab5mhSB6Iw9Y2P4uyJtYJCoPvd4WRuxvbeXDtYVuPoS/pYDNLZf8lb7Bam
+nLSdrrmedTkwiwwsYr7AVrdBeWMLS8reHS1juHHtV7zXHHARsDeRMSiRL8j5DyBaypG3SOJ6KJv
0SCC9WEbM7sIxXbBRAHogqZhPe+p3tVdZqttWfxe3adscw0I2kzOFyWPcTuPH7OenvISAJbkxsw2
dnxcbsJQ60xgrO75w6xFAwpMiNKlNVB/AlJstkCCoLvjwZqVaWnu8deLOal8SgFlRNqCY+es5uAY
BohZ8civunpDAm7hRn1A/Uxj2eiovzbAHPX+gtOdtBpTbpW9oKJ1IPYyg5sJXx0eyDsqYrMjtvb1
8wPqeR28We1YxaGsmpRvtzn9An2M9D6d5jwfc32EgDXLJcv5SwmTs6547+f7V9igLTyEVty1pu56
+PKx6gkfPIUE6sYZPjR640NfMqJYZg3ag0EzPvtDkKhUhzI+VlfLAGgxw8K+uBSgduflOf1avoZB
vTUE/CLCNNIcPZWOEasiCO9u0SEZxj7SbKpEDInnFLrOBoAywsFrXSSSwSMZriKiGenmLXQqcnaa
4fGjH0kVZrHuSKcx4p7rOlHUbYJKsZRLTJ4XOkT3RkiSsuz3gl43OTcIedm/iRdleggT7a3OPQqz
1KssMo/ynEQDbXGUN62DkP6js/Owmco0XcE1SN2bVReqwwUFuFp3c0qafKQYcQ4ynx9/f1VczwA0
wxAhMmOh1LltegL0hIEp3A4ewGnbGe82ScIdQF9SNrw+IESUK4FYxs0S4DCra7ns78AeGtc9FZlh
BPxu8G1cGS65gJgwXkWu7fdg3TkeVqVH2p57Yd5kuXX3zR+aL2PL4BlYUgk1eMs01SZPm7mU7e4u
4lk8enbjRktbMCKGEhAArrixPoBxeZzHiJE7HtvVIPHlBCLma4t5bPysqsW6Re+iJEtP5t0KgPX1
XVUTHyORVAaRmV2tfg1vWsWL5XvfsinaArONHsyhsnzzo/2Iy9Fj6rr3XD4IOWyOrxVS12/Fsdwa
n6iZlbDN7QVdHD9UFFMMSId6Ri3MT36v1vJvkpo485r46ffDQqwYVHBdkiWFBGr1WPzqaETVqTeq
cN0Iimc+8d13Hd8jPrXDK4cchncevaQw3Fg27orVPwwl6qtRpDJykYhyKN8pEkXCp3uWHOW+nR9e
wBOMhv1fnRhzrM6dsiw0aRQsBYj3xYnu7cIr0P0mftH52kfnXtcMzsdGSmZzTezBVPQTDPu80yZL
usTSWMq/7l7HwJCzMQK918w7mD13gL2ZNivb5A7DGZCvtZBV0PZ0tUaJer3wfuKJlNEnxPcO5bao
Zf04F9aab9Mg3w39z8fxGXoO6DtZqU67UxO4PrYxL74z6d4hyefnZ617K4AwpwxbVlN4ndZJvvKI
uPUainJjrJiiqSGn9ZQjSEIHwNwQrlOO3IcBSrykHk4EIQ9KHtKgTbSEUT9mrWiU26x2yd25VVj6
jAJeAFjXZxrWXTUpYy3G00r5niOmM2L7a4A0XPcYCLwTzK8zJY3rTjPFXISq+6RYhvSOAaaJfggG
vNoBVaXpdUMm5GeZQ1cdHVAvA6XBzlLwlPn6eErEV+KB83ltHIiAq4t2gEJ5T0Sjs6K2kicD1pA+
aheQNcBryNJX+IcTn/ybaKArQn2fY3uhhMtivZJK4OrlaJq5pTaZ0F6ZFEpvc5N4T14jjz7zAl2H
RR26YWJTx7oWVajBDq6nQ+rjVgojWBkATxSVgMZVgZ1/hdMcdRZAiPfZM2HxwstrUXPsYqOmNww/
9TlOjvM3JkqnadIgUyniB+gQXri3o2evzo7rvFK/bRAZamWEOmivRfcJh6hpy22YuB0AWB+vyQHj
RS5y6Z8I9ug0QAli0jL8Xjx7LpC+/KDxVUGzUpYVGGOyuXn3Q5osUNN+Bsbh2oblPjGBJ4JWOYxu
eGxExxb+7vmcNCNcLabHVc+RxBqusUwXlUPcyo6dIVB+uVUmaefrF1Lo623d7twf5OUW0dw2Fldk
rlC5OG//Zwi3YlVhz7sxt9DNTdhB9jQoXesm8Q71eGxWMx/4fpWcdbItcTvWrZuegp0mR52VujSi
afydIh3D37X9fsB3lOrl0GHkcfc5O6DiOpc1ae4XS7b16KD1z/BXm3vJ52XrQxPkALbmbdTzZpSK
zoiUQTvaQUOQbbG017zzwP7pzshTSWO0UxV5PH/ksncSvqVYr09HMPAVrJqVyhGwcPZ6MXiWtNT9
T5uHGROryeORiDxQkkIQPoAK5rFXHldFNX01+aaHcuL2lGTwoyn0/iMvL4tNxWTirmYaOyp3S/vv
cwvf1yrMGopbMAo43pI3FqlqtOIPFKhpSDVvAkpbBEFGQLesvBtzr0QbxKJDCcSmuq3+CTkeHLPI
hlL6PTAqMiMnOM4+iRF7XfyCFhugMGMfS5kmpOzBunmfIMot71g2wzPoCnln1PjSkb4aq+U6qxKz
fG+a5RgkbxnuutSedd8Rv1MuiIv695lH6j4hV+0rHFsjGC8sjvodAsJ0XeWPHlQrLnUaOGoE20ZK
APbalWU+WFnH4LSj1X+mpvfU9itEXBqLfWweglv539BzxiNYn8g2j8ZiInD1FYwCOtmR/L/2u+9U
bw8KmYLYQLu3ucv3DuS12AjZOJtOSt2GRII1Ap8mO23+FIzIcemYy6GrToQn0tp16dmbFQKrNR3P
DgqqjMQ8Nz8TWJgrQg8S9HopaqGiXdvxxinjVERwQ4mqNl2a38pFjrGf0Nd8yYPqWG5yBxZbIw8u
D+CGJwPSOwok9moCrX2PCj6mm8BoKrr3KP15kHClizhFRhFaFLcyFfXV4yZgbvGtwwPDusViEJ7y
GHb7IZEQMGMBxai/O1ug87nze12a5DsoIKzLvwayu6x7E0B67lhfhW7DaJk2MIyrKRS1jC3yXV8g
ToLksV9O7Fa4fWkhWx0nw+aILVEzg6Fz66eEC9MawceuhAa4sJfvSqunXs1PxPxi/UvLfL2NUsnZ
p56z4X6I0lAWwJoJF4ztoo3OPmcmzUKj5pDOyWB1K+s2u7SsIDhJg33InTtKGEfiKFToAluQ0cFw
rLr3s7ksz1Ms+lmbg8qD5JTAPDvlZ+6ACpFthZNEB2zF7GkaYBgjnis2HOctA5ydl+EUZM1GYyGS
g4ErhUP53/h9jAkQIuBdBScWnsA+vig4OY6aVgICDNFvd/9NW+VGwTqG/7aoAdkpx9ZKS+RvUQhh
bxm/wQj7XK1q+uEVUVlEtcluz9hfOFZEObVJ9T7Ep8c1Us0H2Xca7O+RPSaCb0iTVi7G3ttlq01x
RXGbttiGIMn8/AFYDJCC40kbaKRY+8fvWd+4OYbQUt71loMnXZ14C2/WF9py1m2VECga5LLrOcjX
4bRzkzi/kNnWBUIBF0BWUIhwBDLw2tSC7FOLua4Ltegol5YSoPT4EdtbB0t798kUkulyPklRV8Z0
shAkmGRz+/ufV3aujkCscAg9tWB6A/WBrm35lE02QHg7ETGQ1WYoupbS84RtIreZCjezH3ZxJnl2
MjSmfalcYgybUJP1mz9cDyHeSGbAd3pVorg53KDxoRmH0XJKj1h1L/FtHSUPFtBva8py8ZxWlGT6
reDYato6WHKuPywqjoXXFc8VjPEqb8P0wDX6TjlHACEpxyHKv2HQ1UTlvlMhmyO83F50KrJKc+CL
aIVy+n30PkZLhsIj0LZOIH8OTJrNTsfutBcplNG88naflyGWFbnYVEyC7sskSlFMawFC12LYputA
GRvv0bs8tlzS994704gtN6MofbYUoUKA8FS6kgA6qzbmL5vL1raoD+tSAUjaetIDM7W0Xx2yZesV
5Sb9S9BV1/9HqbQW2QM4yLN6IHSJQO1NHLa6+Va2c0ZA9dC7T2EfkUpq0r9iFmZ65bgOivhuKyHZ
A8iN8yDfKZSJBIpOMrkSHQMBH0F3e8MuzhJdUKNNcwIJoMEJR91e/C28ijWxBsiO0scm4uNbGrJ5
CFAlpA57iGCe/kOqr4oDWLb8+85A7LRJVn8MwHj+spFCWz9YCFzFCmPihIyaV/V9oY+xqfMRuNih
Iul60RVWsld4G+siRQJ7Hx4j5Y1QgcyZNDlqhADMUqt6pdJMQjznJsXE2oK6sbk0ERgtA65lwD78
paiWWEkxOaMHnhn8t+ORvhhJ1tsg8B9T592vfOWvp06IBlTNt88bPsid9vY3OCjeSKx/n59W+Zce
dhpeLCZ667JkOSJzeE0ylxqYX/RmZxFJ8SPF/1TzacP6W98UlPO4ovKX8Z9146D1TSTfgUvOBbyJ
od1qmouEDRyURMFcCit/raDMMC8+sgAAf0eTDiOGkXYNJemov0NpRNsRvvMQ/YLgK70IJ+grLDyt
ZeI1GZV+q/fPiEdsAhKAeDazkJ4f4vkSnXVo4PD9s6olJEQ0LW+HXDdIecdLRn/5203fcgwnf4us
wKeUYEuMY998JtEXLjGi2Nw/4YBc6tXaVbvy6EpSgMYe9Nxvlsh5blCN0RzwC5gWVKpTrTo93Y0m
IR2FTIhNFB4EoLUiYDrurtlK0sc9Ic6PE/eLr1Am+gpTQgVGQlx4pzXjRPkp928M1U4U6EElmFjM
16UPhvcIT4xmSIquA5qf0zf28ffP/9zwmxIIHKJcJ2K0Vz+ouFNv6Bpm1mNFd3DUAGRd70Yt2dhg
GJFpULrgL3CV7DiBQccWyx+YZ6X2CGMYC0ldBciQIt30uZEJYpZAOdKI0F2pJWXUQypMk+iaCqgJ
04SUb2rITgUBW9GzQdcMAM5MgPdlp30QHUlHS+D9h8Aeir5FI2NR/8XFYaLHI+3d54sCtJTkqk6Y
xz8D4KdzGH2k3wTF/PBrN8hponDEcw8fcJxSe5OZ7/lrVaofCIakzKUsQbhxZ2k3DntqXqODO2XV
iCYKQ/NJ7WJJthaEjV9MQWZU2nku7HXihnnkFA6jHD/rolwbQ2jnGjdvHXojpgfZp6hIRYYcKCzw
re7Xwbkslgx+CjE4Q/46MtI+28fC6LBZohitull31+7ta0Gp/IdRRzGA99M5dCZy7ZsSg4bkI8ug
kV9xcpGDcAMf81HZPYNV+Lxe60Df8N2Pcl5kaEw8XQoPyqttG/NxtJx5YT/pRypbrwGTxFEXjFHr
vGE8KLvNKmhcMh4MnwLF6utKRtE+uMHLU5KUb5Ak4jwmTSrdK0k9gKM3noBq4H10BzCF8BOfNAmJ
7EtP57mbthGyDpcaHp06IupHGsvY+osFFcrBAS04JqV3uDwSMlRW+ru/uvQ31BiU2ooBkQojS5/W
43sxjZbF3bAz52+BPWpKVfuJnnYH1Nr6ePTR0rLNJhFbiWgMWv276wzjN7N0EvqPMmBnhrhHiTdj
HcpZhL3mw8CW3KMMWxiOXbs24bvr97jxRAD36MTRFaw5lYhipBMnBQYWZ0INkTNkqk4MJcvdMbcx
9Vorkg0Dxmk/Fb5I03NXC3vkjzjxOPJgzfQ+3FqthrkTqlr8ksoNbcgrNhrTAWaNkD64yik+rNOP
eqdXNFmuHzlAj8W8qbv6zNpuKLCq2HeHGX9tI2w9max4YMhAH7mQ7USS1flEeeyJISYAB4CjtcVq
Ibfc+4vbTg57lmoyC68HUmNtczUveGrx5mAZYFflH9qHnLQlMcbbPXXnfNwuqo2PWFxBzv7Y87v5
XLrpQrzuF2pqret50a3qHO64Btmp5/ExwkoEybFH84xsLUzBmwdyI/YzbehVTVfwM0UXt+gmMMYv
kbQSz40OQI5xqP31aw3IXDFoz9qgbKrf9u99fffhfhqqfHviVPNDpYKCAhhqy2JArqtECSklndvW
bNRhKbEx6UDO/GbvMYD+KyDuFwhTZhsz22j5tb0rjgC5NWmbCPDt3rFPnaBLcDMccg8SNu3SKqWD
sabW0gR6wXlR/aSMJnomg/AdpRChPILVgJyjvrRb/GhjNngnd2TrgiG43V9SdsWOQO2FZEWDcYR2
rAZADuE1ykBrOCLYQ1JvYj8My0BKBn8qhFQx/CiHVJgA92EDx0LQS8MxKWejyIqesd8Kge2qypL3
393Wg/YLIQ2SZZwc49S525Bb166ltlLsgoziWlBwshAhZ/GyXfSfp5csBr2Dw6DSyteI6oRjCudR
wa1mJDNYTgjiSbhuyAi9IgVZqHN71vTQ6XQ2Lelhws2+AKWB/GXBOGBMNIrkhqp9RTKgAoAbrEs3
8g2b+2YYbKNRAHYg8IZD0TwlAj+ho2Gu2Z3nW6ffBkWJw98TD9hI3a47MwtHD7zknOfionWByoOb
bPKCGxz3X4Wym/pWhqL4/xwMaD29piB6FDIAA0RBD5RuczbUeTLeTfzAJVJ6ODG99e+gTCbvLkzo
Xg0irqDs6nD8eoB0WYSYwI27LnopkdTvqwqTLYxeR8bD9kREWhiNlbEMScdY+ls7uvDpvV7fZYrr
Dxx8kX6YnsVP12DO4IIZQoZx9JMBuWYXQ3ccR7EUt7KOvAErZVesyPw9VFxd6FWjmzQMAngIJvvn
+vXufZ8f9oDnFy1tHI30z/TL7y2Pxi+01vrEQjbLMTpqea1o9XNjJFFa+Re1lPJ0XrdvPen2kilk
/BQuNW+m/EcXpWhIIoxDfsttz0C9De/mT1g/ENEhTadQSuVjoio6LDC39kvwrhCvQ7MISV1ySfEl
sWb3y6EJCqYINgdYDnZvaTdRMnXzRjd5L/WdDE7TFCR6BlyRKGkbEjRsWtMVPg7IjsANk8bD5D8f
XcP9fFXebFmMDvaoXqnDQ4DicDVmq0nYdLQLfABCjEJtU1cWrzxtkZP6GWZanHUKIDqgVzDABj2b
9/DK2YadxKzr9UwG6daECIYQ0e6gEUx+dM50pBQjDRRMsYk66ReFxtl3i1YU1Dej+BjNzFOLogzr
vYa56aUOC5DmaP7pUUI7tjg9F8eY1jtgWqd2KWSjQMx+lLuZ8J2PXZ1TgnN2NJ2hoIRSGhD3VCye
RFzFcMwlpdhugD03PuauVRK+Hgt/rsQxqdOfYgrYjMGwj5b+DvkPkRwAQcaNUdUzehBdnttb7HUC
h2MXJFPTFRkGIR57UiyC/SKC/XQdnGVQ9g1SeYYxdYKjuP5n78yAw86B5p4Krnv832lLb/FnVHrB
C9KoZo14XNGErxgGoSCyJkmeXRf4COPD9ovEE7as4IizxyvMR4dWhABa55r9GqpvH/5GCNEf5gnG
vSidkxaKoE/AVMdr3oB9a6LgwP0JHYzCtjOc4WTuUO4LFNlpPb3baWBGijThN7O6aFXJdJIkSBmO
BCX4x1y1jxGJitok00s0ke0zie2H0I5kc23KPBc96Dei4hnQc6VpiiqD61Jhgy+ZrncXffdjSJnX
Jms5qoitRLXJBtXf5cWCyvgGkemT/7fhpvwOSinSuPIdmw4btlYNVVY/2jdJ9LnZR9nQfGtOtLip
YbbonYt2OBGJyrgYSdEd83PbKHYwa+p+ODLGMdkykSQQz2sbz+VqkVNnmPHE1luUFOqWwY+cpBhL
tht2P/fTx1H2WxWlJXJPJ0VV05y6H59xMIzRjuDunJnBwdMAHxPpdIvC5kC9qemaB6oJsc7m3GBo
8VtYlro/yOi94Jl4C6mL0c+Oqa2rXkv5coU09swg3qq9eZomh/QWWSr549SoKXHS68TscgL4eRYg
F2KtlxuUe14eEP53UGs7IU6oTANn+nMSiI0ZH2wTnKkzEDztjNTEcsHq+sqmF0LkDz0F4mRo0ex2
rdbqXichVQAEhHHDdoZt9jj9pqvHV2qn+LmV4+xjrEgRWGg9VDinDCSDnJV0Hqw/f/5BSyJGmUiS
/h3amZB3bqgM+99qveXITAeN6ELeNlQVgpjvk7XQCjeCJ7Pa67QsMu/IDQsDTrT+qTlTvmaZ3HId
SeRFN2v8ZqJ+Nm5wD6Gfq2FkXz2/yrO+Yqunq7FrPehadZSk30XhvprjDNYMMF14oTDVBRhSpB7r
GoMRQagdzKh/o+anrHqgI4U83+7bgN5LBVKGDFsBDMDZQkZMwPZPL4K1p9WDG+0F1wFgCbcExEXm
lyc/+jrUgF6OLl98gzLQ3Ea5AnRf9+XP97f/w3a+DixjqO/pDyjZoJD1sg+pSYYAq2T3eUCALAp4
gFOziWoFE1F0mxIeyB6A1sGoAryphEkmvyyjVEcr1a/X+/eMPzi8q0s2NUG+BcO4zQEerdRoW1PT
Pxy4lc+HMPBLaiZIo38mEu8S4xkKJGHwqxFFrTr4euxMWbyiF+ySmEGNg81aRpYYs6lKbYep6dYb
4/CU0stoL5jD2tMovSJ1VQDZLlFvj5npxb22t5u5pHiqSdn4y+CquTwt4YRJN4l4JED1mU4LcCTU
aLYFwaZQ/nfbZXos6+LEjl2KE6BZLpq6+mUJPESZij73/lqsEmjC70oF16cLJDPv4yUkEbjMx3ay
z39dob6LKDL9SrpIBZKl6OqLWygT3y1Ql1U7MwXPkqSxaIFpFv1Jvb2lsBfFmB+51VKAJeWGX8kH
0QOwPebhsKlWlr3OHmnVdZlWyrrnpAUZ28mT1sAitMFHk4Q5EEeOSF3v59loK4AFrWNZ+yrwf25A
ktK2vSI9CTJoO11eaF8pR7dkF/1TRjx3FDLFSL3Iw3orAS/1I84C9JCoD/szroBXSF93TggAN78c
nK88vibNAB6rVkwag72A8VZLrDIcq0Qs7wrewrYm48NVJ6cNQ8sSyKhi5uxgw5WVvCYnW5MaqMZR
YzcLpyG1ESv8PmfUSuu5VeEc8TlZLSeUlM5Wjjy5eOGSHLwom50VRq+Zf6uBs8MJgVAqkJCgxAEc
5iZfQcYzNd7hbrb0nzUk9Q+swAC3w4kpbj4H/Ky3p5zuxmW10n+C+kbMFR+CaZ0ucm8GKGNpokH7
Qxr1c/t9bG/xhFbSvoBOQp+12Uqeq+f/X3TvBIUGT9DF8gzwpuW18YMf/MChkpb78l0rKWcrszJA
f2TIUOd5nBnMntrwZSXns/bQ72+l+YC8x4tZhY6PTGRZXiYlucpcSDVaQYqsFraMPsK6kFz9o3P8
SFtOZ8zcye76CbAbQUwZKECccKr1tIkK8vUdkmVcVl3+P+0kFpCTL5oWqsudp3r0Y9DoLJcadnaj
JSVbBGDAn1htXoHlP9vd0HM9yR84SMeFMSuPo0/twcnLpLImkHLLXAqx2pe+6ifp500vxpQA5OY1
RzHfsu9hnV99kOmj5Apwd1XHEruy06zsLMN5/nNvWpFBgLaGOqJ0CyosDutOfwZH8JellFMq+1dH
IFns6+4JnJP82eXo/xXUHR+cKnarnKUHzZHRU4c8nIMa+S2GlGT2BfVOFR23nMIc0uwLGQf/5R+j
ps8TK6wCq2lDcQZb9kgYy+XXl63f41m4oEsio0x7xKdIrSBwtkjCyM4pocA+kKnD1+mOJ3lthjg1
EOkDV865jpnwcbEiB9gbFjxDPoi4kKTrhsFcIhUnhdXAYVX+SXge0buX3pooPFzlW+VH1bz8i/s0
KAuXiJ1ZsUV73lCQ/v5GZ1+vW5Cv2EI9YXyZ32oOPQy6Pr2CmIpD1iMeQC01UCsVuZZnbrjIdP15
hEcFxYgRG445Ccjo2oqjr+gM9xoOXLzN6XFf1cid5sKARDdZ40lCWPN6AlXKVn83ANJ5oSWqZZOT
aHvSEG2oAdSiKjaggB17AYsOZ9ZeRobvdc4HtpjBKaRmEX+d6GGSCBklJZgWQyajfc4X34knrmli
khN3h1xurB1qnfbU8VVx8Cj61+IU7nzblWyvEY0IQuwBh4bddnnxVMzFt3mDMm6xXDZSMYc7Cbtj
xS2FFlDZYdfE5qwwrDbGklT3Cvsb9AwG6nPf/hjpKS+FSwzSbQNAjvORLJtX0S+rzHa8YuiuIaZy
eOO/kX2whkqwQ/2qVdErgKrVc6MdlWpPBYmjEXq31+0JsTKqulvS6U30qrgA6GvoHJgryvuhmRqB
ag0ff2TZktecAOypSTKc3ktjrwuBWlI1RVY4bj5IvWeCHJLY82hGu6sdbtNv5NuZpgb7Tb+E0bdg
cLhJooCBjjlWqV7boX6BeyNwVtMpCCCamcpiNfpB1BfKnPaRjqXNkAto4BIHqEoeLZsDz4jt6Yt3
GoquNaCDVbbG3utQ+5+g2kwYinhfmrcn8+bfbULdbSV0FuvtWB5I90L6oDAKWXYtHrwd8JuUZhIH
WtIDTxvGQN41mpA3gaRfnngi0dtgMjRZxeyuybJBS0WKr+Zg1TVxRoOKa7+6zEMnCQIVYM7oUW6b
UOBxZ5Gh7wOd//cBqyPV8Xip8Cq4IyR5X87ElXoyY70uIiDjLPZKfMNde0xbwR1uCab3gB7d/bEO
9u0trpLPbXas8gsfgHEYWEb0147fbQtgqK6neQNZBDzOxWXYrBzhpGz0kAHsvSAbxMrKu+DWhdpy
90qFvgT5WyTrZ8l5aVWneuFVpkUoILymQ23GQmGxwp76j9OUP6TSjQKRyUN9vm1eHMuMkLP41Ntn
7stkgLk6aG8KzA8va1TUNBCjA7VEp2e10BOl+6F9VdkwLJl9YCgs2Zd5iaZ9J3IFWziIdD2mpurd
3Y2S0eRHcNQ0H29Y7KHMCkxnA2JCeUqkD3wkIxJzQwjfGtSFfmU+yO2KHA3wm26jRDwUIiAa2Wf6
1XAXVcN6S1gZpidPJ7dv9AOTLNI/uPD5CcE0dcEXjCMP0IUnIoviHT58QeGwkwwqopgSZelfe5NV
wSigSBt+QvxfIuyD0uyCWBHdkHqdab2JWdqEZW6Tomt0h1JRuDpJ6WSDbqlNh0INTgs1NY+Lguzk
UGm4MOZQVpF9q6vgJ3cfftUqmhn31NA+RtApo7/4ogqY2OTts25kbvUT6xrQNJjt745mOypgYh+h
Fe8WdACduZp2gnZA5g3ZSUm+Ph1Xz+ZZ0Am1biOE9z9IcBsPNBQsz5qxEJ51TDwXQmNdv71TX15l
nM0c6JQkj36qGtjdBqerHktkwzd+Vfyvi4yurdb/DVo3n8hvojz0Chmq3DQjpij39k/z1V1hejF7
zJ4P/uBUFOqMhbKNIecNMNJwFn9wJImPWIMXcH0Bb4/DuLwr8HLeO3GIbNCytPZdJk0yYBH+9EPq
gkDa1nz0srBROAXjCW4Ngmvaf7f8AnAeGYT2CaotXr/oSRr6T/GfvM+Pf7G+29ZYhDTcR6/5RXZx
B58ZHGTbyW6Tc46ilP4xEJ5GEqLDw7ieoMAlOX8RfssjH4EcSSc4z0ZevwTI5UA3y7tDcp48eujX
fKBrf1Urnzq+gTTWzSsOr2qdbB7ETfjQUaRdDXpeV0Px6N4a6e9PqIzLNr2yIWJ9upW3PBdRdyz3
xudAyla3pL0ISQ9KerVoguKsR9bR6PSSghDfWJxutYNeaL5SWGq/J79L9TwMMb+zvHc3iXe7yYf6
RXlCxsWGcWKayYjNLfl0FRaCJAPUso2/zfc2jmNZQdd06rRHABOcgkVS2Eoq7dP0wMAgr93I6ocr
SDL/el4oDIHJ44oTUqXVLuisIsqtokIFLLaKEazolZ5fAk4knXVojeuU2uylzPti2299j1Tg7eqS
pBr8IDHo2rCdJn+ktEt7Nb9bzgArseX280MqpCVAwzPsoMZ7444dWVa4PmjUvNh9+IFxgWOhw9T6
DnienE2GiNWCi41EMIGHVZkWIRWQGDBnMm2bDLpl4ymcYAc6ymxp6bmac1XF5AZOTH0OOdNK98b4
grMPo5IWQWFmz/yX5Duo3kW6KbHDO3301yzUIpI1QbdOwtfBadTCfL9OHREHo6mAC7Cr/tkte6wX
vjGH4afaTC7dptiVHkS6cNkVOvPpAPRCzwISyG+ZFtU93SwiLbJDjwQnBbsXzh8slIXmV8+mndZw
CUxeTlhr0NOT+VbJ3cjiZZRBGob42YA+n0cvBfqDcTfSZqzNlZiCu2Kf6yz0ahzb1ohfviKblsUY
ZZ7sVrtHgP0nOn/9IL420Sx+2ayFqj8K7RQV4+oVMYYufpYrKeS8iiio7hUg/4+MTP5LXAlRHbrv
icL0kQ/oOgckhbAaPRo5NmGs2NXlDL5N2dZfRJfoKLEWMgia+aXzMzpCvboZiivQmz7u5WewCIwX
LhWTAwiUwmBh9MrecY2kF7acjYpE7Mrj1lMIR7CHlv8+sgZuO1Luoi9GE9d+G8peo2QD16H227xl
2xM+ANJjaP7OJeTaHOSBrkDA/0ElGwn5HsekImsMdteNMQav6/Q5rE8NeYAoIN8W4Y9hLqKQIPFx
k4CjbqBxqI0fI1gtNiJtXLhk/Wi/Nx/PPDgxretM8j5TH/XOEJnYXjaGwMy6zn6AhgBg4eyyfnpB
3qMCPdTD4jUaEIBrAwkpDo72Pcb0abm+BlMnMhELiQ7PpO8qpjWKmgbIHoX1VvhpvJJzxE7cBIBf
il9IbTTYug1KaB6ycQ9sH/nAuaJJVwGRftpiBNOh4vIUYIXmMm25N4dMZwfdosZ0z/6+6mdukpth
zDMw+9kFxrMukqJmAKFhpZIzOyPHpmiHRx0VOzEiCVb2ddBjWoyiow5a0bm281M2L/aVwc2zcl6E
Vxy2SG1XIODFmZ1BUCFAGLcdmqFYmBi5mD+VVQTlcP4FecXu0xp6ZUF5Mq9IKueYZhCWudDpZYDc
a72An7jOsZyC6NEKlZu+Y6ZHkLRLW3qQ4jNHXD1M1+U0Ee8KWyaDbQD2JTIfjQfQRR0Ko8KoF90n
2lIgTtO8yJGWIgJRKOHykK3OHBRUQ+CMllHUZXgEc2NNSeb9wAXjdmz1oS64KJTKcJV9/NsVWdEG
734/qi/u+sCigqFExT3Aw6wQ5qGPiPaD3EsUANv2abaX8xV4nWfKs9EuSM64yhJSMMHukOQbLq/V
/BqcbTr/uz/5BMZpyYN960bCpl1TAgt1VYOFVgEw11AoBfmwq475gY88gTKCMo4cpFcxxS8B9mHJ
LO82VgZ69UY2/v2mE3ojvOAqLW0VA3pweRBbHZrELPxehGQNF0tMYMRkb7t2eWx2r6OXGmyzBTJd
zvVIViOFyDQbY2pxe99dVIaIDVUhBZP3LiSc6GqW+O+Y4b8Yry3ivZaO3hAwDMsxrO0TIH2Rhlhi
onzV6CoHfvpPZVpIRpOW6R/t2EvOXf+42gamxY28uy6GFct2JaHu7s+4BZ3BkIkoilQdQgdXHuUd
tRppHjy5FRKsET4Co71aAJpc0wUdw+liZWukJWBUGRkAb/euIP1xObmQ6/Ex+DbpemmPnd3j9dut
zEOnOOXHb6cK1nqD1/Daj4Hkr9z6KKwJH9SxV7vDQ8VQdcOeOSA7UEGGxbipgJSrKBL1/24qQuqZ
XyHnF5XYRkDjxgZ0+aUW0sblJB0cQ/ar1HaWz+v3PUm7vVyFrghol2qH8UUVmJvSGzeTZ+cBVeoX
ZiPUkxAtjBtf3OTEXIL4MMJCXU5ZRlw3Z5DMJPMLQesivJuyoiFsnu7gykqV71WE96RJsYKu2KKW
2w0c08xn6U8MWPmiaDtbAy8jTiSA0gfb54npoM8VL92YVswP7sVF8decNZRZTAsh8atwkCsRxZPD
7Om9wcMDYuXp0sayDDK245USU61V4x5DaYr3ga5iux+vuL6s8//X8JyGEOUDMLGcZYNVRIGP4gmj
Nux2ZUOaoGaRzER6u8J9cvh6lPJZ9YcKxMa7jirU5RSIssEvLhWfdAr80RlouUFYA01vJFpeHxkx
mnAEkfPhv4pyaK/oD/oXQ+l0sd/3DW7v1FF8XIuWokB0/wFMyjlDQROKWAkwhMovdVkKUAqAdQyo
fRMXAQFvxHyRGk5NE+QIQ5UU2b/En2MnKq5aziMOZDSI1KVV8cHZHYYbY20Ah7VWoQAPkbcwesQu
t9IVIwgISKuJ3v/5W46xy85cA3w9jl6IqGRfgxYX8HPX28VYesASZghcx4XhXl9W9h7xru1B/skD
/4R3ACS0rF9LqaOn1rDaBcwikw2zNfo+s3hreLaRY1EGGf8Cr+G6CgrgA7G7J0md8jd4Eb25cUxn
2XtpaFb5RLe7zUqNPIzEXdoYFXGqze8FBDo7VGGspsMGXtwZF4P3wbjDYrE5rNFi9veBmZOIR7mn
fotD2PLGK6gAiuGKYX9XermsiXwkJ0LI052f/nJ2NgVYdlt7832A1qNM5YnmRygAGOcEL8wAKPNC
QBbm5O0e9odoqpNsca9D/z9fzjMxLnuoale1WxS0c0jIXGuOptX9sCUqTpHAkBW7WxHRlZkBYCHk
xM4OyXzojplDcnnFR/ngrGOx9IkQiQtgfe/AXx+o6FLlm1nj5H8ZXRBr2GEK2+8AV/3TrLqjPAts
timAJDMdwFGbJCBF+yi1jwQW5BSOOhk2ktbqbLMEjN8+7rOF/WO2YyDXMEOTgf0tm/PD4L3gbO0g
fWLDhBkp4gHENj/XknKzOHtVsUrg+YmHCm84dSeN5egBVv4+MRyGBHXV4cnvz4ZVJCTx+OUpBdo3
MYAlqcpyLHdZgolyVGVV4z81OmC/P1MMsPodYSFPMx/Dl4c+x2v8Yn40c5j+6lEFeBg7cujPsUSp
eWDAmKlxnObXmT1ftPCNzqvzdySRNB2YA3YuFg/mOGesOqqWALYQypdl+olKCuquoaY5Pz3hPuPu
oHxxgJo3z/blNsOLQErtk91rbOW21AtKLSix4n27CxRS7KcFEbLj5hfDEbAQDM+gusmzCFq/rNQV
IM3DM9Be83D7y/575Uil9r6dO72LiwKQQ2dP3LidBMeMwXva/iTo1mcldFvE9XV1ighdfN2I9hcv
spyZr7VjGkRTNFTd9EeVC+DShNFvONdXPeucrD1TopDp+vkIPHmyPR6gbUiDO65N1A80Tb+kh8EB
cA2gpkHQN9SlbkMeuvVvxWRrR5Qj9zI2fdibPj7mDYpkw6+/qQWaKo/8MYoxVVuV7cpGxs0ctX/Q
xBYWbZN/tE/3BupMRYt30Pst53a5FhsRYcCvXgjzHLVR/pLpoKfld7SpkWEvqeT81C/J5ySRFaFC
Y/NS38if06/ponBiGlqEfAYL8/rt9oAhQK2GuRR6cUXAqEq3P4nMdS5j9ldkg9WRx3Sz5+rYU82A
JkESkHCYTV/zg/olj4LDlyyDn2VFG0ZSiwBOpnz7J8Tube96JPIq2X74xCi0JP739iL0iN4eoSCS
q2uuIE/aXoPNOrTAz6dVPaiBiJ+QxBLy4+DvkxMgl4PiLGF0spIJLrtaay10eqSDYSA4dWqqTlCk
TTt/a8Qno6ihVRf2wnXC37BxzbIQfoII5CRtsaldwoIfmYj70KKco75VtlqrypysmZ7CTH3ZGHF8
Bew778y/eBndMHPkgtbrId9JKa5uK9oEAc5Ser4ibZbJRkBVWJ9ErTHh9aGIQNTZVW66LKGMnhPO
Iv7Qlxyb9jkmoRkyc5y9RwIUctv0JWsKpVsCY5sOj/B5GU6hWo3tQkvgqUo0bD3Cbu8jlv3wTj8+
4GRl3ChJ43Ne5NdZ6JnTFUDtikk+ZFbirCVcaNNIvOn35V7MhAhMfY/TvrFWk9R3lzUkWa+wDlOZ
Mb/EszHk5jYO6OdqUuVSxknLeAAroK6tExGIZDLmravMD0bOZIaHjUaKEAQn7MW/LmwOhxc+etf8
BXPrpkTzRtlvXJf0uRQHvGdLHD01T+/5AKq5rpgMMo0XprTWY9NXASBQtpz91i0ehwEWr/XDmZaa
tmoiVw0jq/mWPIQq+jvxKZGoVqszcbzu2iUnCA24kxljJu2rxVbd9jMWRKpjAzRt881DFHlAEQt/
KWr3VutshPYz+T32ereFLL88rG1P3MKBhJ5SiF6l6Z5r8oIH3mNdbc6fawVE0f6f2vgo3bXhYW8w
gWZVj5UZceqjTKW1pQRvlPxkSPUUGabWzwiSO0i5grnsrwWNvmCR0bfPkhvcDtBSsQpxtTOyf3Pb
M9WfyifYUXWXbtX8F/B9XrCiWO5ouzRTnmiZ204WsEMuJf9rYiS7Dl8vV2tcUsjvm+ej3VWUMH2z
vhORgB6/lpXPslNaWMCfmt/pFziErSH1telYUQSpoUV+XXF/XotrqCpqIrgd9XCzrI/51G5gqnxP
c40AAl5vCiROaHPke5CE5yVhD2d75BiCewCGWEGdAeI5U4cFUtDu8XG8HqVPufwa4elWLoZkg2QT
vtPZT3h6yDjPW01KU8xby58Ytwa0c/te2dzOXFZJ2t1O6eOwQMu1zZwih/ZFDlGvKQ614gUMEHmz
zn7ZpLtiW8GzMPZRfV6eTRBmgqekym5ZECxDSXn5e24jo2DgtybRLEZnlVtYseWHQ6SN3XZISQ3P
yOGE4ERmgZLo3SHArURi03Ag3N+tP2Ow8r1pl6JULX7fyfRgk78PdlXB8hyHZFC93G6lMykXcVey
U0yE1R1Oq7AyqErwPTciYMZu61m34Vcl36B+VqvUibHGv1E9y16oK2Bs0yYjMSqW5NfX9a5pdo7C
teMy4Lo9/qrNtyChutFuQYkU3SYiehm6+z9K0Qe+g+p8pdmQ4gvkGKX+pCp5hA3VZ1T2lt82+5Ws
mhU6P6dVv7FLcOdRDstJIFSokfe0K3808l3LHrwHMNGw+3EggacLboxAvZWImlK+uhGmJWkBBnt8
2p54QOHzHM7PJYG/fWnCDt7u3kweQmzDTMJkfKUYbiTI5P98Jv4zXJ+VN+pHsmP3DS4FaiN4i8p4
8QVlarlu9uNSD5EiG3ETKWNl2Ix59vY84x9Owe4xnThKcv9iibH+MxMS6xaXcynC5Rm5u1oiHhzy
QNfiVf+3Cq9fflx7pVslGYUXKhn8DwTZ9xAyPMgGwelwJwyswUX6yLtF8G4xuXHTxbj2lWLwfKSX
bu9iyyD7YbXIq8APJU25cUpvJiSLhPpsRDtEVafO0+uApXvMLvwNgQ2/rQhktDxg9H5ixLwlNxe9
7AVTj36RcPxWcJE4SRaGT5U/e7cdS6utsa1KM5Yz0e7wTT8EXZ7v/TsdIlZvKhXAIaaUF+1gDOX5
QisehMGrWB6f7QxEkH+vRmbjDj6fZmdmHJhtzaonXWbAjEU6i/iG/0SxjM1WMxWt5dS6G+ICGg5v
xp36Rc/PJOX7rgq+9RbNKmCzsqK3I7ThwNB8l/qWmKfZwWOGHwwBMWYDiXfXo3HG6qu39qnjGfdT
p5ImDrwm5nKgwQYJkDaVL+QOEvzdwz7tLMPMw/M8xzGW/QUwPSRNxXHcuWw/vOVKcQLfrlPNxtKL
HenyRQdAQY0rmZLBEFAfo983q8ZXGMUQm1mfKAbupcFoNFzt1WYFIKD94ubvm1HPgZdj4XjLtb8b
j54Biwc+IlJtSRad1eNvu+Tefcso1vCzBIOeGczpEREZrDIq9s2zLkf+Hyg9AxAgsiWEz0Ja9RGd
nkcX+ogZbw2F7LCcOlwenDon5FIpp5M2DfBVdVls30C3muY63VYx0Hzxes9Se5WQ2TklNEK6Ny6B
J2Z3441dPu+2/Bnh1EesAquycpGiwhMrCsOwMPV2dMoidf7q4kssN4nVYf1wY6aM2+fVLxc8coKY
O3Q1X4NCHd9e3VNioSfWkoy04a09eNE0z5qSQycf9GGDW7imDXA1iEx4+teZj9S6Go8lxI1HVYNf
ggGvMEPp6Pdp2TMLJ/mxDafZH6wiXMS0VU2FAMlslMliCOqBzwAh+ZgxoTpNSPNAcVLiKftv4ILw
OJW2aNSwOdDntftykHvIL96RVEebqFFK//SuBID/k5i1hbCNC2GKIhisyNj4EWIbpT5N0n2YAyUx
cSXHxQpl9BRHBd1Wuzc8FQEW0yXPGAF9YHHFQ2XO7/SjA0ZEMlAwlcvTKx7mgBLnUQsSFAP0fHCk
+zVFej7YcajErXfvoClHDClZ/TTpIAwjM4rNUOT4LbzZkrX9X5v4w9AvFRjqZwVKdN9st98QSg49
YZFX1RQpU2XnkK1wDVZg+zXBT8LoRpM8iv1kgb2nT3hf3Lkh7set6NQA2zANRM3te909fSp5zCzH
gIeM10mgWHNg41MgpiSEV1E+7MeP0dVuv/f1NJQaO/XZk62pOqPmsGlwEVjTamqIazhfd1FAeQmA
ISeWXg53UzvMfe5tF+U68VZLx30xJ10ftOaDqrRgUymTejp416hYUsUJK53GY4bujWUEQoXrnBZB
/rJhnqqZ5XC8+KSjYQlA86fUaQwh7bHe6HupOwu52HVJF1VtOzG4vFF4kPs/ADX/XPLcyu/vECC9
z3lfsVLyN67rnU9UtI3+aUCDybBvcQqEpeeAwuLpjNTAYcaJn0yk4lIa1ASITiIwI0aTxYt35QDf
umEJPzdFmwdNWg59/EN7kPAL/7rb6AYLGuxNMG4QK0slTvqcSGombWNVBCzMhxEzuzNjqlI0B5Ad
N7z14sCo41l9yxk7FiELiPq5JOSka/KFPD7Y7qchDTr4f4ROlEp9z5QG07dO51YEPOEIEqoA0WWI
rn7n3CJPP1LiHmk5X+G2ip5OQjvq2QAlYD7RMJFLKRd3RdLTSHMSBJ+pp49dmQQ43qquo5YPz/AF
E/oojyJVXrlyKVN2ZzzgNyPi/fPfAv0xoEAZgNfG4vTF6RjHo8v0QOI0FE66uW4y6IBzZvPBwmPX
8os4dfDr8eS7CLz7K5jDLE62hm23lHpguJXfa3e0jtZhAl2HXDAjjVWMeIHegQWqxgc5cKFQ8qrv
z5l4uyRnuVQtc/LeKgaZmNaXvsOBqH6RkfLGBtepim57dL1/ClI3YEiyNAiqEGeBBAD4RzCpN+1c
SwUN8onfeBJlWnBLyaCfNKGQG7Ug0upVzgXZiGADms9xLFEoaT9A2x8kCIR8nj9W0zdxVWyl6svO
yfOfvf//tImeY5m0nRp26y0twuMCuaznEqvDk1EfsQmr50mZ8oNQiKmwN7FCd7GeaaVzWms1SiE8
DgM4dvIwzyTwFqXpb9a1bkWnfjK+I1vbIL8y9iSdqzyHjlFo6TVSJKYUvNOXwFUMJKn1jQc4r6db
Jkje2Xd6xSXR7DtmmrJW1KJohm1rKvdtJ5u7wVfUtc5HIxfnoCEVUjj5NueEdJO2/MF+pCu+7pPD
PIbOPi1ROnXMWrAj1OYdtKJuOjK1JRNmkVGRjOxr3Mgxxyn4Ii7zWwOiXxRLemfaOorl2+AmShYe
P/15RF5ogsqqBcJQ1ADyYQWsg5NQqNAEJkwhnTUsoqTl5WXViGTvqxmlG+Z6shjg3DjtUuGv4oXY
TRB7M19wKCeEi4twlOCwFeVCPRtDPt79bFhQDXrvkcYSF1q8VGoahEK4yl/VpQBc97AooK+nfI3c
5kRzT4GIoCmVzg0eKNCIh3aNXWw6xAPMlQwqpMfKV3XNXNt52aGlauYHvHPOi+WiJI9A/cfzK56x
f5/dGcTF+2iL3YyEqsM48uKWjNZfffHnmRg8cb8ondlMypwkd4O0fGHF2dUK04JkRy4X340tWMAB
qhgfaEXj1TAA8ovRdWQQO41yiCeOnHTps8kSOvwATmZGXm+X5E0wKWhZrlJ0+Qk7IGLUbDzs3149
GCTid6blI/mV9C0H5ljKQSFFvafbgD3uLcstPuouHA2BBoK2k6l6fxXP2ISkTDENgWqVtcJLcLx4
tPVxQR5++VfMJ+vSLRSfJlntu0/hsBPKtSJWH3kgXamlKW8kGK7Sy8y9CIfDOPnyZ8DYDERQ+Gy8
azlTujMGGfDdFSIihmsJhmDZh+TltFdXjJI+03NrOvu85NnG4K4/fK5b13DjF3P/TgvMBlegr3Y3
7+zWkWB6RHk9Qx3lSn00tkm33qUEBgCvywE8oLmy1BxpVHUFJqAetjBJb/ugJgfTHvt78l/sgrdu
rMNyL1wd2i8azmnDpKt1kz4EHOYQRN98KLgeS3QBo20p02YWQ3Y1AtMKl3p5+xOD2HrBc6I15alm
bSf2cFPCEOPDhUeFFcurdiEECkHO3ES56+LqRN+qDX17fFxnfA2+lb6QjOhyvAWbFuzrtDKgiOyy
l1TWlsVbHdQjIAaGA3SQ1sWqBSwSLQsff+I5ABE27/duXh3VOomW0WxxstKHrQoJHC+xe/KuxVKk
CP5oPZq8KZvRYXW1HAe44JFOIsVvlJpd1nuWNcmdio7lSJzF6V9KnIRgcoeHBOzD1fIRnwqMsecJ
zk6t9NdiBRwQjpMXwfEdAMg4tpBZp5hyBcqIUfis4ryh0U0lp8RcL1XH/8Wbdp7MqlRNMXdw4+K9
uRr3XK/YZ8kcJ/iFIXprl4uWuWte/zmv4I3rF46tsHTw1NSnY3Tz6YsAodKALREOQiRQTCiQTowe
kBAE2VizY5KDFGlcsDTXSsTYBZ/SC6Dytkyfq5/smovg0Khb0rFOHRg57QAyhjpbzUwQS+/WfSzB
tN3NSCQbIm+DtSg+hzL68gvPG9A3CDtu+AOCDqR3VhjiOpaoQ6UYMW9O9NUbpoa/1FosUgmNZauw
auYx/Wjwf2EUQ811ATKpZ0YRUPWxR+mwhd8de6ahm+v3jafabA6LBplpQKDlxY1v/N5gPdM8h1fT
K7DtBkIoJJUIHqcOT9hsz1Q+jtII72lc7AAn1VrraOqIoYgG6UdrIuc7NdyOuVC0hHpVRns2cL/q
lEUEKsVqKHAm+WEiwphVfIaVxW7s8uYStu7VEZeYeX8sx0a3tveKTe6sBDhNmhY1VTpiY9U8YRu/
SUYWfhIY7tM88NIfv2GwQnsixkQpG7zqcvNVnBvSSXRkeLxIcDEe2ld5UICK9KoJegaazpFkh3KD
h5UtP7W56uzYPrLXLRJoz8zNx0Y0lalmpQPNwL+Nqu4YgXjiUcQiRnztsR4l+yLfvoQqW8JM5l9M
Vt1aQ6pkpaUHwJ3AsJVL918yScQ+DB4PAdKuPCNaCKm/ExozYonZvKy5SwPGi1yM/4hXLuViTmXp
pbW+xF5AoHmNCxLtp9vCiwFsuVBFGHwmMO2vZnhFrORmV3cHpyXw7arriB++FHjA3fj9AEK2z7Ns
h3Je0NJCEYlDNvyzliJnGH+VqKrdCCFCya6Q54dbiJrecwreDIsC4mUINfQinMO2LLdNal9ssfOl
VJZ0zj0iUbOajcknPkF4xHMGthnLX8cgj8YooeYIO3z1ia0MKCl8/hR9/YilyaqXI8pHw1uOqd8f
mke7+w6rKN8CSLbZ/DqvOiWIA6aEGpCdWq7JT1VZV3/AiSDpmT6oAmSBusrkhDrDyj80YS5ZnU/M
QZkSy/huvd4eL0SpVOSHqzCPSy54uOx6tbAjlJhtIGnBc7uB1JhXZEouVnF7+JfJ5fD8vj3nln4Y
D+ITWG44KV0Xc5hCyD4uzGWqr9Q4QEGgZfxrVw5/DVFLPGmmYAGbJFeBOq6Bqo65f6r23RjMah5b
c11s8QxPBRn0R98ZWJNon1R/eLH65djdtnN/K9EaO4hWr6egepmFOnepPq/mX9WK5fa5O3AE71xe
iq52wJI8XqohqVzL7Sm85+9RisfiVpWX+uLz0Q/XD8AHVy3GjqV8vEsxBRpheHXONh4c/xPszGh7
crew9IN3NYsCzwT1imGvRyZkoVISeaitlUEOg3trQCqRhWvWGwzqd0C+m1UmXvIXx7zQk7Yc2oY6
7vYbDjXQpnALOxOO93Q8LPEBI0I+cONg8cc2U+22fRXhdKBI4qypZdVKimDaou0sOwUCeOZ9fLoS
B0ewbrgl1yk7GUArgXXvAgYgD8l6KAC5TrnssT3JsJnlllIIt8cPcCG+gawxoC+9TPou9rji01Yd
UCweK5Wcudef/UU4iegh7bQph5CVEV0F02x9N/qip63QY48v0vnu5MAtRncywm56TPSltpsbw8pG
tuNoioYLDSuxNo0Cf8IQF4BnLiN/UgfNfRdjDQz9BLxEjJniSvDF3dCqoIPuYNvlEvPlyId+652E
rlXsgXYm4ESekcrj0LVap//mIqHG8O6pkl3WjQxAAxNu0ngpAox00yJtNe9ER0wf9+hlZXIMdLb2
L5dD5vrTnIiT7LT/5vTxku7tObir5YgDMSORqW/h8uJrxkWScXuvqQBcB/3wQF2wU69nVT8FZcPI
ev8bZ7ttAW1Srxv2BT8QIRWt7RhR6pvbkJOAAXwr7IxerpkVvwkmd2AeEBfnfZKTS9o8fxSBW+rR
ArKflzbKtt8ZeI/3w7UCGF/2J8QU4zhO8QWKig/ZjT2cPDh7pLhbKcJ3J+YCxokYei+jAdwdIv7x
YHCiWL7HazLFn1EazVCNmrCLUG+01Z9vldBcp7+dV/LAljUI100+1NdZmK/QCWj+KbTP0Ja7O3QV
SyOkVpHojievR+dMB9LCxaE5XrCO7UIpGm93GU7GR4sYoPGyMqfWNwFaS5kNCDAriyXYppuYVeY1
twh30EcTXmc/fGduupcMl21uuY+sH4GkPyR5DCaXK433npi+25Z1D/qyAgGfbfkmg+qTQhioe2mm
YXr5SE/j1Fu3mVbmmwTWYJrD8TrroMfc6RylBrbL+nPlrhK2np6BANLTv3j3BtNfxBmr9b2udem1
dLl685qeVezLCyOfUNbsPUVGS8p13bdRliqgr+XcW1NxcadfxawA1Lz9LbECPcOjg5zbV70XkOj7
UB9N4tekrsqIwD8zdOy9JZYd95q/FxMASuRB2ed6TX4KEV0omk9k8IHgVbV4zlJzF51haMFpHf5T
tPZ879dBoxZCjijftY8TdHL6N4RHAOz4MocmAHZCY/V1pMm+ue+UUoi0hGiUF38gZ2UI6KTbYu+8
cQnVWvzwkjfYCYlvkdKdXgc5cW8LCfeBhpvihbRWuQrtPvTa82GZhSwS0Jya7kS92ELjaCUhUjRN
5R5COvyBzpxESDj6haec796JOdPmrNQR70xbdmI6qXgSkfH/XWsszmYNDNDxCneel6dSpvscpiZC
hQgS+h9k3XEjTl45yv+ZZxYUy6bVa5AW+wOZyiox0CS3s/GnWnYShpfoQK1e2DZv3iuMu0zdS7k9
SlMXAVUrOrWV9FN6SvfV0SalCsAGKcnG0GWpjH4RNT3nPUYP5RtG5f/bqxMFKiKc0A4UDRws2Com
58VPDzNgr4KNVS9T6zrBRNBuZxpaooqv/fseNWZXRbQ/CLu5RgkRBiYbFN1lRH/YIGATUeEDTG6i
wbP0NsZxb7qx5A2y04tCGu67i8BKvchIugnarnT1EmaHrKAhT0u2TCSoFD61AmITqMezszjxxEXL
DcFuZ4uSu32OWr4E28NjiLi2cNyFyqmILKoEhkB6yzW0t4ugTIuwZIItsdK4pLSxHxxyeejPOEqP
mT2ZbwjYgdbLTdmw/qwFw6usyJc6TJJPZ2+wpaiM1u1Hd7EtyZ89eimkMXhZLq0RTAP9lkcYDlUy
Vqyx3/JbKfXCRZ7V4OpPjwUgpzv11KLFs9y+iky52K6eFZBydTRfq4i+s9TSbPXrg3Rcs9XAU4mj
29R0GV4RFH/f7T5b3sn5P1F1EdId3jUfTWXa3Ju/5LkMENFiryCmisFB+zYpu7W6f4hrOTiDV42A
8s3CAunucZcMPSU2BAhtM0voeUjKToKEJXZVM1CY2pxsmhg3PqC785tMyyEdIADxrkKqoPiU23Lk
i6eFcXvEiS18e2yYtfBilnjzAdgduYctDjK34uav4UulLWV8aeq/wkbvpF1B9ZLsaoROJ8pBptI/
Stl4fqS8pNjeF7CqpWyxHTNkMzCkZwE18X2FzwChKWtDITf8vEW1fLmOu2k2MfcqiFhsDv8096es
p1WXUpSy32dfz5bsPUNwPl/vMPGXyWLB8Jyq4KTtD5irNxTaqii+60t4n16Ey4E1xJbEyAAElXqQ
swRxbI6cOomcDx84IR0uM2KzKmcRyH85bE7gccYdxmAZmng2WSx30+LRZN5D2Jr2iNxSXLIzfo1T
t/cDNhm5OtSw6yP7NyuZkB1JVqlejl2usVBoYFypEStF5aqA6NRY547VMgeTtbJIrSecQaiSFMcq
X7QMbj/7j7mx4X0+PddG8IaVYWUZXTfHiaNQtqqXEG5PlgAXui++QEqQeNkvUSvObzohDdmzNOSR
Sw3etNkkSpuWA4YCSvzF3o2O08AJPcI5MTKTU7VIF7xtHOSU0FIupCU5zGlN/LFolOwpjEME1k7Q
pCUlwqQ3v/Vi2jNm3Sqh7W+CAkBqIgB/tQsO153M8UJfZ7T+cyYs4ynOP1qpejvyF0bVp+iwQF12
gI3YAYqBDeE4gXn/5fcrAMx1oyrM/OWQSTfDEV+sM12Z5GmSnrjR+oIK+C1qCNumbxeDXyl0mwxv
sdNayJgf9lM41k+C0q3+SWgF8qx970nn5K8LsburKePWM5UQdyMLLKe/nMrO4MLdX1lEec+jUNTW
+47S7gJhmhuFeSVnBauy/r6sngCHiWf4zHC4XskZupRJ5xteOkDAchNdZCKG7ZPrAsfU1vZMYupr
zxrbPwwLegeqwdJD+FjPfX93+mz5wYu/pkkTs1l83V8no4McXRM0DxtfmJ7iijkRoJCvBBntBHzd
rk5Kq8LFzuaBcu/xCO6mVl8FPA4vUoBMoPstrATF3UDRxPjMF8odpE6DgWxpBo9jIBdgSaraTK85
v/KqC/+eSn186xx0/+Pn5j/4sQ2FpiwOyAo64BRBdWbbzRD7zDEsgiZhjFmbOjkufuOhCf/DgPnm
ZquVj4DdsjcyN/yahxoTOtQX90q+90VLKw5Vi9kedgBwwIs5GyumtHRbmQJClhi7hqA3z4+9EhCZ
aJaoSdqEEeQPtiENN8EhApNPPt1ZGguwaE5HzxtscjW7YLtwBNrAq+UYe78Kf3HPnHna4YF/1C9b
P71KGMmuli+1jbVJeiiuwPLieAbyVKM8wORdD5+I4KNPRtlfyVRTE4/3ffikAhZgRltHNfSp+rW+
xxAKdhwYX0heMbSi6qB9sVdtxNgcqLJi0p3u07CZ6GmGO0pipYuI+z5nMi8btFApRNfmG81BAyi4
xj1ogAsHQIjDIxYvADIH81joTsBRwyj9ICOgvpwCzOpFzC8otH4s5IUvvvyqqDg2frVsjLklVy0Q
SQK5SipSpuT3qgzUgxLP2ZN+yQNoShct0AAc8yq1wiL+5SWzRUgUZDCmTM3V0uJKQJuVwq4p1cmD
Dz/4kqJx9Hjqs5mTVv2UkOAx9p5qkCprgT8hxqstXbDhabWtreKxgU0hKgZY9KS2HDoUu8vOPkE3
+Qi+28qyjk7MQiJPdJm4pXSAdp6jNXJdkg2lVKx/VbWRQzVFJp53u79lAhguD18eVhILlHN3EAra
ne4y7v5R76GDWOAlTeWSqpocVLDtTM2wXEbrN6PaceqLJ+bdEDd2l3XRYyUqPHKhxFlu593SM/1s
TgzRSVeTRh7yr02uIUO2nH8uLYHkqbASLtTRk1LivODrw7wVk1ZAecTzqirmRUCbZ71P+1Vw99Rj
elYLIH27cnm5ZXh3biGjT37c4rJZcSuNXO3DZxmdWw0+76FpdJLAj7QHqJ5fcraiJIFEUaDbU0go
8if63+HRu0c8kINHDAYIuZM4jNCu7TIv1y3CUKZRUfTzj087Dxcn1Dl3Lr/9DNBG230HzCtbA4oo
qMqkcnQwipRa7gO5yDyBnWsz9USyZGYJMykN5E+o+jEpoQQrW4Wg4KWbb+aB6DxrWFaxFlo7+A5x
80E1jnolmEoCD1t6+ZSUBx/6mqbV+zUlEh6m/cyBl0DEuOV1n4SXoOmJGepolebtPifxsuSazGGE
VOgpTc1IrKRTb/ZxKy6w0h3eGinrvDnyNOqAsygv99w5JMAarOudYbawA/nPRFtWg718lb4myxuW
lLcw71dqcAq9o36jRh5VMfI9D1YG4nQq4ZKfpohR37Q/aa8KS3eV/s/cjpKHYQtxCCgeJGYSsnUL
KFuoC4zQxfSNR/rHKJG7PTYvZvBzkqQaEDaLYt3W+VuBv7PF/7FbajhM5h6WoBCPTHzIELIGKLYZ
Pd+ZoxUtAZnh/5ZwVbIXjenVy9Gq23ZsPNKPdI0zKvuBlivx0HTwEBE5oG0+ZD1sHTX3NS0qiNil
BUt1ChDUk7lqltf9RQiBbCvate/m/tMHLXGobDgXAN9kuqqmIECDCmlFvQGIm8WEsFJI95nafpY4
DCw6oHH6QgLRfJbQ68gXf6F1wH1pVKd0wLqeSmN9oXBhyLqoBE0ZNtYV7NhugffEGzbetClUseod
idavTTe+S8loOzCJtel5dhTscWIhKQrvrIFg5DgkSsu6aETrNzPp982uFlcKIC6M78ABCvxAAlAk
F6tauGS5wpGkLtQ87xp0H9Q7A8gTbAr4okQ0Ej63OJhsDOiSKHkPB8+ojl6B7LqjceDYb7rM9dHw
JNWbG1thhlVtuyai7DQYTVo6AAvfMaaF+pM4xPg04R2ykgCgTeWst+a0M5Kby/115ogSinZQGXRx
XmRAVlRbMeYqBhxOAoZxwqSvKkuQS9a+bJTTiOIpo7uafPWGXVUvnwDLuuNvDeozTDTxcxTWFWSh
TPWm3qQMLfP60qLe1oMjXc0HrihWxc4YGsu/ehxa7HFo7BpwopZNsj+5sN5HZjBbTsfAoQHt2A1p
54irN5npGSv6HWmMGe29dNUAVEg+wrIAVetYxns+NdOBile9ii6JzgdvjGw8fX9C3OPBe02mxd3D
lL1dkWNqUcxBBgfEt7Q/DfQqkczlWObY2II42//u1QvIdR4rj4OJ9mDSIN61h7/X383TuxXWLZzv
aquE9GBOTXHG/Oj6U3LSWAgua8oAli9r8ubTtUnD29jL3cidHALytQEwyf71B/Vt8YUFQO6fVkZ3
NHCmZpUg3JJXfCA2Mncj72H+paWHhMfH/S6wEfDp2EZKDopy9tUQrmayKey6X7YYXv2ZqBZT6emf
0W/FbpkTtb/x3HWwA+LTHWz/s6nqzUV/2F+f3W9qGeC2vrqzcSgWJvrY1QHDriGEP1CfTmiuvqLX
DYnq7y4oGdxFB8iVULJU59TVwQS3zNuLCIxfQmv+ymsDLiDtKZbl/l+bZ2dDJAd0MLjkDPqCHNVy
V3dqbRBISPiVf9nUWeZpGc7iNqQjfWXBoFFrV8wDim4WgnEHEU+SO5MUmmxUSAPpnvWP5StHWqMn
J5Lt7J6ADnYhjxShwfhPZc0SL3H8tGujY/GyKpQDC6lJm8xOeHydez/McpBSli4PwvSSenAuCon0
OlAA/1MlsuyOxKUvUF2cF5l/g/uB8GrNf7AQkHSrhh29sJKuEPwsDOcmudWU5XdUVDENNIiREcoz
Py5hS/9Oks0owDBuNOp+3IkDI64iv2AQzW0wN2OvsyMLMCQSNX5BwggLuAed6khp4340xcHhDHVF
L8BT0ypFNWBkTvRMlBUxR4V1sE6LGX34v7IsLKJlynPe9MMlWgzGuaveDL3YNJSysAnPmaM2NFbk
SMJc5b3DkQbpN7OkD3pVTM5hKdzbUP7Uq8xxDRMSKxBwnHrIjTwtN6+BvgCOknmc/wzPrEQ+rKfB
C884XQLigSH9JgsMzXJCECWBVTYnJi2lOajnfEQxdF0pfTzlLEo84ec8JwMgPZRn5nR568wBvXP3
yOrlI5XeTYK9Rbbv77av8jhfNXZgBtPtzHy7QBozxnj93S21yWxw3kFz9JZxglyM83uY0YYiVgIv
y2BMIM3q5yobtFG14W/hBFpfjYVdwUAQkVxJtLmBNsHcknouIomm4hqr/a4ocYG6f94lcUmboXHT
312fbLKoewlVX1sJdIvgKXjJW8Yugdukgxsppb5wJSLWBQGr4i9MgRN4+PyoGlOkJ96VXxT08Em6
QiVbnpGpdhW6UkB6awz2otaL6qRCVyECqp/78dUwTvyqEqFH0SVXnj8AYez3xNSGlfpwTMk7f6oD
3KD5nIagF+qGBmaKqyRF3RrXWOIV4AjkfAhiiBuuc+BgzVMsNfDFwpUVfinzljLjRISljCKDlIn6
+925ZN9lpATvxdSUbLr9vpOds30c7pHFX/P/lTrryRk2usSa7HKeoO2Cn/PFynlzhs8OVOB1yMYn
j5pVnsQ4ARdwe8BIDztjAFRex+a2JjO3yfN2SNxO3IJ2MKWkHFsjPNDamvoCZcKrOFheZrfhwOZW
QU5wB8g3BjLjhzkUUq0qEku730MqQ9nscz5Xem8uHgfUAm0cLRW8wmfjJI4YJ9xp9v3ttxTLcPHf
BIS/g9EgCJpavjXX34JrFZBoa1xlWhQZk9MUxQeCcgsBECI6O3PKrRsNE0Ueb/NPcyRejvM6bKN7
+yo9NnBebkIs6UxoCta/sVPLy6NO/Y015sg2TY1Jip5H2VpmvHdNiZn+ZzZNhvaOqX/RT9733TOj
jxqYmzou68gEGJEwyNw6ovrtmgRdhZxnF5eNoD8QCySASRqLYABQVofStYu2wh6CE+BBazSH689v
IMjJOxDikxa2tb8hEvCFCiRs7ypDQjaMzr/1sZkrSkLviWS0WayMjAai0EnHMnoI4mHopt9l83Ee
GOWGMm0jNExd4WCoh6knx/14Ujifvf1fJ0gTQ8DFqPmHsXIdOh6BtYjB4JRL7Isu9y4H2sAYFtC7
0AamPpESTthq07jvlcP92V/o2aTKcK+4+ZbGLNvd4lJYcKYVY2LLczDOwGr6UVki0JTvKHlRphM8
MjRZPcUwxgJ5GMUJf4YcsA1hHOOwewgphUi3vl+wvHxbcUNHvNINcDEsnR05xD3ib1ztRLKi0PR8
redVzt5aaFUVqJkU1mMGp8DWs8Lt2axIrPOyPact2nJxrlngHmtYpo2T8UYr91SXalRnD1gts9I2
1T0cZaKAInvXjDSdFlbL2TpqnDBGvA3pQ928Vp1VjyDJsvGVGvKVxbGMUrbtqQ5/ZfRf/G+01r7h
2hgYHbF2OBt+wTwN46YCGpvl8jNVOn7rwXyjdTvHUnGnUUuoYDv0jxDj7prexc+PnZ2MI/T2JYkY
xoNctCzA8Z89GZulAFdKVi2FXN97pMMuoKOQdErGU5LHtGNiLqhhY+kdrYTsYelvrhqpqyyV76PR
n37oArVioBXO1KpHMqgPZ6/MnpWuKNfRvX/MXpDjRE9hp6g4Y5DpRj0UzzYJAlSGfDD46WmmJoQY
o9uE2tbzY3KlpFCEX4vlQF8WESbe25Yk9ztlyDBp+Ql/MWbSPbvL4/fZgs+aVCgM76JZ41qCIVSy
v7ry226bFAeBHj6lOTah7M7F2do9oaq7Dig0BGGPyrjWKoLU5KC6176YOTmdinFLJPIEcMvzrMpm
D4w4jVZo7cIcarnvZ8j/lQLo9x2vMNOvOj7Usu+FR0kY5n2Yl+nqAwEFT+a0QtNTvDOPutXq1XY3
q+Ueek5sXv7wMm0r1iutvv19WBP2vEyOo7u6ulx0Y3IFvDR5lOHYOSFIv94WyG4ftjCGESBzzpKA
U+AVOWxM1PmVwM8m6OXPU1qeR9yj81uCCqEh6ATuFhI1WA1f1wfFBJhouyRbZvXvGJwyXkbyKUdV
j8qs8OqDxx/SpRVCl6jv+MGzKiiCx68FWY+LFJBoqDtINwqElVMuZxlK0szCKLJWRHJxgEzOhgrJ
xWqoNL8SuwZ+Zwge0J/ctHCqlWoXcPRGj6NZOshCMG1aISFF5MYRZZRjscdKor+/xFo1ZOWRLQDt
MfxASxNdDRRT6CDezcIrsi7ew6Mox3bhx4wlWyHb9sgRfPP6btTmT0W0mecI7OZxlrYhwVbcm0AS
eEurNer0wJI9UnZvFXyhOhM1ISCfIv1SID2Z0JYb9CJVEBjg+u5CBCOkLBiM19l80OKoUz+WxJFu
H9z6HGamiqKdaGrmd7ekjFn1aIvPcgSmHZDHp/tEa9pNyvFpsk9TRMODXN0zIWirMtsx6D1bINjF
OqhWPEzQPdPPMtZgoLt0XJwb/m30hcclADyvGW9KEPTKiD7sZqEx5QJaQkL8lo+8AWX8hBbI+Yvu
hP7r2m7duD+f6rmNO5WQPBYrLhUHzNFdaobRqkIAKmJ9ZJ8cuQfuRIDTxr5R9q0s2I7btoIZvv3q
9JL+Ri9+KazSjN/4eJZvKMu2BA+nHEPMsgKtLY7Pvso9D37Sj+XS6krcIfPbfdpIe8dYHWn9MiaB
5kmqpAJ2szhjNavTC8/ZtclOtaYY2gSenSpH6HYNQuPc35NqpJ6v3IWJdtGw7K3ED0DdojlvGlxh
92Da9kYmbSUZ53dNrRiPATiycJyMIBi4aEjOoBRf85FJEDniTSCjklU0i+eKKccNIy8kCe9ek5Nj
0w2MhQ5tBSnXNS+1oRWKBy3/vfUMbBBGkOLWESCs+6813eNdaj3y7Q1Q2kHojWuac6ow8u+vuWKq
r3y8iNeX0Ex0oWPLuwip2K89Vh6GQq3npwNouegbM0OsCkyWd4oXSaoe+OILwd0/LxdijcZoDDhd
gP3/DjfPaBTKyVWy8yTdU82JviAS9f+osP0a3hCwGmlRajwNLrfHW/n29NRlmAUidwyiEjfFiv3E
Kjj1bkurI8w+dWFtq+R6IfDPQABUOB1DH47lX7OX98nFJz8wqsvVzDBFUmb+SEC3ntIadtyn6w8q
P4NCg3tyzq/CMSd0QnJHtNNp/gHsBxrjPJnB3WYh12wYp2BTmflaC33IjvTKtMf7uwAQ9bN9zh/V
d5RuGFvVp9bbaFyA15hQdA8O7zRSEaAczav6M9pwQPgBM3JbJfXwjwq9WqpYfKWezDxr2n4eqtqf
Ty8mwRvl9qVmXbdr6cISn0PJW5Vzyw2OCmXz2QqKTW7GBe/mm/zchUujm8Ln0BV4r1J8FWIkVOOA
7D5+jvtdBWnR2HsHmK97RVjh5ziyvvriFGDqpzH7IzZKE81CSKp6SL1oXEF4CC6+zvZis//dAEnb
3weI37xUuCVssahKspTygCvyqSCngdM6b3x3/IPJ22teRsCtkrboSeI5y4Cu7hCpq8wmKFP36K8e
caFQYBbK20qIcaOCYivNIEpPvkHLzHAhlrqGgv7KpJQ/NLk0K0EuMvtgqfkCz68oVyafO0A60/HK
fiGxVLKXwBePey747drPsVdQeNzD62wE+NnhBHpY56URsU+m4x+Zqq5aDyPvS4J17xUEQZWk7sRL
DwS7SF6zJxMptheA/fNd+sc4+H+gwjrOZJ5PRKiZYdZtMCiB25j+wYVLnX3kxhujwHK6M9Dwwdvf
JHVAf6UbIXy15NhLGiH/VjXG5h9Chk23cLfrUzTq1vk/9jx55eg6SeyukmlUWkmCZeOtKXpoeKPB
lTtEOhOSgqD2gnvBUrevlTYhToXL47a8VSWSH/Y5E4VT0Em9AeO8oUVssO7DUyemPm3c4+4z6zYS
PGrA7x0SzacuQr8MEdfDzuy5+uFRtZ6Br3XAHTY3vI1LatfR+CSNKs+V7aRCntlfhDt+7RMJF8wo
qdF2NTIolCDr4gFSAEPWm4tbVVwBtpbbxEOLglilsb/736r56nOpfFTYe44+bY2jgXblN/7mhmjL
DS69cq/+tO50h2yUmIvH8nuGraCBzWJhtgGsrE0nwJ2MGhsfQdgu6dTKuJB6lDCGAKmWKFljFV0/
QRcaZ90KNMP4KYuVR946puyOxBJePcsBAYjI3NAZFn5840XgKpEj2+yoYIihwn9nBLidtpJM7RZo
DyUF5v3K0KcKWO7IP24ZLhtQGDx/Y4tGTYB9bh/Tv+mJO/ZjzaQkTF2jD73zOIy85GcnLI6c+ZR1
9TxQzHZp1Efp/MPUtMYP8eiuwfpuXvA0bu9QQvEoVcCWAKBYhc6OjHwHHfA9EH8wjGb0gJj/gOVu
QrYWF955zzf6ohTu4u9pWRzQYcODjikmbNGa0xO1ZdHUBmnpc8hjadCX8kF4gaYILcASfMu0Xhwt
/P8u3j135juQUbmIcFtkxpYH6gwElnaS9Oyv6o0OcFUtajJbpNMcoalAfRyfHGEzSeBU6uY5e96H
fklzujmpMM5rSwmwOMxycM1gqJxX0MFm09ERyhDmF5Ao3Sfy10/8rs2maUOteF3snoo+tU4ZkK2K
6TXJbPtop6VMzcFyoeGlvcG9YrZhVRobOAGBzu7aAQPh1CHqfrUK1r+JD/i7+s/aDtNLxSPwCDvK
A2J2kVTGa8aVmR5xHCiinMNw+tGxQCYT5A7XIoglTW+dz4s+5S7EHZngaEgi8ozd7hyO6ODnX8KW
vOc1H8CoDNqec1w//uwoQvT4ZnYyZW8iaT5vUur08BBbjSPtL3Tpqv/eCblZqLgd+Gr18jMax7/u
D+p9G3DaqBgapvO4lT9bIRsMJDAAgc1CXZvsvBwxVbS2MnwMt+ZB7fIhOiLlvBPemmNaMSyqZnOX
ec1d7fE1UE0T8oT7Sf4x5oxLame5LaDmR4O+o6fmYLVML443uaIHVTHTrRmTYdDXezRR8xuh/t5Q
YReHoGx5Lb2hrJ6e5dw4A9kpvNR2sh/qTQhL3bFGHSnrUGbliqrdri/fnw6bWVJXKVuclDPxE4KG
uBgBCMT1EJa1bkc3Cbj3pkX+UvrjGyQGQADj1oxIay4fpa+1Eb5m8LRqd7Kw1iolQRMzaojMgimG
QpSjyjo8QG5JafC14mnR9NfivWyN81t1XIthmCgPpIP40WAHGgJNx9Zg7lQr62kedc7TPEHTGfix
VDRRWduTCN0s7mT/cE5Z2cWLHaQDq9XM0lQyekfBIcj/L5AZBkyPK0GihsmYsol4qHmSbVBnVD7a
UO3KfeMt7xS5Tcw4o40r2HTvvsLGWpOoFNa1OAIwE0xCMdyDxBU4DJAGlHkmMwgBB/rJ1o9fJ+qu
7lY8a9uN0xd79HiA9ljzsZHRMg2gGgWZHPC7zA7UOmm2U/IroKA/RqVAnIjZ8mSxfU2iJGGUbOCS
9kpQ4QFUelcC0o0zDEz0JqM01YC70dy6RxxYjl7PpKExZTBQEmHmtaQEDwWMhvg/JFCTjfbn1rB2
9UedgBkoKPv1u1B56LJFfnHd8mGtT9MoMwCwz0WhXnV8er9FFZ3eSjsxWS0VncvMi+blNtRcxt5d
AQmDBmUPl2WZP7m2zvwjDdDXHoo4mVlARqtd7Fqx+ZSbDu5C4CJO/cV1iI+bK4H7xVyZxBuAvwvT
agZUVD0F1M3T+3l1hf/nOiAxiuKcmVxNtz8mlnFrRjBBGDcoDrdIphshCGlW0DMPk27PTniaWdDo
h5HyPGFCKWiDpeQGeLCqYSnzCWtgxGNhpAeAX50lrBwXd4p8xO6154bk+G/OQI9G1ItsTqae9rs7
J1dOWC/Pwsj+QsTvxH4q8PtQd8jjZFLqIruv6oK026zMh5GuoCfq0POEINOlBbKTBrvlHEOtt1bq
ox33xCf6IUEnEgDympu3MNlgvmrCWufK6g/l7+OLCgKiGyD4N8/pSbvu1C5Wj1I3I2swhU5GqnCS
K9UmMxcfTn3tbSYsgNPMmmAVsbYyAmRQkrs4J+eL1iObrDeo9U7ej8sEfvoVIhvdfCKP8M65KaO7
l3zx6jyHPnLpDojQ4rV5xCFUx7suP5FMzO6eeOC3T4NANuHymSOdwK5aJyiwOZVRYP2jUnFp/hcD
92QuQpbt2ci+LfxR8Xpi6UnsRQC8G6Y8mV06BFdLJUnHI+1Wm4uDzhyd6ka1S2kup71mF8Vwp98b
HuAeKO8k4pGF9vagkaQaO7bPhHfLSYTs2WOmwyvkEvOGkqGYa+RBq2gvN6FfbbKJxpCS+cLJ+LiD
4KsD8vhIOE48f515R6GfPApgGIn9QySVIE2DDOgiHnEcDizCA+3eSXgd3Juj49SomxF4iOFpW61A
LmrZu6kLltmjDPZ2yNznvlzIh4XLwWzoEq4fOt31rrXxV8zdmIQlLO9Y83dvYo63yGoP2w28wbJb
mg4F4I2s6X9AGP5fiS84oxqA3r4e/7bz5394d5CP+c88LKv9MmscYSIRmxkvEKTH/6tz/nIZuJe+
BX/BkggxhoKwfPQLUOkSGP5Y4qVrNQr7NZTO9LLbvtcIqPsyA6uUmy4CDGpzwAqEvMzK8oEK/iOx
LgxSpb09eiQ0HmkWUtqHV7Nemz1CqMnwkthTuaut2oebzfrrC5YN43u7FbANDzn6VX5uQ9yOAeMC
EEmCnlV1SNJmnZzDHdEgiy16b+JZTBPBfYD5BP7D/EcVeZU1V5bVVwTSnKPLn7LzOnTIfXOfWZrN
4QBcEGYRsFornP9aS0SUNw/ak8mIR75kTsahkuse1/r7eLaeXV6jdH10DjWN9QJ+IywVz8IRWXHw
Z821Okf8PnZGfm34yd7o3sPku0PQB5NJrn6Onahys/wj9wM0gMW+gS2ooMHScLHstUFx8dmr5RFB
FV1DHr6rPxWDzf9LHRCyVk7taYE7Q6ImIndq/VyX48LhNO4hImtBQ3ea4R0gxioH8nHVMKZ4IK/Q
ryYSZU0En0O1fKAcPnFnEJIx3be2U7LSXCmFQl6i7ba4wR6qHwBAqrIhHBjJddKagjApLqNEEwb1
cVxZ2QutHGrzlJHcKQcGS1YjtoCQlGnocc2BbJrdMo2ncy6cGzqvIKmaBd7bpZ+vHxdbc4anqDI+
AZy8Nd+joc9INoCkO9uR8jjY62iI7srbs5O3PdOAHNJv5Gn6ZoTZLpdvHfxABrC3sm873SrMCjT4
I4jAHwSAWNnFmsywhaKVkB0SNE17kuA4GLeAbh2DQnxy0tk6UEmfg6JuwQWCq1jBl6B1p+cOMZCJ
9FUlko1ImYUZfSgi+12ptPKRNnt91o41EKvcg1z6I4DpxQx13qry9/7TYhMlhTR3czPIqy/gbCoO
4XNtxKtDOcMcuoktmiXZ5PO7G+OR0ww5MZddQuSYck7k+51qFPONO+ViWeMHq0b5odrnLTRDw9lo
oJ3cPWTx0Y0GzEhqau+rKOUy/4v0s6nJbY5btfSrGZLMi4A4SsMrittIeTkHEs2gUQybGvc3m/QN
lCDN+I6JiHwEpHU3g2A8rfiWYpbGGeILLDoHAJJKsVF/YV9n4N+zGwiV38IXu1Dv5hKtL6w2ZWoM
rHyDmDomZGnPy/Q0huTUYD51bRA6xrOiOcQS3pL6lVl82MdjkXyFBHXUGr0rzFmDf7LECW2mejst
aMf/53YpX1XI/TJ8T8JwjRfXuJgryKJWqIlx6A43QOkMJjugCgDUN6/hyaykefExJ6TAENXthP6k
CauPp7iyPD6eJ3Dkl/P/iOTQFxTMh2fQrdZBAYOE6ex5c5DX3m7zn3on44OKau4sDt7OGcXDhq9R
Q8/q8e0ERDk7aIp7Zap13pw8AdIL+FVZo+8aDIR1ikIlbk7iPjWjmEo0dosd/Xd3dKgFVbdHDOIj
XeyLE2K7F6a14iTxAyAbBcWFJU+iaIx0qR7Z7HrnEgRuHY6HWZXiAovHrCySteroFqA2cMI9TMLT
MNtHWwEYZoVEZI1jqpoMf15k529WyfRw0zfOSRa/+YcTOTmiPqkdLnlthb1LxckdwyEDUr5zYqQd
Yua3qBAGkR8S66myNh+y5+N9M+PJ3Pq6pPKyWVM4Acs4R5AcRKXXqHkOqISR8+aLPb7LsdfpfVQV
PMHoQM1IEF/uugRCoBp3XkFz86NAt8KxfryeiX3D2C46pSj2Py+4a82kBNZyLGzI+j7dG3UJaYTF
uKK3l41plWNFbNI4ukJD1AlfSCiIC4yXmb8KgM3ol+JLKYMScuV7mUKRsNXW1C+IPQpYRCEXmu8r
hCM5snO7aVMAg8u3lZpNbOk5QaDPeY9+1FnjlOa1sJwSzUF3isa+8PsTl1irUxstU0NVT18CfFit
H9r28DtDxN410JfDiIgo1CYwSQu7713a8kl1kRwgeU1oJiuigTbdzyvMFFP6inA0+q8jnLqRgkMO
KdUj/mqqiIi0W5ba+zQ4lYmJHGPj49mArOmU9Sd6bzqvSZ1xf7hqzz+5bqCpCS3RMBL7oNLGIhHE
e8valrqlF+4vYzWg9UAbRZl35y76g5fuOUNQ7fPgbbzf8iFtDKSU6CeNWtxj/sA4ZQ/TuWb9bJRh
pDDnVjAJi8pGLYz732HNv+iNI+O5Zda4TS9MepQ6tZbQydqAqkl+3Fi0udhJ3xpCqtKN3axIhpR5
L2eIVGvFe6Gnq4IngBpgZ+FaXzx2anZ9r1qYVhDQ7yXKH1JAW2GEOaqJG/xEmNd/z6TSKaHS5sGJ
Yq7vFZN3+amFIF9UJWjTdhmY4h3Dx/yVHEJluA7S559nXYjvbJI5ncVZ+LYITCnNHeE3KZPCzk1D
tD85WI7LhJPp2ZWFVeioSZ7EGjGJOcV0M7RjX+pDqd/ZY0PAOBGmuwyjAZV4Knf5l4wzUgY0G+UY
I1Yi1G70rF3RxDQMohIXd/cAiNPd/gFP5fblgdBDGM+FW7mbHVMS6cMdCVJc/J7HHP5PYYbBtDSX
QKrmmrMXh7ueAfas8XBySGwXAUiXRiyn0h48q2Dey3q39JPIyFY9K3ko1gjHSthtF7z3Gw2Anwh5
onUMSj0OudronwsQcqIw2hOx+SErOpOkH04xhKZWso3fT7ubRxrXLgwM4D8T5kYMlhrHNdFl8W5c
mA7fG1h3pD29057AjJjThHO6ZTI+19hSPVCIo2thrXca/SmFOF9/C75GxrhLph1mfoG3PceCBKw4
dAJmqYTy0m5fjqI6xJytgv2uFP8S2Rs1OBKrdB4s6SPQbr2uTEOwkwnZJEBCCCmMUlnZu0dVReId
wqOYOeS9aa80ZZOYRHEkQKgAy/CY6r3Lrn2vOQRivgdH+a6uSRS4nQOnC6rKthTDwD2juxCkbswQ
b7C/WChiq1vbHL89Go2udk029TqRA9I7BAu0I81oKrpRcKLSGP5bsIWcs67bpg3qcm3V7jeqjyvr
N8glgesJfPg5DZyUmhGnejO9PVtNJHCb1lPIbYbC49PqUStV8oOLRGgqoXwXyPz2xXRfd/0Oskee
UUwIXrv0zio8e9QnJIpRsroGLKFE25BVFK5nTHgHcFO+1D7ugN+/aRhUoY9BtANEySJpWGbTcYYm
vHdbsJ0cS78FJujffJw8v5LXyQAI1gxa8s6mutr7QgjINdSILLBDlud7xULwRREE5BitZCWDe2Lh
AhhOrdX5rEC2+hHqyxugGLAXfNxGPAUNY/MJWh/xYOqlnEAPY7v5lQN+/KeuZ8Gm44KRwlC20CS1
P6HEf6uYWXEDLQoGfapY2NpjE6vQS6aXf5a0pG4dlW35uvoKAIuuYTg247mWUx6Jk7b79gysYTIb
WRvcPWE4S2/Sf2MXYjfgki8/WbYaqVgCd9LxM0s4saiq9l8oAhWT8QwX4Is0v35M88TsgdGyhqU3
yQj2/e++VPxZqzHQ7elMST+L+CFatS8KYKFuOQzMusgj1CfssCZVW+O6XTMWpmJ7muJ5JxydO1gC
8RiPeRK3ShZKyamaTFVKnaQDIcdw9FAbr85eJok9q6CZn+mDb8Le2KA03e9tEkbwVZI0a4XwRmlc
5tf+UD9wIRsNSoFZzCZID/cgiKzolMh9e27tixYKmvo47rPwgqR0jBBxZ8/dcyOgWDqfTKKQfRyb
qNI8poAQL/iFd6QW9GCV3manUUnErJcpL5/80AZOX9YNACZXnKOKolMRN+FSjPZmHiq7V/1dMV03
hlowTcQCirsk7oGjyRe7N17pBRugpTTJqGNdUqgr2MgzEDGxclAkf6fieJY0jA3PIaKrrIyGEA1c
+BJGw9h7XGRrXpAQkvDXmkMsklpjkwtiXzzZe+2QF7O41f/soskkLahOwyCbbugebfx2n4Z8L+9k
OcTroQLzyic1duR3U5j5JSRAnFHqaPecb4YKJKILQZmkxyeAmRcCZvbwxdZ0cWyZTuZkxuXXEyum
jXyLaUN9c5rX83BH28QORudKSaD7Elidd6I6xR3KGL/owl70ESL0OYLMBUDmbPei/6l8HGGcqzD/
tL3iM/TvWqlCpTULutoheQhzedfOyaxfPc5mYAVc4U3qHHOEAKFttnUn5tL/yWRyoryrwcvMMGpw
jGXPI5nxrWg3Jxi54xgGa+nxz+X4D8B3Lee0kQIu/6pujxmzjsqYmt5H64zWo3oq8FhsrEeomxbu
DPMfslqWIwyqqTptCHjxMIAIpy+5A/zI2d0ov+vNincRwDgGYx3lziFHSbGXHY8iz4OCj34z6PfE
/DA9BRnlYN8liZVkfzLpK32kF7qlPoimktBq4LXY9v+6H5o0fv/NErmpAEgmdoB3FQm9fFmhKnAD
LuOjfuw5K7PkxSNEyFfRTySJqpKJCNBeBrdUI/lKczeImv3F0IONDut+jbVA4vdchTMWWVPhjgpQ
3oHSNvlrjts+wLi8KcMKuIHYUpj8jS5wluqLE0bcnO6ExaPF+8KkMlhbX4w5sR1k4Yd0fJv1rrKc
2WcrldepCMb3mFurC7huDiDeO6Nv6SrK5w93usLbvLv/q+DLE/VoqOFunrNEvJ9hI6U7IP+hsSVQ
GCxin3jwijFsqzvXxOJejSiQks1waNyKuiWePhehSAnN1RxMCAmBJN0BHmPLtW1ry9IH/sOamDp2
htvadeH09j0SWsp8XAucEMfcI/6G3rDi73dq7Ic+SrMpnv5fruBMDbWJA2pH4tObWAP+++ZCrk5l
AuH1ZcaK/aCnYTabbwrnhM42ybQhJy04EQJ484T7Oae7m9mveaYmXm5ub9d5LmvS+b1HJfwrh06T
XXR3jTTSPrnky9rB2RJVKn5TBsRlXTlQ9NnI4zewLLc+x/PSIg05T90uZs81WahueqV6R33f5lQa
rFznwSFRiPKX75dLAWFN7X5uXZwYwbPLayIGcRcGWNteWQAof3pdw3kxHYfWWy9nXKNfKxMcPd8o
iNYslmRA/F8ybXU8NW1+95SWvZbFW4+dH7LTCoQ3jpDmoKo8EluMjf6pZNeD9oPQvN1rJ7kFJ3H9
tWsx6YpY4sjYTwNJGag5c2OPew+UeVktIaaGEQw1/nS9kMCKlq0z5sM2UGFyVMO1Gy0rM8vlwqRv
QcheqL1aj4NjYCkdBdfgcC60CiXREFAVdghx1vPQCLA/63hmzd0zVgZeilquFsqQvs4jMRhVPnCH
auhP99j5yWp9XWwbd6u9Ol9MG6lk8lyWcmVjK1leGcuL4UzBFH5eeF9buTXAL0TFBehokUbY/Wem
K4QfSTGrqBsw0T2Ohuuy+ykLAxIEtF9JnZqSIGNdwBhY6LlHI6islxhi11Vl9V4AP+TIpfOwgGZ7
K6/61c4Udxpx+CQEL+/XBM+Gl4ovC8yfmMESQIEs+jqvaY3zMfx2EV+xpRVnkx+dpSwvQaDBL/vO
1doJdUZe34OFci0LkCPrTgoL747cWMvpKYR7H2xvTvgSMMN34Yv/fV3e60Rpad9sbtAnQZ5r04S4
eZs6lIWJXSlahtgcf69YqHLXqj6/9bZ9fSzq5bVIbcTSeQ3W4i69zookIIRoJ4Bp7UQDIWPXULkI
Xk0IjV3XfM2IEWsX3iqVjSMz/E3IOnvPLmJfnYXAfeCsy6XQtFN6K5F7E6+5c/h+U5Qo8crltYBm
Eu3lRRMHqWx2sGA26BNqFIT30hCOx9b2PmoykoEI5pscuCQwCn7CcADgIwu0/NlFg8I7dxN48k2R
6bEx8VYkBrqE2bMiWezYuCr9u/Q/hEFIcPi6+d1DRiIY8WGTemKJ0JJTGHvEbW/PsY7YiaEuTifX
wsJX2jwSLGPakKbiV4NNrn2tpfsK2R+UefBDBtbuMq4diHJVj3/TYzJq8z/cy+91cWVnWj7eVG2/
O753HJwlWXl0rLmC9HMA2+tJxkwctEw97czevDCL2fipy7GRNWbA0iuNAp8CW8gVGucOG3OYCVVy
5UnCcijDVfawLBNaWXbu/mz6PzCR2w7rPswsXx8Y9vk1OKUKMJXc4M93P2HGg7S2rTDYniawo3NZ
ebXyPTz6XU6lNk/Yy+FUliJsGCFZp8KoPp6yzgBcs0kmQ3PaoKbkYB8oW8CtHHoIIDQWW69ysu+m
iEMjrcBRWxIgCI3h9GLPwTyNNaqMS49YPEx+MAMPhgmORbOHVxL5lTXI+mQOl8O2GC1Q9nsoF5QB
XPOaNll3KtbCVIBJUrPN2bR3cDPRCCCV3rL6SZV3VWrGEdt+92H/UL4Sv3Ov4Y54wsYZv/tGFOy5
8VLAAkLBCoTlzkijFkG5YpXBeAWs59YhTSl9DDbLptWTNtK/yBAe94OSUlZ1ND30p17NUhB0vruj
NC2EmN0uJBz0aJB19vZ0b4Z/PrYjubnKv+8nncaZGWVRWtYQ8zWZ4I2gI6SVOeK5Rk2J91KsQXoT
d0sCRBxsZ+LmBZBAtgQ362WSz2s4X0IXKjhNQVgbrNapfA+w7p0oEkvbWxC5mCis+GvkChlqMAU5
3ySH8AMz+LJon0rpuRfWUP4N+TP2vySdKIsUHnTJOEmTOR4dSTBM9IZqoGCSKIwzGMGOGYzNx/VC
01Bjc1ZXu3fsjCNS8KyVSbD0v+HSDi6zHqgTaEeMvdHnD6gkNnDKih/lozVyKUiL7iOzfWVToB+8
RSwwmEj44F+GSKbehJzScT/DMnQx3PeHeDWfzN/COoZXOH/drXfambFFe6bIfSiuL8d/DR2+amNA
b8aGsvFpgPEcqv/YtkUjWh8J8LmbrljjLG9qRp8L14T47eKmvDmIj0C0AcPd13ihOokFvxvX3HZf
vYwp0g7Sbz49MsdVImOkNC4HWkunvuV8drq4AdllqEHUIb6Yq27V03q5AGEbDsW/0YQcG3BFFDCj
5klvCea5up4mpq1CpDQmceSQZGzO2P3hT1hRH3Ej90Nk7eYbvw6nmjuJVarG8bynAB//asHR71Oi
wBSecpTa+k1MB0eZlP8bK1WkFI6+dO4BJ2Wpvz/+VfzmTQpjD1QSTMKKevCRy5wBpNBBvxKXC8LF
3qCNAFktZiCNeRhhLXZfsKCTeebHESGFE2EK0ScmupTmpZNegqqF3ckU795O6BHzxE0M3YWuJej0
FLu4lsvZ1wby281of+S6cpszjiqZy9LiVuocpc+H025IGR5wINmzfLmkz5kbnD+xpazRIS1P7eLV
5zvI/6u/+ZJ9qNGIMcJnv7PvZ9lPPRjpjNUCqiLM7FNK0wBlUCZ8jMwMTPEGIZfUNvGzEETRYJTW
JyvarCZpC8n3cp7qljPVp70xekwk8HR79eG2pxF16vnCIDJnvxtjrOzW16uupXG/oHdRhR7Eso9X
lujHjwTiopxlCQhUkoH32/cDsJKwAinAEnrPSAfTw85LvE4F9TmiLJWjtxasCx738p+ildLHwMOc
Aum+9jQtc183HIBGAVZ70XjkIYF9qJPrPUq1jj8XLpHVVJjwIZFKsIVsMh80FLAtKTpcBeirw5RL
GVqz/okdeYdAFzxWHDDfUCIHh39kBTJ1MHh43LDrw/8KaxMYES0w7AzpzN+qC95p21/0yNC+xOEg
kGrWQEmcxrdxeFAID3ROswm8CwneOenKCBohAZWTDpMpJtjbuecveslGDUO1aHWKQda/ya5VtaU7
L8y5PC/Aqj7xv7Po9bgeAXzqkNGHs7538uKm7JLyE7anCX3U/tdWyKLkyYdNT3eWReIk6hH8KkC/
RGAol+H2MGyfOYWCGOGmxPCbyBJSJMMQrlmRR5zMuRcxrxNZqo9DR5YkVsULaI1asYbSxbOKFHsH
x9jAuWGfZ4tyQIYUrAUUmthAdd2NXbMBnxW+oideEPgPLNuD/bFf0lxTQFgXV0FXePUNkGSlR8fB
bPFuODD32/5ygUoZl4v6fM3o25UYQbvyG/26XA68Vj3laKsx8o5A3CsIpPYCEIkRikzftBN0Qzb0
4ksv39suEG3+oowI40BzUZSfKPIAXCJK280eKr7sINWocmMX/UDlb0V3RT8VoW6/ye9aSGld5HHp
0abf/Cm7JD2pp9g3rgTPhPQEHwcemGMu3iecztkA/vwkI/V1Vl91QoNBs+cCXBot6BDRb//dQRe+
paGjYqT8eDgGMEfLE3X0cMOAGjsuRbgZpNQJGwamSAeFoem5bQb9byW+ZpVoxA7VoGYbsA/QPCvp
b4/lx7QwNLZIoApd7eiwVOLjmAIKjdYeCLEmHZq9TN9CPy6acEgHGExUfAqu4izo2F48HS7o5BkS
vFl+bNZmyA2SMkZ1xXBg+Y+fJElWbrd7dMTArDIS7iNo0bjxB0wsT/GVow5uJcMTaM2CQSiOPxC8
q8kHkpIOYV5BgTRhJoldxEtDHxn7j+6JhEMn8hMkQilJ9YHc40Lq5tOnCP0aQk1SVQx9tzTAdlo1
HHnwu315Cvs+JuxvNuMPzKaMZ9KkXYOsE0/k42i3e5ie9zXZx2dhCyBfsrdOi3GUupwG5SzylQPI
TKbJB3rSahnNV+rRCcNMEnq1h76sJ/SoM3wzTiuPh2FRJQl6xswo+rIlu6rYsRJO0edYopNc/fSK
2Ul1JzbJet/tvMXXlCOrwUOgHUsEmA4jmW+VTwjt5u0S7QP4AeTURaRlaLmUrOq5Gl52+Htm1p4w
WMD3GhbMPHU1+GhhgZFw4iK73TIC8OnWVVHZQcVgNJFq/veqDkSXHv7NIWXsyYm7EPRrLS9Shaui
pXNNCneabMNq6RgecFI8mxkqkIZ2n4HuYz/KN1EfOPkNcgEUiauCapRI2sW8gqGsMjz+M7prAfc1
foByizK20VRSylXUDGIsU/3Y7IphWkIyO8g9ZhAaSe8YgqvbnYMyB2u2GKQwWCkdPUwxuFGob9AX
sSyF8pg4Ipj1lJ1slBt3ty5oaE/Fi8TNdc4IiwtZWWDoryxqSVfl3OYjhvUAajgx4/yqu0JK0p1z
hPqz0+/+OHruk9+IyqwjQf6CK+fK/c1hdvgvY249u4p7w+Y/6UaHzfb8+O/TbFr1QTTNeyWp3rc0
A9E4LnS/+8ty4BS633s2EBVImO0aq+xul5R5EijUGacRRMNxRBlg7L1JOvnuJOQ13JRi7peTpNXG
89sAyVjJvw3hDeWBCm8ib+HZW6YNg4GYOoS3KOnY/DDzDc3iVwpRvbVmKcBbwWffncpy4dtdlRps
+RrS7rCF9fMvIvUneGy77y2tm0lhDQF6VEk3vUS56rWgfbdQwIUyIjWhn80U2DoUpyhjpWLIOAdo
MbIdIzj/xJbaLLL9cN3p966lXML4xGWaOVBHHfoRXKwS6XjSg+1vBAAfuPtEvsOfR+AGFcZn7dRg
4VZ7B1gSdlxS8XdtIu0e6au9fLwUcHQgrvL52lKfHkbSvz3IDtD2FAF11dy70nVt4stvsEHV8FqC
u0kKdWZS1s9ODQYsVeX9S3/PTPEB6E0XrrF2EAimQzmr+V0NDxeW0/kgNrR40+2MhABGly9ErDci
Y8qvpfs9C5HSZ27mPtgBnhHC5xL5rLFjJd4mnT1XAROwEv8A7er7SeNHMremoxsDbmr8p/NI3NGf
vhlXNI+SrMhMbQjXml3bY6w9ac1hSbIycBRqeKA0x9882S0K7xP4AGXCSX//7L9tRntMlh6ENEQd
Cq83pV02LV7CISwjsfViqJNORUnSmU5kj+vhRP7ZJ+WwTxZE9XUo+Eu+puSTgPzMW5tstzmZ5p3q
MhLj2CotN1rGUDrF/d19s3KPZm8CW/zRQMN8t7ig9/MVBWliKbzo7ZXKs6bbcG3kzG++8fuqAwWR
fHtvIuwrOu03pxfbar274VzxKJtR0MZV/w3OhSoUsBKw/40R8PDLLBBn1v6dYWBhqHq309Br6vI0
qO0+PijFo5uxHloJBdXPq5T9ik7IdayRRRqt9RkT+dfXP0rOXilfX8SIzQvXSuvjGsUCkorTDWiz
0m4zh/wiZ+123JKPR5uCxmrkk0CiTCR6G606E5shhWX3DPXIsjeV4rKq8IcdG7OVsRlaalrOFV43
+u/PYw40naCyvkYiGDuz/6vBjHK57PeVlXTT+OvJG/PNfETPXVbggVCaNmgvV27mkF9X7srerPxn
AIM0G6JxM5adxx/HpH4BtUU3SXg4KNFygVaZ0owHa96LPuvWudrwCZWgH72fYgoi4/7DwUF7Z3Y4
3KzreiVKinsfRFqeX4oViJB4JOHFWvmcjArv3JnaMc3eNZHftPMNwcBGv+hvyjZ81GS584BtJUVW
OkD2lt2SL2vo5g4rEmLp/pGpaGtLPxqt1V3lRkW/kie3yN412xIymfeC5ngKeI+h834tS9gALCXV
8Spb2nORiAevM5P01qVYdmaMvEDLARGEZL1NLeTJfmzbux3exNlJnf4CZJLn8mmoOf7ogZM4Dmfg
QFQLYrrSvLdIwOYxJMkAMtJ8qFOXKdyjMAC0l/H9DjRDqDXV8mHy6P1OmpLUDGryybkeDVjblPV9
z13oSqXOj1VRsLtyNRovTlsgV9Q0L5aN06TabfiJE4dshYJXB3pvrYHnqhnvAUmXfRjqR1r7fdm5
birWfxYCxQ7QrhZg95uIx7vonhgTZmObkBx7CKHCLwMaVGLF/DHeyvxpBPwBgIvxiOarJAUgb6wy
NzWcxOftR4OoGBDU1QB0BWsCohE7xRNvvhulIl54mCyNEV2B5insO0HeMR6ysLGgd22CSCbztxIc
wQhSaRKz+er4nFa6nEDYNu2JHs7SpxJH9Xxx+pr/Oo7fPTyQbgfl8EwgQmC8blffD81JgteeBsQd
yks94cmOyNgVnLhaSQPe3ZjuTiJ8yh7SVqrfToq3ixp10O4LiLSAUyc3HEKXJneiBrWgoEXtNc28
lKAee3WmxV/DO/AH37/VpfkstG5tQSz5EPWnlz4MXklqMmE71B9hYDtWsU8e7LgOcbaGHbjXXxD8
Ngmty2FA83p1JmJhojRr0Rhnb+9tJudweQ4m3hSF8R9M7g2GPqMVLXADPxvV+u8E85MlF3g3OcDs
XWLobanXH6wfuKbkE4YxkXNXu4mDmO9V8wg+DrYJuO07DB8793MKaA1v7nSB1I9ZVgPYlPEoDBe5
k25hbqpvd15AzWVjlst1D3GWXNwmiuL7lJ8SkKhU4uRVlzW8/r8cZeSMzGh1IL1qgnKMd3s6d15l
3e3YPD73x66dqZ+r9bAWPZBskxMgrq4u43LMRiDXkAOfYcjhilVU1CR+W6jPPWvpuc3fZcQavovd
d8AJe4+ny+UMIxsfkikRkLw4dSI+NYoIPNY5aFviYLrZTu/GVDNmh3p17pV8nwBtRBLVGHA5+MVM
Ho/zd2IhVQDxt/GUSLW3Exsunuwqo8pFBu8q2B6fOjA8zLP3/Md6vh9OwvzB40Gg4EHGucE116+U
DKeu8H4MllaCuwM1c+T/rygdsTwTw/bJg5tHyvOXfbAbfYTjXhlqTlRVZ4avcpOFx65e62WfzMnP
xAg66yx2uC7XbYGcRgjAlbCAyQNOs2qpKuoxDgVc01f4FRW395P6YMaK++GUgM8CCabKRI9231Fz
rMDG/a5zABYj1u94qFaC4LQWb/dBXdDzmqxerp7v+gjfhPzypyy/QP9K9oKk+2ZrN61bjeIw2iyN
GBIZNRyEYHIHG6Ql98aN0YSDr8ulv1z6AgPwkPB0PWcckQJ+vFn1vqn2uvbtEfiyvpaG59il/3Hb
2dTTXPM+6/P67DQW0LlSXzhn/BKDvTOlccdOSl7q6oQ5k+s/lPRBgS5pVeIUx2TkXIeINsEFp/f7
9Vkf4xOUnkXYiLWOwKt8Ofw8eiTcyn/meTD5xt9ozw9RxiM1hdalOCunCo5QDqA1GPPhyMvGmMrk
YR5HcfEUmN8ayzasSXWauMrylJAtvuuceYmrI6H18o2yM/nQKZ883yymuSInkrQLHS9xXwXLL1zo
8iGJVsskmw71pHLtyztRGOBBcJ32qHc+fQcy9xtlxabvFi6+03fJDqulUSQPWeP1d5sQWpO4x8Q7
+6mFS3UzY1Ot8a032djm3ny3GMZZE/krFrTey08H0146OSjRDiAPGkf779pmk2bP3PLCboEiyXbG
8NO1YEQs2JAilES4uut+S+t5qUjAnTp0uusmSIwAERprwfMxlJ4yEBRuj3vT2zP5d8NX2LXeT6qk
QrwpGEkC/5PiyMi5kcoi8qatzIM+o0Ubz4l84WixWTTGIXM2HCH3bnmCoGNsesbBtYQwrfGowUV1
N/dLvbuIEJNDz3xUywGc6YzQStPvon1xYFjvRoGOxMMizBNNV6lYzg3jqR2W0gCcZppvwmLfKsJK
6pKEpc8uP3+K7xl0aynUw/h11Cf+cz4wKBKcjvcUQ7myPH+vkogm2tt/ZFs0+GjCRRo0qabpm2A/
29Dl2mGCy6VXJgbG76iuqFw9qnQivBjPx/ZJAhMN92I1A0rWY/nh0G/z2OUrR71SmUqU2HQC3e1c
Y75R8IyW1Coti2BuyROQXNGO4x1LjNEMCqxkoYRdMeAQ1+vrTlEgXqMwXj8muy6dRRZx1D95o3FA
LlmsCDs7h9qbgTb/yYkNXMJyXhAteEcsNxuryIMp0qonkNgCbt06sKOnFMKcBcwdww2FDydG63hZ
iv53jAPocj3tmISX4UYZouR2OcjvFJXfYvUzC9S8JnooCEtZFyIx0tfVDOJqT3gtkkqFIABnZT5a
C2A/D8EtJ1uGQRiUDBFGu6WoDcyG7UcsV69jsA7p2DD274bgRKKViZlfT616yWosENp/Vze5WpnW
uQfl6UIg05wgSALWMaMsBrnKMnXKFyfBduAlE8jPslJxzHwLP10IV9Kf453wdOjSnfiy5+EbRf2t
wQrCyMc8egL0lEHokDKQToVK3LaFeYLrBlOhDzjCxxcOxkG4N0zK79nmQTyGYUFsN7bZw8YkkcuD
SA7rFGA3y9Q67LbqKZ7uiM/smmGfSuqnE6kUABQRCOvEMTemsWIQIycIkXrlwVx6sfmkynibFMyu
jCU79Uc2ckVI6QcO4e5ub7DrTCp28z54DT/W9iaSACY/YoTDKsNgzKnJOF/iCdOYoOtgAlNPp0pM
24O1i7oRt3nZYIJ7z/9/vP6aGs1F3LbZZASiFNdtEJ9XcjLU9eT2qIRwA1smvDK8T9t97IjQkrJ2
dr6FLJ5/xDvJnNirojmAworJ16uUaHmWou6tjlRjiUbgQghr9ZKqayJjsoaKdKpiJjO4gqT+tJKb
g/llxn5ZRrXCFVayAojVhWPqnFgyRrrbxzaafMzMlRfcFzZUInHHvFZCOk3cVdPOu3ZFVldxu46/
ac/nNCqWgdcAeuCbGFnwdgQQz+0Pg4BeexMNF7Ro2WesS6xNRvWSsohCVYrMqpo7zCrseGeQiIDb
NzBuF8CLQYd5aY4AJqQoxvZtXsDb2tlJoC22TFRY3nYo4sNP0kuroLReXUVjgzsA503V1FXHAvYl
04/O4MfEshPdOpZ5xj+H30nP6VJ2xFe0uUYPlpSZ32Lx10Uf66ne7xiOd/kyPPSZFrXOa6LfGGWa
2Sc2GtwPRNPHYC/o8PkOg18MeGzPA28ntRmMa2zVR1WdLm4QbW6UkJPZnJYuXNZG6uTXCC2sGwrm
hXLFY1Hvmg6hPnUmjWp7/bNgd2jJU9H6+QJxe00gE85dGbvJVTTVztSKYrSnrukjyuIE5WF4K99j
a/cWoj83Urb6pPOpY091bY0XE1oHDpdbYmDUBPgm7nNCEKkmrtYQNnttFURZJ4qj/7LfI1vEczLH
DCUfh5qFnnjzwRVXlhpSC48e9F9Twj8s0/2XE7H+I2t3GhSuYL410/H2rGZktsP+EpHb8tUpUdf8
sV0m1wf1Q/qnRcvo3dxOASgmj9EUxjlxImybaPxeOS3VLii3l6CtFS8NTO51lQx+HnBWVwLmVAct
F2X5+n2cGDJDDrsTUYTpXWebYF12V1ZMC328vUBAJ1J2bxh7EPdnzPZ+3gw30mcxCHvVxORDQnif
wHfP/2w3IFGUMF/dO1LVpigI9x6nDjaVDzNuCqkgav5cdSF1BV9XdD1U21xQCBS4AkLEQv56+pSU
nfbAF8o9Fy1Y/quakFJwEDrw2LMiba4znXRXFBrRAMCG076cl6fybnrnjaAKoBrl1lvCDWhCs6fZ
dOq/CRP7EBCg+1kxoHCILryy3f52pjR+KC+MuiDbMiMDVCfLI6hom8iu7PU2fCvyVvZAg0TCi4Mi
h0LdOoW4RqV8nopr9HNJ8UdRIUnoQyJanmeQtBdGM3unxl58yqnfnKY5WghKFSbPTpwuujDZ6Yce
pliS6XXnfgMhocO9Y1oJ7xtQVWbZ4YOPC61aJ5PzzXp1vnKriEI0+ut3RWRs+qF4Qk+HpPFQrKCX
euONpnD0wH7ipMUtWHy6G1sZLwMi7vnjtx7Y01ySXE/sPTMJB6Byq+eFREc/kILwELTSRnWK5fer
/EqNEfMqu7HKXh7/BaHdCK7sgRNSwSKJvzCTwRUSF+NtmD4GPR9d8Tbj9uYQK30UZ6PGVfHCtSm7
d8rAXHjPz2jKf1SUonnWf/Coej4HWr1oxIx6rRIrqg82iyZ7VLW+ecHybdNHBUkMuwQt+P5CSlrN
4xAC1l83FzmVTDD16JTg02/cKA1tN1iUWieT+NrxiL0RIcCKPrN6hiIOdhGawsdJXYjheQlfTs4M
cuBHJXFgY9VKMdBtl0z37bVIvTL7AqaJVmI5HTFDUp3nZ3NzsoxTj5ebXqjdpA07on0wBCcReci+
bodGT1vJGaiPoJJeleW1UKNg0Gavf6Q5MdSzl5Ae1ppvnknByeHKQJSVnyFTkY7/y9yJPtiifSZR
5bVOxqL78nysIKY2a349pguIaTNOMdE2h9ssIAZxFj+jURAT1SHOLQCYc5coxm85mfoCcdS8LSdU
c3PjgSfwRA5aonhRF9OYimjpURiuwnFZ21+Re6M0j5gfIlZT/RWF9FnYXZvSpyhBbHdVn+HemvNp
9icLHI5JLFER4mYsDS6ekxXx14nwPefUT69cEHEe9E/zccnMwF9+6qGYD0Dl5/k6anxwAn35Ikda
6BE+68zvVxRY3RhCbYmrDj5aGALut6BwZCupHFXEi/WjT/PksL63PL0r1B6pkfjEJCYJ1wwR2MKS
OYMWiaWBbmCQ/RmLUU35AhsQqHxzGxsAyFwVDrAewPvRJhdZTmxbcmKFIe4hS7PUFmdlOldyxMkz
CnRuD0zs66PB2PZBp97T5ZUXI7hLbseRMLGL/r1ORL/hbMeY6i8Nk93HqRM4WCSlDowVmK2PVd1K
Jxsah2+vfl5bCLZ/9wSnqtLLVl3i5UPXbGmNdII6UlQ2qmXCq7Pyxt1SCzE6Vcc007vIMTZgJ75Z
hYpKlZFdNsPZSXLaZ+gyQu5W/Pjb7y3adUHERoXc4Esw2M7SFkXhboRPEMbe1PWmyBJ79ep6ySRS
cUbmnc6JPN4x3Woapo0Zt0HdGQ8+L1qYh2mXtIQaXMvVltGkl6wVyCMHnYKNfEvfALNn6YBws1SO
UoBEGswTvSKJfJBcheh00Qm9sLTI7T/PMFrrBgcrsegJ5uA6aFkTt03RXy67tNmFaIr4z7XuqKRN
gLjnMl4mTdJtpiqwibrteWH6AZGT1Pchj2lKB9QN/0ghICRvutAJJqaRKLs0TLhZT8456oMDitZG
Pz3wVFpIDK2UZbzHvDahTcntfIKGoDQuVgf6An+ZKNJPJX0TyOX+l3Ve4U5oKMZ6DRtWr3FNq9oH
YR9dCH0chdkKuvSkp16XYCGJu5wk6QjuS+xKZNw+OClX49jAfrl7LzGtnTsbFe/e6R6d3KfhLLdi
DCas/8PueDOT27M/BqTx6pnVDF5cbGSacEYLsB1Gz1ZrUbSkz3d+Gb4CdgVgz4FJvClezBTiIKM/
hqmdJxRGZsQD0eQ3OvOGLsn7UNrrb4maVTkurxp3OWMv1eGf8Lv6uCtuvHZWsBJYlHyXiIlNkTit
5+7RNI1p01iL3qrexMkwzgcxba/bYDPaRkh1VsXP9f9Rs7N/LRd7M40dZBF9QfBLX6R9NnamwJIl
q9QaEQzu6v7CbDsUu/RfRey76QiM02D2za1Ne0CScwcMWMCgQLzRqRPy7fGh6k3gPRMR63OFb9au
WggguuyjbJATTJt2tKSoLpmTplD1As7RNbtsvankoKFACdNqJJQyQU8iknXe/ERE0hAOKfjUwQiq
xDUFPWelkRtUaheA6rsPJFlSkwUJ9tyE+CgOCiyEB1CD54IscsIgfgXo0L9tQ6duBudg0TGx9l8G
ahZSP/dOfJZqCnBRlFCaso5Vh7uA1z2H4MJZ3i6jp5ZRQb+ze47VhZ4pKbaGDk+hbKDsbtJ/DqRj
Ws5XVaccHFAxp7jC6BhUresykJNJZPtkUX/ZyIZ61aNqLAXHG0P53wjroOE4IZHQ39H5QKJbR1oy
ht7332dn80BH3JF5EBtRDJMEcZ3xMw5ecdj/UkljjTZ1ndjnY1SzPmxKz5C58vsd5G/3DuMpwAKP
Vd/w+QSTDvgIAMG7G6+V4KI05BZ+DBXlKBaF14Nfvf8CBNNTLoUFXrnCTZu3fbyzrc1G61FIc+q5
eKcTXU8VC6G+hXFsPAIvm24ZRYk7+HpW8JdicdzSPZB38b4plN2Nfx3LEZSQ/RW/OewHetbLFHz8
eYsr+ghgdNO1ueAvMouUJ3UgeCB2SdwLXWx7XDumA4NqQqL36Rg21BU+k557n+UuQ7XgqFQQAbmG
pUTnXxhvkvgej47+wVv7cbmfiiTlUzH3+7RAxImB9Rvrc/tGirYnGFBGYa1zravov2LHjoX9M4/v
yBI+jHuqWXwndIAna3FBIZ4Fek1wPZiEyMHvY10zuJ387eMRRPs8SwA28Gig5DDhUERczHXL5Ju0
r/XbRa4JfplFmtfVHV91MWb1SHOHcwOTkz0jjBx0TvgoElcIv/ftdTof5ISqVzA7mktZt4xPP6zH
AcW91RRJsj2g47B46XlVFFCAlKWU8xDfozkJalrZ5Dh9hr2WCyJz0fQf2H03BUv4iA1ka2vtxF66
1t59IMJZ8mcEgDANeRbZp1E2W1CzXDVcvBy+/wMgYmy/m5wCgB1L2HwTFOwSGfKnyFTUF5Atj0p1
3MRLZvlI0zU26W8xUp0it0p120t/Kv3P6tCp5PvQPUcLGnSY3JhuJyM6CaEuBsqnbOGYRegb0pDQ
21mW03grduEtORYs0LNe4sLNtRkgLCBT9rMjz5P1JH847b+byrTnGFiMCNw6Ea0gF7Lham82fvk0
DuJAIP1JT8XjHvjYwCo3hgPdJZnsXFsnzeuNNyxM+P3/CUeQMZDor0Ut2QBeelRCswhXa4CC/ARt
Cd4iXgAGHzmpN3o8DuHaymXgL49K2FlgqpTuVWZRkHRVwqt+jycsiZBqj0mzXX6EhfZbExYwzsFW
8e+GNDBr+xHWVWOsstuKX/zLrlLt5VAcH4T6lWweM/NtV7CVc6zK/2LOb5grgRc0uGjkVvDRDfYm
22vkqj2VSg6IPa9eRrOB1mGQxodxSF0ccf+p7QwP+NBxlD6C2yUQP1L10Au3DzaziqOKluT7ycUJ
JxUVyMDlopzGSI7ADe0BMm7oE6zdSQUqJNwnymxDMuC6o+MvhSyEXV5M2nwbBW017pf9/rGjAf1c
O3bO4GYzORR03ufH+O2on5QqXKCyjkzQWtyKABLUIt666gk/NLChqmhoQinG+6UeP9gN56rcUWhP
iGBBr3heGfBi4NjVAYQyIO5BbAqHqp7B2lREbNEqz9sTjLs1bUWGSkhr6mvT0G4SJqjgg7zQkLhG
NOy1edSt9t67Gy1yxAUguUoowup3011tHkmNXxFtlVyCc+zCeaTj1F+jWcHZhZPRpxC5jPtBQKf0
ZN0Zm5lpcxXt8rLpWh4FNsOVpJUsXoNpY3SyfFSmiUxrqw5JZj5b+sqyh+KgRBh3VA1tpNLY22E1
jZvv9wZ0xUrYumhtCT/XCgx0wS3hCNiwDu2AsZfyaEcqcaRxqh2ioqKWf8vEs8UejEDrCOY3k7QM
yMCRfqGoEMltGnicoHA5mErd5ETe9P8uGT5lvP7BeDvWStoozCln5fKEKPje1crEbIjfXP1WU+Lm
QeuhBIwSi+BXLjxp2kxELBaMpRlzH1GYpHKh/8p2iALFoXW1s9SBD5EtE0d+xFHp4cilBZjN2Izq
RgaJDknAnzinvsFOwAZvbjI2LN5VT1WMoXRo5T6x/dic40HPlb2wsmpd1gAYLUxgdE6iSLGdhWLR
rc2cV4YolOc50Ag9aIzKgqy4+OpQ6trPYSsOk66TJgPeVQ0u1r5WFHsSnmpbSnXsp1rJMXNPIolz
RYmmaNp41LUFowagkCpL7zEqRVGzQ4luU0QTl9fJCV15zPk1Q1JE/bR0lavCna0XzZVVtCFsEj1J
C82R8zc0XnWMQ7bnkmbY7V6z0w92k1Q8UNVq5g4/igTs+HGPaPLaonr4svoPiN6YsKuA5QhABQ0/
oc4/vcBl6SPvSmiEUwbCC1E1uEx0wjhFkSBdOxNbjME/O4d4Yzyn1iYTn/0aewAMyMxrrCfFqYXk
TSVhZXv4yq4atISmRlNbZKczsNmc3xHCv8czZPnEIU/htOFe081KSg3FHh/P/bhJMOhkZ3c6COGT
9Al7ONLqx2aVt58dlYTNEbciPsP7lhm4kfYSL0olPR2tTo4Uq6HaNvKs6LZqWj07tXsSG/4QdwrY
LSFVq7Tj6pDu4GfRYwoJ1pF+jS18kX6gfRzjODfpevetf6Ni4RTAC2WcnsGA4tPiAruz9eOd9lRD
Rr3cDyHvW/mpPH1gW96uezCLoTz71LW0xJkFz0b7MtFg7v8vFUxi2I2O+N7Zq5s9ZUNVBQ1u7+5C
FyeyM0TorF6W4WGVjNJ9jkfq0zbuUam3Igj5jUdO7tStG/zVaqhCniG3gLys/KubfEXRXgGXzjJs
ElrPgr6Ye5z5Q0mAPjT2NlV07vrc+KVw4LqsSzKcOEsCUptHJocsRDw+5IMIJVYfRYIkNfV4/blz
25QKUQLLHX1d8CJWSqISQ6BI7eo1eyB77L1YgZPefD2ifJBuJC0jGy9ikNN+v23d5h7ajTRjz7It
4wzsh2v/FdTQuJ4YkLvxK8hnLelCdc8IlSk1ulAglTSZmLSMThyMr+4XGYYfkjSlRN8hlXbiUyll
t47MT+M5/x1mKM7TpIaOuc5Wu2aYCfc3sGkbMWaWzZ2KdK+6r3K3N/MOn9o0p0/rEA6Iglo3R/Cq
J7o46trd3N5s6o/MzaDslgFQV30uX4Njw09zXeXa1pqJHHzRbAxMKumv0C+En4U43NKKz4lQuovm
Cm5vspUW51c+jgV5BH9aY6bJCJxiBb9Ta+jYF7uFcxsfQ68Ut1/mirxq8ZGrm/CL6AsORJ28paZZ
7uhHMB/GsT32WJcwe7uokrcNgD5BNzH7JMceYa3zTWY4g9q3r0i103c6w7S7bDpwCgIyzNvlIvec
su8UQTu6ERsdRO/V0Af7+T26/RTkYkE3lP3HLnSLxKFAGQxnSfCMsuY1rfqnXFkn9eIMzos2rUo4
K5zTjFsfPUHQC6QHsKJzYksnKmmhdAiza/VbmTRuTGnj5xiggaIGEAMq3QUISUm+Wmn9vMT0PDBv
QZuzj30ArQCqKFHK6s308q96CJ3MqQO0pEiZ7rCrUNkXCCwxlarh6u0Att5cUozpbfjHWB0L4RQt
bTHabk2jyzUNSkgq5KK9988J2fDmMBx9ZqpWZ+3tB2l3SxpYJhwbXupAWewRLy+ISr0LuY8wYbsW
BNjn+tbb3y3ksTqcD+pJNCaOFBan+WBtWjtl7svpRWl37KUPuctLXr5iD+M9ikbOnIYqmyOs5Hwz
KtXnMmACHVbyb6QP/zLzO9zz7IrNYnXakz1HnVn6wxYNtfVbVFVlNsU7YAXIr868Z8TayLPFBT48
W/S0Tl5OImpr0VrgmWhRCuBqMlhM7jNKfKgE2ugq6/SVcOL2LZUO0quHoNq+8HDUv2gJ0nBQVP7f
wEWYKb4jEFJZ6vA4R6afQTwD2vZL/0xuLwa9iu9feKuEseoEjIivN4NWTS3y8vxPnm1BdPF2tjX0
3oSoYZPv8vViDdlTpiMLg0hl24bOtUxBKQEgnGXBopHuDzkmagdi3GVh5o5UkOYoKITgGzhnnNM+
OGOyFi25l1QpJa1P/N9WikbxlHKAYtNnBcpFtjPH55SJP87CF2kiu/L/tUjagVtlA5gzMoJYtHWk
u4NhSdmgVE2GL03yoknH93r4PpVL7o4ZkW8UYAjuRFfhuaS75IZ7zMDJmGG++SJEv2F7E8CadgJe
5LyWDVW1MuE2nQIwsdVl+qIcSs0dZ6I7WbMPEyt7s64qgLWjLWiwpEmYVfaWBJfN4UuQ1WiDJS+q
hMxW3cUbhesQAKSZiydDWfmK1fNyK120WxsAEuxTo0s0o4PC+rzAfunb41rP5V3AYWVRCxqfSFV7
UeTpaXV9h3OzKMXx/nkbfXe0SBpThx96ar9FrB23GDEFN9Vq6qOrC3rh4KtrLlfqnCecMeOg+vy0
GDDYjkp6vSaGfgQ7jKZmt0HGRFGPCFIFiZSU6udS8Q5JyFxNBX8i9VFAFHCUxkqMc+2r6Ly+hRHQ
Mx2X2DmD8x8Dz5rRJ8+Ii3ZkZRQMeSGeL6aunHXdUKgcesZa/2qmgmzlM5M8t56kZOWUgNTf5eZ+
ylvpbfjGGUC2YgZ+lw3Q+ddQj5F6lIR4Xx3x1sK2ilSAedNIQm+S2mnoQdCcVf6GPsayfDS5C8Ph
GLm56zTsbmaiaBgnFbIeatKxOGpRR2EuH2XloeQWWF87g5whJ8p4xTOULwA/ezaGyzWvYpEA5HDg
IRIj7ljjTw4/CjGW5KgNp6SDGyizYZYjv5fdqkBahIBKLMC83izwttkij/fTvliBEZkhnycEpyeY
Jozgt9HCXQvMRI56kxf3l8AtWVIYgeHVZGpIKBLdL/Zd3EUoX4oxsN8gcLG3KlXthFTqx0jco9kc
43QPYTAntpPygSPNgdCqKmfxk2pZ67ZRUKAoNIS+wSHNK4LkHEA9YUZtEQAeDhgulwngI1Um+ZKp
MvyGzHZcePVFD0DDVfQxwjpyHqeoobRc4wOHas1lqpw/eFes6RII9+oOOtcDWDWRaAzf9VIbR9P1
c0fOSW2NwWJf890KGfUBWKLFHqUJUlFrdLW6aVI2aweEiBp7Pmm5yUQ/8XyDvbNdDm6vwvgmmAOt
yEZev+07xcGjaLR3p6SewWoBMsRX/lvRa62PRrEjJFI8xo6YT3Pm71iMp/M0F2KLy8sYafhbhY9O
aEiroA190ASD2E5yi80cXy3gS2esaqTShQzzUxCvgW/ZaFdU1WYW2ql/k1Ehs32I55gKJ8IQo0rV
N/XXV2pWlRhVPDJggEgPASuwpII65rzqCdvBkJuKjdmW5G9TlA2aw/kGd1xnYOvizV92x/NDeE8S
9+XMh3PoBq9vySBxte1kffIqArhPW7XvTNac3yjm7QTTCJVdYFOl8eTSXXLaYVDXarMb4qanotdT
ylBX051XZ9/6TJs7wufWA/fHvhIhLCLJPnziOBFbFngilKv3DuSqVzkd8wyuMsJ/8GZvrUrZAyDS
LWVKd3OXrlRbcTJhlTGV9PAU6n+gEHIsfnZA2oW7PYoIkYkFXDkhMTRnAZdffhozB8hJxi1O2CF7
GNeHLhZZGXoC2Lhj5Twt3p+68cJwIZjFcp2Vz0peXOt19+Aws6B5KaxN+Li2zkvdaGRaKAJmYXEh
7cj/YWueEa/4eiwoWRqWih+u5Ca7w+MJdZ2Yl3tFpuXwVoPFUKlGPsqnLAcaU5DaFYAfJ3fQvTyy
bm6Djb8bMo8kEJ0GImWDGLeX1IWiwxXgLDIrYz7EOCkCVs1kJlQrHWQRvNAPhLi2/U/6lkHQcelZ
3xNBRz2XCAzZM6dtyU2XZhA9xVKgecjaGKoGcmcePqo3JbN1OM9kh89BRr14KwXAAgdBbCsndmxH
p7FhurtmVSgI2alBuyRqpV+kGxDSggk+3Z56p1MzV0zYlvU9y6Arxp1i5isf3lwiaH1KJaJR4Bjj
zFWsdDE8Yi4wbWGo7vGiaSIV9AcrOf6ZDAv14T3w/IAmRbUd4IT4ev+5OLPOmGEB4ID37ix/4plW
8l/rXcd2KOjfbDHqMAAl63Bjx4zoHm4airx9DffwrkWxZxBr+/k91hLcMS1sanwQU7pggko0rjwB
fUomlAP8gaj2DN9+q2l7oDDc+e9ahzc76KpmzuetEq5eHrdy/ED3v5BcG6TNEJZR+nt94t2ZeVS6
3BI1WW2D08cloBaVPAsvwGN4RBKoUT0eePP2p3TTkcrLJ4CakW3T24dlafCed0zhaWNVbyyNuKSd
A+NA95I+1yGvZS0CfaqK/Rfhqj1ApJeGv6UwyLbZj8RD598rV//uazpHsg4bZRv/wZF+/sxT5ie6
neJNZ5xifZjQvfiJr6MkLvQsYSYEJ5zYNUGFvbAGwxks+FvYu05R30MqhvfCzE0L+Akcxn86DzyX
Gv7bppKzGkA5gbbFkjrCJAgHFBotojWZhbj5nhW2GLul+qgNAUAJcYHQEbm5bZr8bxvHNNLU07s1
QGEDbq8mxS02vFLd3lo0Tu5aEM6ngC/yEDlAfETMe9+5UIn5FJ/jUsOrs5V7bNq1CI1Xx3NhJost
qZe7o/7Uwn5qTGZHtRzpjMcfmR4BFi0yd9hvrh6Iu1hKSc6U68+fISEHQii3H1o3pCGab/lez8SR
Ne/ngRnTcWRmo5f6cOG/ceOEakotIApnd/k2hDrDivKylO95Z84eEUKrDQR9FtKYUie/23tYEKx1
NIV5pB0N/0eJxQuGjMc7CN3xHEdDPDBrr+iei7zdwzpYhDG2B6++O3PEyWBiFqOOcofOsL8Fa15Z
ILx5WEK3B/3zK6loJOghaozmOoH97MGPbh4rmmm8DbfAKuud45ptDGfmBqMPBeGVQ7Bp5Pp/uLM/
qOK6k5SRz5RWsupG11i8ow/bt/moax4XLl3IFj83SUKTxcQJcamEfzvKSpeRDkZrMZeiRkHpay9n
VZwylxtmTCk0IVlnH/0L1rPcCsUisGA0UsQqzER5fenNh6lC+Xxm6CwGD0A/FgMjACHLHvVIzsfa
nlZhU5VzHW2SfGdev51muKZSZU7QVF+a6ga6RIcbjNLmGZ5rgX6WYEhQdwVxYezS3oITR1CvThCA
B/7UGziBUntECv108MRic3qHQ0doxfX9blv4aRhVo/kqkYmNJHcyqlOlXfuZF18ZcJxzmoJ9HM7Y
oq6btRJAGSKGDD/3Re4kiJSGHyIDNi2bBEYZOQgChoeANaPCvs+FEox52fAp62XjAQgPC0t77nwD
Zwx01jfd8DdQizr52vuvGYw5eqPfaTzeHVXA6IGo9iysExVcmIF3PWBLs24NqNYxudHrRi9f3RyT
hvVYpZ/FrsjWrtToTuh4AjhPpAvMSANiwsrsX0lV1eqCngZwmi3OQz2YlWuTPEL6pXPipPeT2cC4
OMtJVBWDYuhQOJoX0iWLrv6Lb9OkjopGuC1i4NrBs59kNpDlNvc4fYAioF1Jc0M/8lhQViSJw76Z
m0sF7MsHNitlfFyO47g9azAT+43lgHbvvVh26qZwY3ABlL2GKPD86TRYS5BwJjpeYfSXvZ0tdWUG
aAdARBh/yRlbkTC/mJ/ynfz27Et9+/ULf9xAKqXZEbX7/ZvKjPdDhWiPHaHwOFZrOsmidGZoSIrX
6wUUqQeVdGXIb7YVoedRSh8upEVn2DmuTRaRktl8rRnehDWDIfSN+37TELyApRes8btAdnTmVGnL
BMLCb/+xHTbXc+FX99RJhjSz2zVY4PBS3xTrqg7VIDl0PqZKTwT1hvRwujwssB8FLwEB8VSeDBbZ
HijIdFVNeeGIQknWTTSbzi4BbSeuqHIfPQ8CvtHeRe200NkppvzmLhLM2ZNoaHBrCyZagE8llqGS
4XWN5yL8xG2lf9L0Ozq3MRHnx06HCYDYKEyhciTGMW6Z3sXP2sJXwGrS4F/6ekrNGubJnYvv8UDy
1REyYLY9iUPN8UWDFiJ2OYa4Z3AZdD7H1Q8imYJyAn3+IgfpF/zXRyteHdHCYlQVPNZKgmqxxVeg
fPCejdXeBeLzOt9byXeP3ZuAuQpfwUANx4HD5i+GPNaeG8eQ5Clsia/HJLOmKYyIthInRXj+iCd7
e2Kixy6CYMtfUTfT4dSYGUn1mdUHERP6G+KrHLDDJw5uAEcOI986gR0J5mqJmWChz3ia6w6g985y
pvQAZJ9Xc3O0Amy/ycmG0qlRJAIYTgcvOrm9QwFRMOZd6OqqCebnbbn9CH3Jq0mQUKSs2Dqfw6bl
VRHSkR92oVYfKxmdBpub4tBU6TdEz7N/Ju8uMadjxECV0mzFs6+XM+pS09X8KH6DVSndFqQHLiXV
6mB9ROIB2vV9qZnNPZujz0zpokIbztc+t4cWztdH/fU7tvQuSyOMCsJOKvVOz3MonpCZXuYIvrlz
Mb9X/jTHiXegp7zGL8RG9vqZEu4MjXnjw4v+g87NQR65FcxOZG5O+oX6NOOiOmOrQ6Laz51gpZM/
wfiACWhhI2BizSmvuYgIXsZ7blFctIUYARKuQ/x9TRvSuYZs73r40eP3mkt+z+PdmsfZrn5X2cvx
vMWHtU2GrcAYXKdh3XmUDEOv80ZP2CLoddVWd7GStDNvxE1nqQIxnjiZBxGMUoRss2yj+nZxEM8H
ZvOZsM66AtFAtFFzKtzdibXuFLXAbJMJaOESM4iUTooei4yWNA9HgHqZBm0oJDsnrQMHO/RH8SgR
zXoOOJdWobWjI+S7eiDg7fmY1TW4Zw1StMcJ+Ow6Sd5mN61LPiobe2TtXfKnO8FHPjBfJ4ydPDc6
rlFpa0PRJeTp6qvLD0SZTf2yyH/F3dXMA5p7WjEJPLSJC+sOQv81maztoVMHlTITb4+kUWcysouB
/275UJzEAlwluBu/7Md94yfwkMTuVCFRDOrd7d1yE6ZCI/T1dh3b9jrafpKZ57N104SCJlC24h7z
hAojV67nvk7AhesrZs2mqUrIWjJccJ9Z+Z8RAtWIfvmtEw67PgSoQeQDF0PTzeqhQfbSEVZQC+cx
QTPruYsBfaurQh4X0jDVM9Bcv2vJhWcYWghH5LFZP+y2Vqi6djTcT1QPF8RNyAdlcxU8v4GXe/No
wRpWr/2A8VsYiy3O4qXC4lhAkPNkzBeibz//01CUXTBysiq52mNrMCKDjO/GTOSOEezagstNH5D1
TGJ1BQWW+jGtPtg+jjiqqzQg8FGPqMCsY+S+MGAEhnhP+hQqsoW1LWVKcK5s2QH+Y/uMab/47o+G
asq4gLzc+zc3hId5WZ6tzD7bsDHwT9r91hlBSvhe3tjjwNhku+iQhC0CN7B1pd0LCgUGmNgW6ovq
IGu0S2ySPUQgsSt/XjpR+ctqm6XAMNt/dp0hT/kbuJNxH9srgCMsTyMvgxEdyK4yWYoWHPIx53oJ
Ocq0Q6zFMEt5umJ3wZXfn+5nuxXYR6n3SDOJ9jp7HTzpKMj+bdUsCW84mCtx3mjyeRmv2uPTEukx
FMs8jY+t6PkuCEMgL2UHsFYziCg6DeLZHLrJ3hgnUYGhps1byATUcfIj3L/x4a0WptpQ0NLojJ8X
YYpw9psgsrOQGVmxjJeQ4FKece4Gv8h7+eF9ul8ll9aN+bekehA9Ks6R3AMFrh10KtZh8p/BThGh
6nebqDU+NWe8aQDrcj1BqVZrJOHEpsDbbb6AVoJY+RMq1jdt77KxmSUoi2fU7D8prak/WNEchnmr
SburzdphGXJEZc8q5f7KhdP+anG9wT/PtjRLEIEyGCkSLCY1hyBvuZfAnLfOE9Ippq8mKf+fO8JT
KS96Sk1HQj1uIhkt2jFiHVE0Wria2J3QKxw68swAl8+Mzs/ubMlZ1T7CPL/OBoj+3kh3GnK6CkoX
4FBAF4ASLi0XrxrDDYkCn97opZzee7OT37d6w1WcNwhk1a8x2Btp2UadB2C/O0AWnVD0F+IanpgF
MghLrURtsRrydhYa1bLZpjF8jGQ0hEgr1nzIQ2RZkXboQPRvRKZRSwsXxllcHeoSU15EgDPpZaAd
iKcHDkARDRvx7Mg91kjhjMadJ9+1EI+xxMKWtYFIWHG1ZvKb0VzIXFwoQ85LoJ5dPCx27/0lvgPs
vGjLck1YP/FktFhvnLKEF8LfkarRI1GiQx8emklEc5RsgVUdH6OTKi8YmehdzOg+QuGVOuPNwtAN
8w4p6VSdhpAsmv6S/l4lEPHb1oLMY3gDOOVGtb/jVR5wZhqOSgraqlknDO9Y9LXglCJmEjyoMTIU
TFW5ESGlcVEZpB+rr+B053gcC4PzUQPSo+V/pkUWXeWt+C2AQhW73tOM4jjWyoWJd6Whu5wZl4M5
1jdtFetXCISfWZxVz7vqfd4m3QGDJdlOyhE3RfjuxrEu6tI/S7SnaXxtKXUzJyM2nNoFv8CpH5ae
YgNaOka/kdcZkScaWrO64eVRT+zyll/wIIHkyi3c1wgwBixQCjPhn1en6yVMktydjFbFB20kHt05
Y79AJmB5/WkaJv714JmOcH76T0p8g1yC0Y/VJfoXBfxeQv360UHPeREdUvotQdYheA68FGA2wgxH
6DbOkbqe+MM2yxseg8dzzY2MdH60EThyq0urjaewLL/sgJUjSZhzcCvo4qoFBrouWhZeeMxghV2A
Td/b3tHJr+I7A/z0xrtC4sB4BlYewx/V4i8juLA2kVOej1ygExOvtg15jCR7llvLQxG4GlEQqqu+
S8ETs0bEnIv717Yt9sE+eSSY59ue6LuNF/NTw5gtJzZCTvUHDf4ReR/4f+Wjjd4mbWaLaRVBns3v
H+en1UeJCTyZ3PofJZsaw7LEh6IWrL4Pp+WKQeucxTKUTR1IPknLH9ifx9pxPzCF69KKFfPp4Sz2
3BP/FQcy6fwSs2k/aZ336gZwxhpg/0M5Rvz/Nb53eZbyNuTe4iD8fZP+4aHucEft/TmYPzrLXWxi
0xByXfKpqOL9wT+sg5OfOOcBJ5VIVsfJ14BV+uMI9quR2Jp+oOTKO7QszRA9gIPZWztfreBzioOp
UoYR+VVWrQ511SIPW/xldHXnVb1a6uKYG6uq18Ux8krdELUye8pWME8h/KoPLzs1xk8q/1CoLVe+
t29vm4tYlYl1MtKaHDP2APyKbbdeJN19YZS+rbSKah4IXr1I/px2Y08s34hgRx00HBm4TNO+oK1p
akVxMkD5GzL14cAcOYFtXPA+l+A29fDl6tg08BEsTLTPPykb95lEBovY3xGRSbGkU47y8eeFS/x9
JkYZgahpdb/V3gELgHDITX0IxhZj66Mhdz2EXFTlu6nTc4VO+fPZjhgG99KpVwz41ht3qI0uOMU7
bx3W8Q5gzwK0xRA5N461ZfsohQU8jGs6xy/MIJv1s9i6QSsW+vrFhbP9MEXHGnS3lDHk7DC/w6xa
fQvXjLq8UZ/RoUgOQRqydxgSJvBvdDclTToW8d35dTuR5fE+zPktaK/1B0vnnrGLAWnJRN7ZmL79
aYVAZm+hT9uM0SxdtF8AbZc2fst7q72mF/ZHsc7C44Uu8K3dyu1r1q8mc9YyCkUdXAZcUpyeFUiO
TYlCH9QQ1PRFpVxqppdT4wtFUBYHOhtGqaSgK5TghmPaZAxBOIBPT9qpo3A87uicvdWSM9Wy0ddJ
+FblAR82x4XO54x1p1YxCIndMYWWI2iWrlPJVCZe2+Y6h67X/OrmK8Mu0O3C63FLbmGyTf75/64j
W2HYGDDcD/Qamxd22BG8YG1IbpGAaSJ8dn1kUU69nA3+JCFEJ4OXR/VA3aHzP7sWN5PgjY/JL/B0
s74M/0IsXE4Wp1zRt7HO9NNN5BSXTuY1h33Qq7tc/EcJ8to7Ib7SK8DnCTy0IfRJbpEq5qe9iaaX
/SwAW8Gal1C/UVK1iKRgcfTf+aTZpaV95lreZtF7dT9LofQmebeKQhP5zlNKRQCQVbwghVCobWF9
5dIVOWuw2LbjmEycC6T82FszR+MXxE6b75xatKJJSP0sIEqxott7nckhqDEA7gC1wYXKB6FiqMm4
FePp93Fo+KoFPCrTUVbP/OYmS6YxWFCKK2qDnGPSsbHP2VaB0MPujo4XmqkRBkAGX+GrtvqWT0ea
tYMilTE2IotAwwioHeyYPlkYW+nbz/TO23QGouTwUcmwX5yMr41diVO+YDLKPNRMpyXrvwfqqjoH
lNoT4EAFCFm7ZI23BH+j0yb8z4Dk0v4gTsFsl3blardYwUbXYPer6F6b7P0RvThnSmC1YeKc4C22
x3HYui906AyV40Rhn0uMMA0GwZB6wxZ0pt/+KWQILyzmZW5kTakyQAJBoFG0V2zR7LZuYBFDUNEQ
YWUfAxjtAlyg++xWVS1arAk32sZFW9vRZeADYWFGVcTPcNAJQ6B5CvYhQtWy4wznwO/b0TtSnCnS
n1PvlycRwNCG8DUsUKhczjB4YDBz0E01tSQT6j5Bm1N9A3tD3i4aKlGB1o510VpU5F8KceieNKdA
oGwUKDgS+BVc9bUlmyALenoXjb8hdF7+tXBSohafC2PmORchMrS0bVdrbn0+W0w63STHeNL/4Q1G
mxulsvPJus6gSWd85C9J1L9fJ98HldgkdbgEW9ZFiUz31wYm/1HpTQXntzMfgZHjV2t27vjv83QK
tMRH8jBDfkmT7niV0Ao/21tg40UQGCPBwrg+U/T/hSBNFhc0+aTcSy7PvtEs0Y7Na9LsjYluSbuG
0NFxWEnccryKj61Fx8wjTAw6dB2EacJBGXmxAdZUliQvXegtI9mboL8nXjMxw2IZhVdzwnjk5T8o
l+9c+ChoOwqNOcSAMyPi3N4ZcG1xtBrF0XofXuh7XrvwZHSERpYlclRPgrevT0QnFRgfFikwg4vI
x/bvUfsHpFFQ/D//WOUk6uXa/RXQFloDCyuXY1QHpDZ35bazUx5Bm1hJc35csqnXcv78Nkg6boy1
663cwGAaLj3ynvvu178dnRWBD481EBQ0zhrNTYSzNKZjcquOpvwVzClmYFoLJvgKVhXAMbpkFRS7
Dz/8WhsqCRXBmGqkP+2kPsgyUmMaEWHGS8f5VXVvQEBTdvxkkPe1mMGrLVi0JvxWUizq/yg2Rh6C
Uq6rzIP2ZEFQaB6HWTutoWmXb8bdQjxMt1RP/gppoxslk85HVZqvaPrQLHynw/ARfcNI+32vx9FB
+UgdzoE+LmwARyhhDHNld+1KDa+OwiiXihcHwBAuiqkIY44W/GNwZyyxpo+MIUIzZygEVW5vG+GG
U9OKLYYXDKHqAI2g3qLPzUlnYlcnxQ9tgQR7oIVeyBd8yYZHekt5KUO2BvNY4VfboyWRSW3Si92S
r5sKOFwRZcZ1aKQR4Q2uhZPXtNdP6Ai+KCd01JHwR7R+eO9DH/Ra90L2fzF0Bpm1HuvqJ0E9h/uE
3X9WmKGD03lCLJQWXfIacf554Y0u+da2JbRvBRqTzehFKFj+Njj5Gsl6v9kENrNLdjt3CBFMcA8S
lODwBJMUvVgj4TYfu8AI0BX7akooCQ7bykGwpBL+Uhl3TiVvIgTE24lIh88J4aFk8JDjsdGE+eWJ
dZpZLsGFGjFXNLlfJIEhVVbTokEnkSx4dfwcL5zRnpYGK6VaeE6mbA5fGbRkBcdRs7UnaMjykTtS
iijuBz+DER1AbmKmUoAm4k04h7YrPPFEYHQlMrCYnYZ9Jvb3pvajScHSuseFcHpYnBQB+FERvRFB
dG9UXxGd7I1g+BgvyYKVhVvXwDcPbZ4YBX9mSwMmje/1r+Urxx3LTXl+O8PZ4gZ0+tE8ICIFiSCs
0yv1utcym81ppXTutniZF45PRxzflTrs+kReVfvxVZvAGe6D3T+9ojPmWBFs06VNUHBAmviEXIxO
vtG+2uFU5nSneEGVcZxZP7FKYcPUuZkNzx/9fY6hv0UbY8Z+kfV3fJT88FjTf1xJpTPOTy1vSTno
OeAPnr7wAU0IzND+1i0KG79M+Ot2m9IupGHRZBAb3aD4zl2grmAauRCwnJdizvLFGDVXhxpbtgsr
GyiNjqYNJfAccR1o+RsdRWmOQauiPq0WhTr9qkoXUz54seZqffEmXcuDJ8J6MgeFQMN0Q1rA97on
CrAwcHWiy/mEIziz5Hmg310AUf2mIJgABBrlJRW1XrPS0nkfwP9JYIc3amghe/HinHP41QsGNKic
q9LdoCVSfOV9ksR3ode6x6Ryjj+b0piz7YWDVVsv/PXMo69dN0VBny8IzScFWAjiNxNhhUOjBNuh
r8CH2rg4mR6Kbd3xqr+/5zASzT+i1TVijHeISnrCNcP4SofoNkgcb/sWbOX1KGD1Z8R5KxtRxKbx
Omnqg0vccgCf0UyKUus+PG97+4KrTjXH91B4g4XzNH2K1JFmJ7cKocz0uV6qkau3uzOn/iX8KRRO
ADfqsfPJwIwtNYw35o+Ym/k8ZLGYlHtI6HM/GdqcD8tmn1nAayGAngUSJ7nbw8dMxXI2MuVNrQxf
4ck4DL8tit6YGR4kwGqN8iKxVzuI222wMMwJPxHxIqoYELfumJheQE38+uRJWBX5Q9PiFjV7+2NA
hT8deSArugD31Ugcv0CXMgywIHPq7jLPeO47oCCwVhSqVArcUSMqvrMyVzDp2q0pNztWMDFbLWO0
gRFci27jS7iPLSIm2rzfQyMOzSGWSxb/TpRng7SIsHGsL86b26p+LYLqXI0rpMcDj+q3eEpEAhjH
VWbuZM1Z8yQ29EkcYzH6b7FJMrhaIbS5ji3/zK7fB0Fk3Kcw2BtqcAZR+90g4uLJH5ROWZ8nIaia
IgeaomuNUkWKU+GYv/Aq6etV024qVtiBkt37H22ly97heQyQrraxICptwfvvqOFByzNjoKefldGY
0HS7hOiboUjejL+e0t4YXr433Urc7mRKXNKoavEmboJZSz8toAvcJKkM8Imzf+UqXs0y5NBlsQFu
+6KCxNdUF9dSq2wsHmn0zll58jmfZnRFoh+rty32jN2TPqVoWxd1tRukvQEptBjMg20Fl0GykUrV
0sRpzvCXbjffFt/GNB5COneUydfeU/SPyG7fuRVy41RJh3ZMfZzMGESfJs9r2gBQhHRPxsYJ91e5
g2/M/Fr5jygASKQ/pawa3r0EdAosWSa3GDz8k2IvoMCtH3rvC9btprtbob9qEFA+b35j8cinI0pZ
WPL0rBy1JS1J63TfM4ftwd2paQf9i854oPaAdphjvqn/bec3Cf7KTJXEDz6WvhEyto25IiJOYuym
W3Tzhww4Xc+yu8PPX1rTVjAcNkKAKAWjez8xnZeuu2XqB7CkhJpwbeNOEwigufKbbfI1xaXCK980
WdF6VnDYTOeOpiaQ72jFK1xgTDpRPGkEpAtal/fBQ2inxRZ+n8TCZqL1OHtrNnsc+zH2S7aXXkkT
qCEQEb0fRvJNev3tN8u2KAnTbPIUbJYAW4AJ4Ik8v/GKzHUEkAryK1dtixJf6rEi/xig6FICM1ql
tRwBGLrZiEgVyMph7cTpPFebz+kW3frSbNCmFL3k4l9Us3lIa4GCmq42EadhEsF4pDwzAfVRVPqw
tFOr2xuZsUl5DPooWHOMkKQJxsMpySxsuS7/91/4GyawCVueWxInB3RJzCpE6Rkb9gBObsZttTqu
vS+z0Bg70AnM1oNHRg2+peywsVzr/I3HLYpphawoz3d8sHUNtjor2UWKRsr/7ou1phdjb6QyYCVe
Qm38AnGwoHgTbqfZwPz+uxUsoKvBeVrUESwNWqosNK1TfYUf5SLwxnvyV+pv7MJ6cAEzkWUU5vOU
VNdsnUWo5Rd3iuDWRm/dydWCfNkrEXVVfCV+FwZ+AooSYJJVCUNfDsxjKHTUew6Li+xIjEJhKucb
1ff8ecNmJ+Kvbgud99HqnbAhr9+Rq+Orwy+beQ2qoT31cRU+eLojDr5tnwJpIBRJh6JOb2jL95Lg
jUtdf5C8WSyoBTv2VqX8uPGc9k53UbJitjyyjk2Lx23lpKGIdh17NASHZ+V3Hz6WmSzd6bNqdxO2
ki8pLiJfRaBNrI9X+rvDci+Fkse4KCuigJ5MVUjx6dgPn4ZfGRUl+7uQ7cgv6G7Ws/QtHi6xuD6q
HcTsVwINtEPLNXYPZETB5e0GsNii+HBygIefjWt6o2/BjG2wsAhW0GYlisCPHlWyGAUnB3Mp+FIu
aofeCwGf1FxccP3L6uv/CWIyEng56rAgRAdZPSbmOhC2dNb89snLRf3DI4dILxZj5D9yxiCv8HFm
CLk35802mRHjZl1WPIsVeKuPg/JjuiOiWjUNJuxRh8E9Y8ShWMNYPvklMH1IFewaYggrcwx2oost
YwLX9eAUTa9G9LsHaZBo+t5fkmGuqBgMTLfCF7Lf3LIBjPQ2Vpc/BVgQkSmOb4KNw4XmPNJyylLO
XWLgmoJxt8Jd5YTKrqr/4dPanue1Ko9aT/eupcSlkxJUdc4szmnhfWoebFkuKvrmfMVFWbvQK30T
PGmDjfFpGDl2dF8nrct2pSME5tkTkBmYIWcFs8BuwQH1C1VbBKH3R3BiW9Nvadac9GoxlHqm7Rrs
0k4lELcgzOKJxzm4o03SDlo+ZanW5kTHWZDKzqnRa9qQ09JafN/Yx1uxq8mkUYNS+ijxRzW/LiHD
9bmskhT3Z4HCk8YsMejimbefESOXl0PaS58+Y34tBFnplu4ZGGplD15xhX3Z9hGjxWf01ytZ+5nu
m/m0fGVKZPexVOd8JoZVv1lDqMa+bJAWQ5Xi+8LL2YxrqLG3oEOkL+yPlmJH0l6QJfOw6rBbZqOL
C6c1qXGC9Zle6hkgUuZ4HzVJ8JHGiTBbs5/rX/rg50zloSDpYuif2X9DpO/csM432Pf3vmgjgNFd
aqRL9E3aLcgXL+YcY0vdZ9kJ5bJAGuFCGrOZ5V78gNj12yY/WcWjz2/sohtp6gNyYx9i8d0PcpLT
tGoJuAVh1mr/t1XnT8ReFcJFrPpOE8LyQ0S59HMJM4I+0k1tIYla5LHLnN2BFRsmuWO9sl1C/qXI
bZKC5BiahQGgerXpk/ey9RhS3muq7MzOrVJgPyaAt48k4+/LrrLG6RVC6YLfOH+2nrthrwW3KobR
0SG0gZG5mDaXsPLzGPmyZExIBiA5JZmEJKCwjMmBJU/bO+rRYHJQVxTrWF4wY9Cw7J1s4lVpu2Tz
/w375Jxz4oC2go4k0/KKBmIZn04tTbfRbyz2tFYCLx80zfA83vokZy5yUrIIX5CbkH4tBBdAuMB9
vBItRKYQWprfeUJCptcsS3f5bTDDcM4jforB+038fPIDSD6MSdV9D4oHB0NR7nXLfn3xItCoVgK7
z8wwIsE5NxvJKAVKqkeN1+fYVHYPENpXSh8JXyfje9KB8ySdoyKxmKRgHofOWl6HHVkZaid34xK5
2O6T29i99rzIbWTcfRWBu5spDbH5Pradk/Sg3gXDxG206l18wsQSph4I9M1H6PgbrQEw9j3KInc1
NO9aQxiRm0RNy/vE6IPJNQrzWElfXvm31Wlj05rjB9olWBe9W1ah7cnkxEA2VWMn/+kPkYr4IevW
Pqa/oWju+XsKRPd1oBX5nlW2Sxuj42WIcsyFUut3RVbMoOvSrxCNa2WBWyMySESpWsrw8lUMQjyi
NBevUMFDPK0a5ed+i2+yDes0Kaq28BSWvdx10PueIqjHxy1VEhVwD+xLCRedUy1mMQL5bO5HF22D
+hNGABjJLs52P4mpWnZvXUOyqVaIGRINu0JxLN0Ze0Of1F0gk3DrtiZA8uxZV7eZMyaCpjqWeDLf
acoh5yQ/Hje2tc6JQ4XQe8gVTecjNHQfNFulhPi1yM13XErLYb6jVQX1ELAckbwSDurV1BVpI6on
bO0KlFui7QdrHxcSt1RceAk63StW96JjfzyKh0vZfn4ReR61pjJKOkSmRgg1oAt4KKQaHDYlShla
Myvln5XwD2PjQkiH9vNFAcFGCWyykTxHUmDbdFD0Dcia/R+f+aAASEP2JcAPgNgUDArqeaUAVkpQ
7SprkyfoCb/mwLJfC5ZZ+FkRji1PkB6vlx6iLsfA+XS1hmwPPSO2jXzhZ5Chg9oC3nM2NMGHzZ5T
zc2DLK7eBw3s8Ez+EbHeB17J/NfPvOsaoVfO4Q8uqzM6Q0qZ3hb/gZaFO8qrw7n7k/jK9GxPjJDC
5GRX8flF6QQLBLE8NozdlSUJa2cXlMHEgfPlzmD98ynuqk7yuG6qSLtT9OwGXL3KNki0hRKYn5Tz
UhRalmDt2hmFSueUlqaLTQhSTm+kr3/aC8CryU6u/sDm7k5IGI9PHVdGW1oJ2qB8mwyREx1HcXEm
QCYK8/W7qjrVNpI1H4M41Ev4ZM7DlKKKlUsdVlF315GQEWWaNcOJoN+Ssi1W7bk7b0tbiWIardTK
Zq2NpkSy8rBVmIzUSCLpt6up48C9UmlftTaE1zcqM5tqmRnFuMuEvG5go7AO3BoXpneCGVDI86mI
+lMCkawCzxXWvLSxS9QxZV3v0oRkIUkpzj43g+0DBiAaNZLTYVaKWv3K4TNhdyb5GL+fLFCT55cB
bS6pNqqpH+ZT5lvdZmdjHolYag3prSQTV/z56OwVvtCslqHc8aK+la1+xhfyGoURI4OdDGDHGR7V
HXb9+DtMtwlAPCr4QEzd87KEWkq4CI6xems2ZcYCfW6SCK7cAmBmMhvXYDwoSLTCVwdb7CNdZTEO
hQEgK79NAabt+kbod5tVbvoLVfubWkAJGCkKd6CcN4PA8vDzh+gDjIyOe6BJvIkoAxUl8YVsuhRD
OKGp6KmZSGaEksG5l0znBQnisHD0tiRoMjdoh3C5kMb8TxXEqN5rVfC/aCOhHPJhYd5bNN7LVKmX
kMdLzfeZlbZHDjRfKrcHMoetkSKmUYW4paBixpJyLeib4NxVGGQNwUVOy0VFyynfaKLQzAe3M2mf
tUJIicG6Afe1vlUmlKOgwBZpmQh+lrmcxUxdGNByogOdIDKJo8XmYMKrNL4UT8O0cK6j9gn8F474
z6rXGK7ywWppw8miqh8GNyaMCWSG9hieYU8FRPSgKn2pLzPCcZGYpJUst4PaHsFWqZ8o6ICZ+DkZ
rw6JokSnq4KKnftzSd6yRxub38OBUTsW6Vnqe0Uj9+qOWIUUN6LneAXqent00uZFliQHxyZ/JP1/
P8grl+ANNBHwgKFe9cLkK+y61XhzkvQiEQn2g0lr0e6tv4pGUo9ycI+xdHDVwOGl9b+0IurTUEkM
oyDaod56xDnBLJTAqE7XyHGF+e25oAxaanzJ0Y0OVJdWptWHDZTB9OcnOS3+mCWAjPDjSdbfkgFc
zGhiYsYiVRxshsFxUTt8DxXVtWCzFp6onYjNZ2rCAdIScvkSwRCHhBtDwUzbXypatRQN8JrLqNWu
qG6tpywy78hemHWupOE1VF/9JTErQ3yyMus1rPgXvAxJremf2IjRSj/LQIvsRHBq63SMK/WiLQvZ
XwpBEtjSfCL9RrwWAuBdwRaiAyfkborN5WfDXldJU/R20tk0gmuCorLDz9CZtstW8OcqAlGOzDjN
VQ5P588dGNZJX7+GEzq4UCvaJRBxQ6943MYo/VIsWpRQdGGqb93C7dTTwHpxQAZJ0zM6D6+2LYya
Gp04QjDfNbN0b9J5OJNqn31SwKof23ZHb+rWIED+z6Knx39pMviro0+tU1IcA14rjmkGwiDrK6ib
nYTjd8VxtbkxRskY5C/dMivlA4wNMdrDkAa2UB8S1X6wsKM+WFuacr1JDRlzboENZZVJ2HeREDKC
nXbNpPry2Eh8xuZgykaGTslMaDZPjbbArjAJuRSOB9G7wWf5Wc0oP7dTqbyr8/aC8xgBH+akdPO7
ptOD5B1PGQeGW/LHTy2I992EgE71E/OzfSWbF122gxqPVgQWCIiZ3A1DTbZyLMGpmkx45EabMIsD
BW0ovXuT8RS6Pd6fStIhXSOm76U6AGuHwaWa7/rDvIg5IhgueWMUCDd/O7lie9b/9S9T7/ix6o1H
SwXtB2ud50d4scGwghjTqrKaIZ0zM66EtvxT2gvhHlkpFGc3HQSCyzJSfOpeRo8rvez6E2EfWOlH
Emj2qU2WSEgJEjMP3bGDy8stlmdlmnZ9BPX2aXq+U/0Tf1njayrSjkMEEYwNf/yivHs9uPGtqsOQ
gXRkbEkh4utXjY4NcZbt5C9daJZnD/gr23zcpPjrGImqem1Gr6IHhSeahtuIUV9mMqRWLt1VIDwy
vPXEjAIGyHTIyHXYIQUWaXQmeKbH8SvigPCZGFynrLVrNsw8uwthfi16ISlLQ/b2TOW4I4XO6MBR
MJkEB3y1a4b7y4cB0dU+yFENQD4Mg9GjrleHw16FlT7IJ/lu3OwkxpNE+WRA2GSeDsn/ZJuV6AqB
qFu1ZJJ3e5DFUvnhzRlHBGiV3NSuJURtMXqbrVtllmKa/WVAj3UWS2fQEWSjmrbdffVoRuBslwEu
eE46nYjVOr7ghYBExdw8Spb5mKdpSMPIPyL/pqqf4UPBauSgzQYl+hsKxMX1RKlShdyPpQFUBUdk
wFjjw2q5UWqRQjkVTrRBtOI8SnhoWTVU9WQTe8HavJEhKQO4uS6IiKhYoQT0CpMQwlKup+p53iS/
1HAdCAD3PeWvyC0ial0HmB8fpAzXYeJmRmX6R+2n/QQflHYL0N9X1yd6dHwtgl6kzOlK4NMetTNe
Zkv26MHYgjGnD1diNAYny/SgSd+gwHy3fySJoiJMzMsQ8ZVY+ffZZ5cgRGwAFuYpFqND72+Tp1cJ
NMTpeatTak53vkbxn4Jqymnal/pKQ0dQCERNqL5ddIMjA1uR/ERvTGjPnXAGKPXaqjrbZVV+LI2O
X9V88dEdVlOJcwHGBb6KICdXy4jn7zIPFT0qS+iygxrYFUjVA5LhvyK0n3CTwmn9YfzN727+jHRO
p61RDX7r8BRvnXGYWOWTSRqbT52JATPpQDGJ33leLVgiIteVV3fRb7XLwQGvq156gIRNvnQuPDlG
0wY8gSsAmEOfVql3MLp04NTkX/T6WlI0QjKZwnkklj9sg2Ynw88gJxsc1NMnWZxooJ47+RovJRkD
FAfiU9PkfZcSS7WgHcd32jju70BMc3cw6Q3BIRnPAUCK0d6ZyEb8ZGpuRoD0sXHf+qVGbBmK2Dps
wVLqg+YVsKmdPYBCKoY4riZt4NjNglThUaXcmsLRLc1NEYQSjV7NLz+AW5P5UhEJYUR7/jzczgsX
jC4/eRx8ERHx2jSWe0ef0GYJcCthfSbJERhpTF1VGPUpafeIm3p2g0u41sYC9bOHomROIPZaiPnF
tdk/q3d471ZaVhnqf6AACc/ryK+XE3+ZPR253jRhqG4IwG+YmCeeb6HGFd53eCWfIHxya6DY+dyf
sxPzGfwxXHphXbmWIwZMiEjx0gv56Lv48IIJgLtsczKGbtKc+0KHUQ9uS0yv7BHjRbmrpg2D7hX1
yXe8Oq3U7Kg1xuCOEy6nSTkgzuZ/v9YpNQFf72qi2tmeDKYpw5W87nFFJgwMGY5Yamgaa5c4LntR
H7YKP9jiUDGY0VJ2/+oG9CmfKe7BHD+RqnqoGTuHlF8HJEzsdSQUPpOk2H/D41LStOvzX84YXxKj
rkOtD6Z1OT28pGYqDmi0m+NzSXFVujb7cE4rRj9JsTNAKA4xqNSnGo+lwRTxITiMl1TTMJBHHwpx
DkQgpt/kpkd/ky9+dIlNzYt+HhM47yr3LSQFZZHDvpWBRyzdeFsG0lyMp1AoLaBbT3OyuvClwOmi
Eu6w+pQJE1RaCI07lPi5l5BuhnO2dXWZuipKtUbcNQ7miCXM0+ooPMwaLt0SQkxlTRzw8tZbxn/E
/PB7EjkCwTL/i1SA7WUx6XQrDTlkwp4quwwo3KMFI2OaDUYjPa9rxBJqASnTJQUMzxtcFJMVQVc7
XZ5cJdAZN4pXCGyCE9TzBpgiYNlMOEv5JJusFd5I+DL3Pj/LXUYjabPqXrShTdGBGO8/SiS5wALe
gCkgCdPWRXG1RRSHMkZ3lE5Ym7SdYDKnDv8zOgouZH54BBf3uLRTTQikRFKww+ZqGDNTg+kq52/8
7pjtw46HlzNa9YiZiNUMuDzuEeuWyBmczmwoMEUkMIeP2ORNVWsJR9mQ6zamhS3I+r8qKG+Pti+n
55NoV+MWq2TZoGj7MhpLCTJY+KwJhwh/83sX9jooTA1VFJJL7Ub5+EJNTJFLGLQPzolk8mLb2nwP
B2dKwgbnJXJAQ0reY8KVQ1RSQrxFgLQAfEMulfeX/65CWdS93Pk3O6eTtceJ0LGoX7PqApJYQVQj
1V41StlEROejwcm6x07vYlBX2qsHX2+5pLS+xIUNY0R9xX8PYROYVa/t4qAF9NJgOjEN0/s38x6S
/lzB/Ka0hp6Q4QuSxrFOoTRXhfAc2KeA0AhAFW3kn7u19qpm1K92nSYKtHxBwiRHnV/L32VhNQRZ
iiAk3fKkA/Pm9EoKILk3SVIl3SK2FzQopJeu61drp4TdTjpEFluyoTT3gDi02qX50oO1bqJ9Su6N
nnN3CE37Puo/JUy3rUVduwGY92fvwpfDYyFr1UQvZtPyPIXalny2TL2oK2qMFhtEKClZQsy1/Wb4
7a42oYK762BnwSGZmMKWTZlhj5GWsxd2IyaWSwXrIP+NIv+jhrtJPZq1GEdawLZYC7gQ2YVZ2N7h
UoSGKb2ShGbG9VvyuYwqfoY743loKwSL1iE0bxpa0Q16PYCEvMdwV/tnlUlqOdPElJw/7s+4Qa7t
916uf8cg99yr4gQiHT+mjYL/KHtnyX1bVQHBzH7YnE7R8SQJXMo3fE7OGF8twvO/enZb6GFacLGp
8osdHwdoZWmojJBrMHUb8iT9EyL9uwOOCU4cSlXW5aWC50kzfDlyT+eyhF91EKSkjdZG4P+4Ffkf
2kUQFuWW+qGSSgrc+POp/1nwJWOzXufFBg9EQdNeKlllI0BdqWJUFpb7n+jKKWLRDffy5RD6GAuw
n/OqfNNp3yovAIgtMLdOGIYzX3NOUGxWukr8CrFUOYI4YLRbSEUmKJ0W+hFIwU0lTrWWKpZAWGNq
pMuJZ56AIu/LJvlMy3Lx48/GYCdadrh+1lK/mElZo5Zkr1XU2vosmyX2kwbgKsGXtAIJBMSPsSO2
kHZugzVEcYQ8LEcM98UnIaq7ltqwyOs6xHByj6BBLLkKrn5cP8a/PfMBNdyYwVlNaAzKDn2n7KLq
zwrBsk3A14ohmv1ShaMYIp2P866kVwFosjqML9lm0UrDgUQZPEGl8RzwhuMIa7EzCxD88/pTGx32
bRi4RPdpz7NdyilU0R6QzxekFsZWEHP15EGPk4t0dFdjA4+5JuCN7T1z+HLoHhzC5pNzGSgS0k4Q
4FDVzLUoSfXQ/k3fuFdjaTnbwX0gaKKYq8Hrzrz3k5Hv3TSZEO9tSxwfy+NR5hD2+pFfnMl1RRTE
mKDjJvYZHWIUh+d3QYEuXBIHwXLiSlA+aVkz5AbPhCB8NJWBdQ2g2/eoZPtg81YLVhCIObGJdGoK
FtsdtbZ94aQPraQNWaPKRGWk1FNtrR9jfXYpoQkTPdRQiRLfvU0TJFLA9MUZjFJFNoIoQAHeL3/y
XaU/coSO3gWP+Oxv1AkHKAnXj4VDERziWcuBmCdqW3eEMUFfGMubxXb/YsF/ZJZ9w98wBbUrW/mq
EQO8brxY36IcCfVMSuzquwIaKbHD5GlyK6kGQpgKkWzJbU175Hg3MmDpJhwAD53XguUzpEJ6bT47
Yh8RkTl9nFMkO0hfjtjLXdun70H11rdVFhaHrOSQL2+zZdbUZ4MGpjy0RFRYx/At/DNwfeauAW4I
a7lUV9zNWILisxGII2wmVp3HeOhxWLcfveBUWZ2sejfvpVcFaTwLNVbhSx+3DgdtFYxCYJoFrKx6
uQAeuvN6UanLW3YCH4WqgYyHPMGhO0AR5GKhrigNwGL3hDB7k+Ft2tbRrPDh09Z7UFpIsCv+JiHr
peB+TWL6GRt2VRVte8jg2vJT7P7DMbKN3fUoVxMvUcsk7oaeZrIZ5qHz3f9Hpha1UiWGHhxD645q
u7+/UMl0gsa8M0RjHlSlLeo/OiphsFxSCenF4sTKrG1V2ET4c+TL4N/rU+UjZjrR8AT1s9YM2HEf
sy+XTe+rFzLrLF3C2As7e3zZzciLLUEr+7nlk0WkoWZjcrhIEKLIprKL5mLQhPeOpvODw3swox/3
9uhyX23mIDJi1mZx6suGD1JLspMfdfiR7+/Kvm/NF8r5aIg02WyAssy26Spru0y36ZGOh7mBOgSh
R/bJ8Eo4831835RrBALF1YjaEFd4iy9tF/m1KnqsA7k/ss1nb3ohk4PnPQ2+lFVjngAL1uDNqi50
cODfy+ebDikA9tZamVMfui6nl9SOEiud7Saw5Gyva6sgO0yQE0WfqjS94xxvg+fWIifMN5wEaNxz
TQLIW9neugxwO2AASpn3zLKEniKIWPP3DRbQxm4HLLEKlZqOdo2Cz/8Q4goAnIsLFwqb+khVReh1
ifhdM/P3M7ZhXCBArihpUdVjHjSje25bDM5RxvsGXufXbDj3OPmbtN6SxBDia/xr0Y5P/1UtQLaP
oAmWPRy5BPoaY6ItpW4OycAorWce0P9kRbL6zAAMf319gzZ5tIyGDzjA+B02TenHePasvBZVkO14
NiqPpGJCkosttDmDkNlj9gW5aLSTNUI7iRB/EE/HKuv+/2wCSoedWRT/hNf9t9NTwbukx9hddm5z
SJ0qWlHg0jbh0RLDkSwurmn6sArQY+b1oMoYK4kO73kPdMqRNogG5KMja47uCVQOHy2WW85rjr1r
QVuSkcOTw/y89svaHPB0K//P2l8FA1/gn61oX0WsUnKIvPy2CPZjuRjTQtgoLMLg2OWU6VAID8AE
MzeqPJPwdU39wVB8U7qycaCN+dNNn7uFBOzr0y3Whb8WlIqo4mpFZ4k77UI1lULdBNNEn0Nb7YKa
H0N8biYbDnnoQg08xvZpuWNfd6Ft7diL/B9rgf9li+f4tB+MU4V5CR4Im3+0Qy24z+sObhD14LWh
FecfLXT9Qr/ppJ5w5Gww9N6ecob+L6Hk0qfaMde6A7bcAnW+Yu5Zc2K/x9MlTlnJ6VYo6MAK3Z+k
3MWwinmIUDOaevmnOiaGkhUss2JNxjteEq3g+3M6dFiNSuhCV2y4FAyyp7Ac5CC/Ih80OwVQyDY+
Z8HgozFheWStqEc1E7CTBZ0NQo//2ApJunAUb/rarmciqRMdxx79EqIbXRJoNXEF1jBcWaHPY0P0
+fchTVjQrs8yCS8WNuNytg/61/R6whC3sasIrXCfVYQbOuj7XlsJ3YQFUpk+lhtUKoRY1GH6bt6t
oIbJTDuup9+H5alfzBCqqHNaE18Dn2bsDB1LSpnBBFQdpj664PB28dZYsoyPIDc82uW6xX7NUP7V
UQP+MoH4wbYdz0VHU4Mv2XPMo3ex/56sbS3DRKeO6vp4Lh+yeAogUPRlEvKQIQvrxCl7TviAq86x
lqhYmeChfffXCVJ7ES/icDdcufHPX0jo8Z+pf5y33qppwPqloJI4YjQ3F85jEO5XUaca2i2i4bcV
wDTQZMXVrksHdcyYbYHkRNtNTIK0XExWez1AJbqT9Lbm9/NDst/tc3+wCFw1PaUIl0t3+3Bl+LNy
j285CVRCiAwT32KeQdUV2Hk2OX4j0PpWfAhblq3tO5wPQYFY8BOtarVmjhuZSmiqawXJDIqNBp8S
hCOlKJ4gSWmpFQOwBjDw4pKaSN/MA2YjjHTZbfthEi/oLl9e37SL2imLZN3i/rQWru7d0B3BWTir
fhAMaUiBJHXuoDpmxWelONzNOGFmuM8i7shIs0iwVzL9v82+a/hWveQFjjF6xS/M3tXXtETiQjA4
+ObtrPUSINjgvOsUTcbVDHMydxd4zJPNjoq2Nrsj/7vcpYcMniz8pK5oC6GAL2o3A1sodSm1DjRz
MfUNftmcGZ6wBGScwfZJ8Mnd8Qk8VmD+DIqdlo76AU4dT9AUx/ewcGyF85HOfGh10BpgsbyhTJEi
FoJECQC0widdmUgwtqqQi4oFekV/qkvqZdvC5245AsuBUh7w22Q+3EZ04GSnzOJWy6TykV01E/hj
nsZ2xaJwBWKltvvfqvZ0V6oNFgG539z3HeqH7IMmpI7amuriLqwSdor5ngGy2cuDTyHqK1edYvS8
WkkDD9o2VYpgF2KPNb1UJVNgZ9F9tMLJvRgyZES3Z7yMoKr7ZW0SpOjPyzTIHynsAj8Lrm5QajSI
CipyszUGPJmBJ1aHV6K9GmX1hq0YYPxhwsRzHyVQVr2M+Pgxuly5ZaTFrKgZ0AGmAT2xxjqXok6R
/4VUaRSWf5joCeCoyn9rBCEch3TNpMdizOF1JZMyLbw4/Rr44j6m81582qSLYRNrXYisxP40XsqJ
X72Eudhj2Isel9N1UmjHaHb1rA8s1NCLLKM2IxSS73+7ccZrBX606yOLHzg866C2a/gE0+VEPiXK
LqmUPwng8pXrQCW5dRudxnWXq+McyHCFgLxbQBWH63nPYdUOsRZhHC7CPo+737wA/mF2B1PQRlUM
H1iCCGI5h58X9wnh7Vd+ZiOOdHaNjU9a1QlN+yJb6jkePsAl9iEebe6xSbpPW+t70T4a/DvOd52j
gMUCm0gwvMF6gz2IWVgMWLuKwqoJP8vOaya1btuvpNQb3TluWBTcBbNjU6Puafjo1r7Sf9WGalsX
sMtvQ5P8crU5zJFBtWlgijQKejuweWVHIs8p4/asV8PmK0GSZbZb0yVNw9TvfnO1GKeYJ/iEEVlS
ub3oM85+NKjNkFUn5dI9TCWBvsuo+ZRjUwDk8Ox7XdhX+acgFlH3rKpqUeg8Jobs6d6UpWzxTS3U
tRfHtno+cfECK+MHga83VU0UIByJXCQ+X/loyqFezIymySwC2VGYLgqzz1F8bnBjudFnxnZRaT0e
JidXBN1XMtdt5tmAE7WAifBKio5dvFrcjYJkwXhh1CZib0AhY4SfYBZ4VbY2/u6Jgf6G5sFBtbJN
L4WrrfWzThEN0pk/l9JDwyvXZEZG4qcG+fo/uGFC1ln5f6/iG2Q23mwfnX3FvYaZi2RPi2fAPxWR
ak54VhrhwWQjTU2fBPfhmkucpI5uA6DArVcf0T4peiTV18/heqgTGDGFsfBULye43RKSZZZmI89Z
fprIfM5rSZr9GqZ+5Y29Xrbg/5fDljZjGyDJ3l5U+p8ed4Awy63B79RipA8z2c79R65QNl2l+vWl
JWdrIwqa41UtbKZ7a8fb9Pbsu4DnFjgsifYd0raED4btlvWx/Up2Iw3pOJb/cg4rm9t9Qj/lYBDA
Vya/dDM4HEBAnTN4F0AGl7mk5J6eH6Npd8oRk8cDXirZR1fXUTMSt4T4mOzoDBxNNFoEpPWrjq6y
65gRNE39SvDWw52nzRXB1I6FLn62HswSxh2lRuD1uJuPVQBYLwIkWC09JF1XBvuYlOXtI2vu1Go5
yH/dlWWIDirxv/qtmC4F0MDtI+MLmUYrp9sNsRRNUzuZpilxjmRbNSns07v4g0gRs/L5NzQD9JyG
fmKPdgvcdz4Ii8zDknJSAcyNnvrdV8xIOP7U/6lSBdNfdbU7GmIK52YCnwhWqWEbcl9d9VCTsVQP
2/b0hobgIyiS9gZlveJDPKkSvmNU3I2DL94PrsV0yvKXEifr7gOUNiSzgtyr4k84TZJpBUOLmRXt
M8WovG8Qu4ZC0bZ9HrKsTBN7EQncQITR4ZEyjxc6zxwD5zQlGnjnpyYv5gxBUI4ut2PV/ay/PwBb
42atPNJP9tEKwglrKiOl1uuB+6hY116fVQ6dOh4zS56AyE31+oWbGBpo9x8vfzrWgQcHmsvf2YkK
oFYdhigF4PbejdTDG7C+zjmFdhEQZ0Kv0+vb2ygi3jU95x3BaJfZgidulqFWWjkg62YKPYQ66ed3
P2ALZ5OOXaaBRiquzVrNzq2tGwFveEzewaHzXXgZDLlfvEceaUmT+UfXWax6mu3lkZ8La+xEueFB
TF7NqHv8o3ZrwbuBLkMxt5K7P/11B+hAq24gz8EwTy/tFW2oMFsZtYjCaM8mOSyglMZoQQlQpx2j
12IlEfDKdOM+roKPkZN2MJpMLBmp9JtnrY0UKr0auGuWUBHod0Vw2OM+VfbiBcxKeIkLMoD+FRKF
CM/IOBrU4EMRSueLx0IZRMa3tU7GCJbcTKfEwxwbZq5qiy7rv3N52oEmoT8duGhRDox2G3ZXKp2M
MDyXnp2F5YKyC4chP8wprwgNEih+OmQWfemHEWJrftm7vMwdv9ny2AtVJKNTOjAQz8iSqYLAA1Rn
8meE7+uAL4oOVYuiPkJ4hqTV4BDKaXdRjd2uUnUhOBW98g3YrUzw6lI5ZsZX7f5J/a1qIRXtiW34
1/MNuAIej6rf3fnZMrzeVI1r0T//I8J0j8OKbLsBqXJaauQUfiEmNQkemTTCpRLoq26nrEP6QkrV
TGh/0YDYx5FeOSsZT9mgaNKS0QQ4372czr6MzWKfwTrTqgCH6GMaJqJloaXpiHqMzzwGQRwDUb7W
J5QXRRExE2dXIbkYUakjKizNi6TyqRkHEQBXizP3r7gD4Jf+Bjlow8R0pyw0QcM/XENke+SIEzZc
fuLb4z+WrmtmGaMFlFxpHdXFW/yZOZO3zqCxDpEJ8uZQ/3lQidaum+Ckuo9tjQY0R4TAiyzVP2Ov
HG4GE6l5fQ8lXuXL/loDUKgxqEPKoQVslZy5/Ul59Sq0c+f1PcKubPZ/m9QgRE9QsCX+aWxzDVs0
9MBxnZn7Vfb00YFo2keIhm/SnKWT4Dyf/oIPsM5eWnlsRi+BSgpCrHShw6liY3vbdU9DFm7PM9la
jHLJTubkyfoGfnbOLC/FFOakhS8mmMRze5rpnPzR+sjdJdWi+77L3lGNR5RFo5tG25Nq3jlpEhry
lmziogU3f9vAH58384BEtF229P49wKFS7Jvh6hlT+5VRP5P+Vhz8TO7tgUHHp+lCYXIaWw3MRbMn
iUqvlKp4Jnu8N/PgVe/i0gWpDaLfm4WhziCI1WZDG//FwkXWKO8gRqVUOoNzTcrPXim2cz9U3M/2
mpgPFIpOOLfOxaod5uDJUdBfNWlxe8M9XKdBrqFDinD1ExZT6ghYsi9nK2Q7up7XgoQkfTpN8Hmv
DqufJCLMRcwVWaBU7F5JbvIbYcYHpZ7Zx34LxquwbQA8julBOvfyX/2wna+uIBhXNWuMcXS8Y3/e
id6DPrSuMq+regnhGwXbukYvOXChlaBRfemxHG2YUWDyLFVb16oUuUJOTFypiw9lQHJfBTlDXQYz
A65veTrnFx3+Grdt/i5sPvml/lxe4/mWM+gtkAvBZlbv4Hi4noX4WAL/XAyjP/KRTTm2PMwwRZi9
qNIK0ZpsYBNlNfp9KpRInwlEt7EOvt02Jbr6PswHtCLZCuh+vU7KTr2PeNXL2rZe1lr0lf0gRo/6
fZfGdxHmBCqBf/H9CCpPddvcjnfDY4cYI4NsVpStEFGXXLmGub/kY8iL/K7Mff4vO9ai4oGnJgqa
QhN+09hwbQ3Pw+UPcBYMZ7XK1CNS5xT87FW8g4jXvMiwpSyg5YtxqdclG0U24cxCCT3cG7Cuid4O
EO4gQmrDFhRZbrViowPo7WD4coCyIj9DRipHzlCPDFqCIH4COe3JC9lBUwrzgo1Gc7+sYOoGcDss
gxF92mvgC8A/PtyEUGX6Mn2iBssyETJhFhUJBCoZxQYKrkrJQEyL29JT3Oy8NDXijsY+u6HHdHFK
0X+eesTKqiH3Rkxsfj6c58GPocKrJkPAlk2BcZsSvvkW3W3s7nifZeigo1h5174NP/yvKsioNDFo
RFrVZhTpLmyB5eZ/of1AGtJbtV/Ixw8CuxJBJ+2bWe+nbiRjO4fmdhGlJ04+Fv9t/qZD4JF7mlGM
sMk62ABnCIhHrEQ1k6v4Vm2xVmNlIJfL25h1dgAmzt5/Or58f+Mqqw23EwH0D7O832x0SXp4vDit
r1PNFDIt0wakTQVa1Jjjs0P2Lajt+ehqCSZLQahlMbiew05gnQ2eO6q5Vml9eO82F6V8TebwUnW8
sAaOHAbbjYU0m0NiLfDebA637Gn+VPudbOjjBR5LD0zrSBGxCdUg6Tu2mpbfqTqXkYW9ieMDDVK3
HT3QHqpJ7DG4mfRtgwPciVUPYddWhEqZOEvAIaznwyhzHlSva8oTZ+dziPW91iYdXsuiTxi9eGgx
7m7SBBOp+juh2EHiozBr+VBGArDWjZwcjjGzxxi9q4D9Anw7TUpAmR5h9UfUdG06XhzNTKHb7s2K
tMWlGX7OEO++YecyZl2Mz5B/4C+xBdJPu8gloKNLVX96Z7Ejab9oNXdFWvXy779FlX5WOPN2d6L8
+Pn0gFa9PRfeuJFG5sZaMV9k2t03o8xXn6cDDmkvJ/D/SOSbuwJoOmXUTb5TS6LzIoZcbg0PMfMK
CuKJ/NKqYg+/snBL/44R+5lTXXW0FnUNE6nmD4iMltnJfCvHEgtt3hX6aIEhf3Cd4wrU7R/DKUTP
zgMbL6v2io0V/+LeeceL4qgoby/ktOm6J8RwL9pHyOsm6YMhc12KgjiUaOOuPVUJqBzxz81DiDby
yIW6rbATAb2GAOOlrOTe8TzKSeE4mwdVkTSTXndBJexcsOAytaWIrJKbVJIcxWlXwOBJfWDvD7KE
K2/5M4vk1U8JJG0d5dakWsfBCsf2R1BzryfDdYLV9mIEaOVR6wnPb/gY/hAgSokdU/qibnngxquK
DxHRrsWHsz9GH47xEAUHG17/QtQlau0m4g+lifY+o0FAcH+nG7a+OEypBUHjh7iN2GRQlGqIPExr
0su9chfWHNQ9JwxxSp3SFwr66mIvK2kX0Y8vBnI7z+E4kGvqWSni9o6810jcsI8gAm3oRdS8dKhf
+Pzh5NjZsmPEGApTxmbOpibIiAWOhlxW/PzI6F+LAqD8Lp05m+f1ombFYmbxOyPIUTRbhLlfq3uf
LqBqJBJcxJ4M7MkfLcxCbLbTGElb8MQfXXG3xBPJEwpNOvqJnI98HYOuPSV+BOjY89C4YiT195n6
2tM2BlFyCdOCtea1E+3sQ7syYVEzsgTJAnQfitDdcYoOaRyu8mORTCTKZJcVgejUX1/KgiAeEL9i
0Y7nT3a0Sn8COiEvc9nNVvgdiM8GJCXaickHbBTQo5hWHJfKmGfdhd9bn73LE6DLRVP+jpTYaIx/
MN5zWzGpgeN2tL5aQPrcTIuMFXjdvKeEhKpcDyngbDWEVAa16EvOgDaqUVg3M5Oe9GrnZ6NNp5bt
wgOrr6n4eWhz1/XtOVZhNYIZddPwOk8tDsCDiWhn3GBt+7ex80ka08F5NoQDP2IYqHiMkuqfvVMH
idr6eYUXG4ikQ7VCwKpveB/ebT7a8KxDEosI7Z5fPUp9zZccsCxRZN152phn3hmg4SARX0f0RkDn
Tvw7OqKEO3jhuLoozUu9IqqaqSAkcsuk6cveTThNOd/Mh9wPiMnOb3dRh2h7jf0lVZIg02XNw+io
bJHhIBc5siTf0oY8SoEWo+36l7DmMKLoagM6IVxFDwGIu6+rXY3bMM3uwv+JJQJ1qv5uC5nCESiy
s+aXcjHWsuU+IXuGGslQOlmM2qy3gywOtNNjM+kWx9N2a3Q8Blm4zCpJCowc5sadE7/3CnKBjNlr
iIdt7RyVNQWsgBuIEmg12gnWkI0+pLreMhybYQVs24U6DTcpSbTCMbs/GfDgsyy5SqFCMSlN22Xv
W+Lm1et9NvGifjggPtyyQdyjjf/et1fEDB0Wqa04oGUUVbXir/dMxHA4mu3hhAwMhrNsMuOQu7Kc
STWlZZMZzRXNJmK0Sv7rqh3nqJUkq3SQZ0dnv2t7ZvWtALc1DFew5fefY4elKOWw3MHIfdLWis48
6WqYn7nk0WcAnugCuTuSRsbPai9t+HqRMW4vJY8Z950uYekSBG0SHyq3/EhzqLsvZ9XhPIZ00KXW
dYzuCjcOOb+qUWR4xkITCAZpzLTxCWGTNf5QU6PgJztAw4ngvGB4Zn4qxqvNi/29q1wm4TFk+v8Z
dZqBtak6dv3dxV1cmog4frDxBRDWnanBXO0luZ70ahdECF7SLIsoKwEz98HzlXVGcO+pZOkjhNcl
Y2B7/SKtq1Yr1mw5lIH9ZWLmjjMrTocHo8FDZhjOOcPDf/jChVfboYREPzk57pq9ve21d/oVq5Gl
NCDndXNOw9wPdo8tGqCoLiYsIM2K865OiyFQM/hAr4GmNIhHdxBBdu4PVizkEU9Ipenck8ZOT39e
cqDbjbbfB9EHn4wKQgxN6GtBOLODOzpP6lYTW5tDQY2dsxyKrM8YFlejJGANdxqS+yNEIq35kPub
FK1x6ecnVZx2FlnuYKwtSX1e/p13fR8j3MSJVpR9lS6JRUSCdEeNlJXhlAnn6aoX/EZXzbqcoAaI
0bZyRVsp3kvc1EDtXF3mHl9dkmYFVQg/thRWrLSp8f1jK3fYvlpKVWIeXc1hnYtqngDReRb0jrqD
uU/xlcue27c1u0UL8UonQzU2HgPXOEk2a/fgjDRZJdw9+b5XBTNYD+V2FRnqIq/0gVv1gbYIT3vv
T04zXYdiAeLaK4b2i/wKnwVsIMHMmWLyFBVAT9uFKJXP2mTXrt7FpQKU0FHnh+fExUmB978VXbJV
axrvKr38rwcribZgAkBaVuGp6P0Kpuf3/yoL1Y5B9xyasnyFDlbojmeKVyoq8HXSX5ZhUKrd3XD9
ymA+jQZWoU0N79zW7ZqGkVDwOFBAHDpr/OW+Q68A5zHa9oGIS7IskUMXR11wZVubwsbyZlmE1fHf
XYFm20vEA/OWJFh1kXKv1UyjWw+Vsyg7STm5xeud20S8HXgl+xC7F0S4Ez8akgIxGz6ln3c0CiMC
LsBqNb+9gyIDkyk4vygvKNwOSo0VEP/WOuihxVeCtfkFxlF1Rgqyy0Gp/qtF1KblimylPmzp8CUm
u+Dt5z8hm/fVd3ISVjtcIuTxvNOPFYQ4XVGmKkXZiXHB2jYeD5eTImEZmq4tor4mHMkVHcxYTGwF
OfA1XU7wUlkeHvHS+7HpVoqJ5IS6A4HqAN19C6/Ciu2X7LSjdzJRNq2jCxQPA9Oni1u0wjhWJdd/
Z9+Xr26FqtYrCizqEtcGbdkxY3OHAbC8dNiQdcH0YvlQKfN7rUIPuhCM6GCITIwk8XAyur5fQq0q
7F1MtJtjuBq7NK1Gvh2c6fK1rJuxEPcrk+Ssa2E0qjp+ig89I+QJV5lL29gkLUQjVmTMxUoWzpoS
xRcJW3XEsnGeQUJe2ThATJ+761IVuw899FA9GJdrE3ZcXB7U0L/tInA8MsnzI2ngACRTEfc2jXvN
VyeAKcIoTmb9FL2hR9gZMlWJIOi0ukwny48lB37zHxhTUofXP4M5vap7ALIiyR54Ff3M61zETR+u
zfna6tDqX0hwYlpG0Ir/fTJLG5NAyctCvZcfMi/2tcbxiIToYExwiH4blIejnqHJOBgD+UIu+VIG
Dzl+CKZBDfBj4H6VVKHz2JKDGcvvpZKGcFo/1yHWsdjS/ruEar31K3TGE3ZRfYUHo4lI2whxOUMt
ZVbDuVTxQkGUc9Q5gkWoElrUbpGP17ZsZUYO6YqZo255/mwZDsDy3aE3TBRpk4AhXJHKMyFnTACk
ODj3KvtVb2TFcXyG7+ljRoQTEQwr8oL4cTstT0i0QOCVKuuyaD317mDi0h8DR9Ba97yVzU/x6dEi
w8IyUkdN/tgyLr0XZ0mieZADXpx68rFiD22/856tbLnOTy7aDj6Wo6D1W9vpm5wteso7xDn7/bGG
eJ5Ep1W1gIb9weRnPZ50OKhnEhbh7ANujQ+IZ0Ka7AarDY0IQ7JRIGmEEtDNkADE07iMyO5oLh5W
H3QLDeZPb3usHWe0EsKI0alSLgeAdveYDDD1MUfYrkTiPZYopxRj0MmUZc5SCOGsJexR9a8xjbXG
5UJBD148rdcwX+x2Gh/qktXSNeqVHsF1OUx/CvGre7FrJZ8weFbGNWyGXKX3R+n7Zx34kM73fwu9
pWEtaAyQuQ3bwOeEMV4hQ4CXlUC6U2//Gspbnpi8K/s7xCTqu3m8du2EHQabMXX9tUXEiDY3R8cI
T1rplAJzMtlrRefE52Fg9uPD36IlxhXguG/H6I0IIsW0gHmVDVvyvvm0hdabQK4DJ99Vm8ongf7f
uKNBtLc8ENUE8Z+3t5lOSn8fqRKcE8D/Ondfplz9N9EY+xZG5X/k8I6fPM4MX6my2tdzAmpojFxc
yqpp9tLEqq8tOft+qWd2eneoPXNenYtkVsR+UX8YeiLixsY4kyhakUIehmUGOzuy5LlTjatmuLBi
peF0rXVJFMHT4nrsHbqiXky90Rkzjgo+Nv6jv8irSThmGl5LpLVlkLpmVgkpYhu6H4fH2EVmDaBA
xkSI4qYau3geaWob49k5bAVZ9pdgjRe4YO3eJMt7h6SNmx0wtLyLi7wQb8EFv+T9G/PVG7iyvxPu
BUI93oyB8KDb00Q2s5y6Apz/4ULStEe1ha9fCBAQD9jQFFsxacjdH32KZJ8kvfKVk13dp3VTSSV/
VrZ4bi6xSajFA0jNRTNLNlNI8AoYE6kRursjxstHTxSO6pmKAWciRaIDbd6yt2cIFm9yBTCxGvyn
tWCJBbWW9wWShJZYeG6m8oXfQgHV2vz0DfzO6DLMqZznh+lJcCvR5kM5WG79jiY9gbOtnKc4Yipn
TAkxbl2Cuaur3bu4opGO0JfiyZFQ6NtS8X9H8HWrnGeWK1geVw43JFbwkf4j/MVJedELSslFQEGm
Uk5yj9ozg6SMUmpcjH97Td15jizAHZwcJxa8td1C9U3q7XiKqWjiOB0JdM/o9AV/K4jM7b25rF7n
WDVXItHCdA4EpQR8LinL9e5T35XFmNLES1kfOHOrDgCGC8/noBLWsCaVv2tTEbm/wrV9sJPQf8l+
FicIxnIcQX1yIrFh4s85qcn19EPSZ4ARV/5KXVkYVDcRYvcqoFGPKjHlIIT/DML0fB8wX76V+Mue
bwHdc6ygEqgT5lorj/UjOdKmruriTG2nzYQVaaDB/ROu6LaVtcuoFY35WSgmvJmmGc2O2ZY0+HjJ
CjTYWOSIc2Z449qp7V4p27DkOJ3VOEYdyA3tYLidRApqUQWx7p9Xm7sl5nK8Ay+sj7hs9AiLdaEG
DqaXkcW/eFkJdUgJELSX4U71VAwGBmxhQtbXy7akr8Ml9kc4Tqn3G5bjZQFdip4sKPwadv8y9J0R
fVWH0DUIV4rQRyNpTntkbGGJN7O1GehBEDitcgPaKEJeObnnMJzYn5Ig8zKvpvgr7wTiGT6vnCE/
ucUbX0ZW4N311MR2A2C/SQQ//iDvZoCOGqQW2u5dLsTUM+0HOEoGncogM26qxIzhf48SJM/iuS66
UtEk/qBEdnBWh6RpfgmkK5jMAs9BoksWmjEkid0dGAFMYXYpT/ZNJQAWtEpWxhIzCqfMdz8etEsE
CDbdG2iLwrkQxdIbvrQ=
`protect end_protected
